`timescale 1ns/1ns
import mMaskKron_package::*;

module mMaskKron(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Bool_src_d ,
  output logic \\QTree_Bool_src_r ,
  input QTree_Bool_t dummy_write_QTree_Bool_d,
  output logic dummy_write_QTree_Bool_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1acS_0_d,
  output logic m1acS_0_r,
  input Pointer_QTree_Bool_t m2acT_1_d,
  output logic m2acT_1_r,
  input Pointer_QTree_Bool_t m3acU_2_d,
  output logic m3acU_2_r,
  output \Word16#_t  forkHP1_QTree_Bool_snk_dout,
  input logic forkHP1_QTree_Bool_snk_rout,
  output Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_dout,
  input logic dummy_write_QTree_Bool_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Pointer_QTree_Bool_t main_mask_Bool_resbuf_dout,
  input logic main_mask_Bool_resbuf_rout
  );
  /* --define=INPUTS=((__05CQTree_Bool_src, 0, 1, Go), (dummy_write_QTree_Bool, 66, 73786976294838206464, QTree_Bool), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1acS_0, 16, 65536, Pointer_MaskQTree), (m2acT_1, 16, 65536, Pointer_QTree_Bool), (m3acU_2, 16, 65536, Pointer_QTree_Bool)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Bool_snk, 16, 65536, Word16__023), (dummy_write_QTree_Bool_sink, 16, 65536, Pointer_QTree_Bool), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (main_mask_Bool_resbuf, 16, 65536, Pointer_QTree_Bool)) */
  /* TYPE_START
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTmap__027__027_map__027__027_Bool_Bool_Bool 16 3 (0,[0]) (1,[16p,0,0,1,16p,16p,16p]) (2,[16p,16p,0,0,1,16p,16p]) (3,[16p,16p,16p,0,0,1,16p]) (4,[16p,16p,16p,16p])
CTkron_kron_Bool_Bool_Bool 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,0,0,16p,16p]) (4,[16p,16p,16p,16p])
CTmain_mask_Bool 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool 16 0 (0,[0,0,0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool 16 0 (0,[0,16p,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap__027__027_map__027__027_Bool_Bool_Bool 16 0 (0,[0,0,0,1,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,0,0,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_MaskQTree 16 0 (0,[0,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool 16 0 (0,[0,0,0,1,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  Go_t go_1_dummy_write_QTree_Bool_d;
  logic go_1_dummy_write_QTree_Bool_r;
  Go_t go_2_dummy_write_QTree_Bool_d;
  logic go_2_dummy_write_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_snk_d;
  logic forkHP1_QTree_Bool_snk_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  \Word16#_t  forkHP1_QTree_Boo4_d;
  logic forkHP1_QTree_Boo4_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  C3_t readMerge_choice_QTree_Bool_d;
  logic readMerge_choice_QTree_Bool_r;
  Pointer_QTree_Bool_t readMerge_data_QTree_Bool_d;
  logic readMerge_data_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_Boolm1acL_1_argbuf_d;
  logic readPointer_QTree_Boolm1acL_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_BoolmacD_1_argbuf_d;
  logic readPointer_QTree_BoolmacD_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolmaci_1_argbuf_d;
  logic readPointer_QTree_Boolmaci_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t destructReadOut_QTree_Bool_d;
  logic destructReadOut_QTree_Bool_r;
  C14_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_d;
  logic writeQTree_BoollizzieLet13_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_d;
  logic writeQTree_BoollizzieLet16_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_d;
  logic writeQTree_BoollizzieLet8_1_argbuf_r;
  Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_d;
  logic dummy_write_QTree_Bool_sink_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  \initHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \initHP_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \incrHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_CTmap''_map''_Bool_Bool_Bool1_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool1_r ;
  Go_t \incrHP_CTmap''_map''_Bool_Bool_Bool2_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool2_r ;
  \Word16#_t  \addHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \addHP_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Boo3_r ;
  C2_t \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memReadOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memReadOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memWriteOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memWriteOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \destructReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \dconPtr_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconPtr_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  initHP_CTkron_kron_Bool_Bool_Bool_d;
  logic initHP_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  incrHP_CTkron_kron_Bool_Bool_Bool_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_CTkron_kron_Bool_Bool_Bool1_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool1_r;
  Go_t incrHP_CTkron_kron_Bool_Bool_Bool2_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool2_r;
  \Word16#_t  addHP_CTkron_kron_Bool_Bool_Bool_d;
  logic addHP_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Bool_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Boo2_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Boo2_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Boo3_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Boo3_r;
  C2_t memMergeChoice_CTkron_kron_Bool_Bool_Bool_d;
  logic memMergeChoice_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memReadOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memReadOut_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memWriteOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memWriteOut_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r;
  \Word16#_t  destructReadIn_CTkron_kron_Bool_Bool_Bool_d;
  logic destructReadIn_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t dconReadIn_CTkron_kron_Bool_Bool_Bool_d;
  logic dconReadIn_CTkron_kron_Bool_Bool_Bool_r;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d;
  logic writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r;
  CTkron_kron_Bool_Bool_Bool_t writeMerge_data_CTkron_kron_Bool_Bool_Bool_d;
  logic writeMerge_data_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t dconWriteIn_CTkron_kron_Bool_Bool_Bool_d;
  logic dconWriteIn_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t dconPtr_CTkron_kron_Bool_Bool_Bool_d;
  logic dconPtr_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Pointer_CTkron_kron_Bool_Bool_Bool_t demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d;
  logic demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  initHP_CTmain_mask_Bool_d;
  logic initHP_CTmain_mask_Bool_r;
  \Word16#_t  incrHP_CTmain_mask_Bool_d;
  logic incrHP_CTmain_mask_Bool_r;
  Go_t incrHP_mergeCTmain_mask_Bool_d;
  logic incrHP_mergeCTmain_mask_Bool_r;
  Go_t incrHP_CTmain_mask_Bool1_d;
  logic incrHP_CTmain_mask_Bool1_r;
  Go_t incrHP_CTmain_mask_Bool2_d;
  logic incrHP_CTmain_mask_Bool2_r;
  \Word16#_t  addHP_CTmain_mask_Bool_d;
  logic addHP_CTmain_mask_Bool_r;
  \Word16#_t  mergeHP_CTmain_mask_Bool_d;
  logic mergeHP_CTmain_mask_Bool_r;
  Go_t incrHP_mergeCTmain_mask_Bool_buf_d;
  logic incrHP_mergeCTmain_mask_Bool_buf_r;
  \Word16#_t  mergeHP_CTmain_mask_Bool_buf_d;
  logic mergeHP_CTmain_mask_Bool_buf_r;
  \Word16#_t  forkHP1_CTmain_mask_Bool_d;
  logic forkHP1_CTmain_mask_Bool_r;
  \Word16#_t  forkHP1_CTmain_mask_Boo2_d;
  logic forkHP1_CTmain_mask_Boo2_r;
  \Word16#_t  forkHP1_CTmain_mask_Boo3_d;
  logic forkHP1_CTmain_mask_Boo3_r;
  C2_t memMergeChoice_CTmain_mask_Bool_d;
  logic memMergeChoice_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_d;
  logic memMergeIn_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_d;
  logic memOut_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memReadOut_CTmain_mask_Bool_d;
  logic memReadOut_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memWriteOut_CTmain_mask_Bool_d;
  logic memWriteOut_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_dbuf_d;
  logic memMergeIn_CTmain_mask_Bool_dbuf_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_rbuf_d;
  logic memMergeIn_CTmain_mask_Bool_rbuf_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_dbuf_d;
  logic memOut_CTmain_mask_Bool_dbuf_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_rbuf_d;
  logic memOut_CTmain_mask_Bool_rbuf_r;
  \Word16#_t  destructReadIn_CTmain_mask_Bool_d;
  logic destructReadIn_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t dconReadIn_CTmain_mask_Bool_d;
  logic dconReadIn_CTmain_mask_Bool_r;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CTmain_mask_Bool_d;
  logic writeMerge_choice_CTmain_mask_Bool_r;
  CTmain_mask_Bool_t writeMerge_data_CTmain_mask_Bool_d;
  logic writeMerge_data_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet28_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet9_1_argbuf_r;
  MemIn_CTmain_mask_Bool_t dconWriteIn_CTmain_mask_Bool_d;
  logic dconWriteIn_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t dconPtr_CTmain_mask_Bool_d;
  logic dconPtr_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  Pointer_CTmain_mask_Bool_t demuxWriteResult_CTmain_mask_Bool_d;
  logic demuxWriteResult_CTmain_mask_Bool_r;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreemskacj_1_argbuf_d;
  logic readPointer_MaskQTreemskacj_1_argbuf_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r;
  MyDTBool_Bool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r;
  MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r;
  MyDTBool_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTBool_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTBool_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t es_0_1_1_d;
  logic es_0_1_1_r;
  MyBool_t es_0_1_2_d;
  logic es_0_1_2_r;
  MyBool_t es_0_1_3_d;
  logic es_0_1_3_r;
  Go_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r;
  MyDTBool_Bool_Bool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_r;
  MyDTBool_Bool_Bool_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTBool_Bool_Bool_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTBool_Bool_Bool_t arg0_2_3_d;
  logic arg0_2_3_r;
  MyDTBool_Bool_Bool_t arg0_2_4_d;
  logic arg0_2_4_r;
  MyBool_t xabY_1_d;
  logic xabY_1_r;
  MyBool_t xabY_2_d;
  logic xabY_2_r;
  MyBool_t arg0_1Dcon_main1_d;
  logic arg0_1Dcon_main1_r;
  MyBool_t arg0_1Dcon_main1_1_d;
  logic arg0_1Dcon_main1_1_r;
  MyBool_t arg0_1Dcon_main1_2_d;
  logic arg0_1Dcon_main1_2_r;
  Go_t arg0_1Dcon_main1_1MyFalse_d;
  logic arg0_1Dcon_main1_1MyFalse_r;
  Go_t arg0_1Dcon_main1_1MyTrue_d;
  logic arg0_1Dcon_main1_1MyTrue_r;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTrue_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTrue_r;
  MyBool_t applyfnBool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_5_resbuf_r;
  MyBool_t arg0_1Dcon_main1_1MyTrue_1MyFalse_d;
  logic arg0_1Dcon_main1_1MyTrue_1MyFalse_r;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r;
  Go_t arg0_2Dcon_main1_d;
  logic arg0_2Dcon_main1_r;
  MyBool_t \arg0_2_1Dcon_&&_d ;
  logic \arg0_2_1Dcon_&&_r ;
  MyBool_t \arg0_2_2Dcon_&&_d ;
  logic \arg0_2_2Dcon_&&_r ;
  MyBool_t \arg0_2_2Dcon_&&_1_d ;
  logic \arg0_2_2Dcon_&&_1_r ;
  MyBool_t \arg0_2_2Dcon_&&_2_d ;
  logic \arg0_2_2Dcon_&&_2_r ;
  MyBool_t \arg0_2_2Dcon_&&_3_d ;
  logic \arg0_2_2Dcon_&&_3_r ;
  MyBool_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  MyBool_t \arg0_2_2Dcon_&&_1MyTrue_d ;
  logic \arg0_2_2Dcon_&&_1MyTrue_r ;
  Go_t \arg0_2_2Dcon_&&_2MyFalse_d ;
  logic \arg0_2_2Dcon_&&_2MyFalse_r ;
  Go_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  MyBool_t \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_d ;
  logic \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_r ;
  MyBool_t applyfnBool_Bool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_Bool_5_resbuf_r;
  MyBool_t \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d ;
  logic \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_r ;
  Go_t \arg0_2_3Dcon_&&_d ;
  logic \arg0_2_3Dcon_&&_r ;
  MyBool_t \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_d ;
  logic \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_r ;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r;
  Go_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_r;
  MyDTBool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_r;
  MyDTBool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r;
  Go_t call_kron_kron_Bool_Bool_Bool_initBufi_d;
  logic call_kron_kron_Bool_Bool_Bool_initBufi_r;
  C5_t go_4_goMux_choice_d;
  logic go_4_goMux_choice_r;
  Go_t go_4_goMux_data_d;
  logic go_4_goMux_data_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork1_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork1_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork2_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork2_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork3_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork3_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork4_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork4_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork5_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork5_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork6_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork6_r;
  Go_t call_kron_kron_Bool_Bool_Bool_initBuf_d;
  logic call_kron_kron_Bool_Bool_Bool_initBuf_r;
  Go_t call_kron_kron_Bool_Bool_Bool_goMux1_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux1_r;
  MyDTBool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux2_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux2_r;
  MyDTBool_Bool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux3_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux3_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_Bool_goMux4_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux4_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_Bool_goMux5_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux5_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux6_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux6_r;
  Go_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r;
  Pointer_QTree_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_r;
  Pointer_MaskQTree_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_r;
  Pointer_CTmain_mask_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r;
  Go_t call_main_mask_Bool_initBufi_d;
  logic call_main_mask_Bool_initBufi_r;
  C5_t go_5_goMux_choice_d;
  logic go_5_goMux_choice_r;
  Go_t go_5_goMux_data_d;
  logic go_5_goMux_data_r;
  Go_t call_main_mask_Bool_unlockFork1_d;
  logic call_main_mask_Bool_unlockFork1_r;
  Go_t call_main_mask_Bool_unlockFork2_d;
  logic call_main_mask_Bool_unlockFork2_r;
  Go_t call_main_mask_Bool_unlockFork3_d;
  logic call_main_mask_Bool_unlockFork3_r;
  Go_t call_main_mask_Bool_unlockFork4_d;
  logic call_main_mask_Bool_unlockFork4_r;
  Go_t call_main_mask_Bool_initBuf_d;
  logic call_main_mask_Bool_initBuf_r;
  Go_t call_main_mask_Bool_goMux1_d;
  logic call_main_mask_Bool_goMux1_r;
  Pointer_QTree_Bool_t call_main_mask_Bool_goMux2_d;
  logic call_main_mask_Bool_goMux2_r;
  Pointer_MaskQTree_t call_main_mask_Bool_goMux3_d;
  logic call_main_mask_Bool_goMux3_r;
  Pointer_CTmain_mask_Bool_t call_main_mask_Bool_goMux4_d;
  logic call_main_mask_Bool_goMux4_r;
  Go_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_r ;
  MyDTBool_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_r ;
  MyDTBool_Bool_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_r ;
  MyBool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_r ;
  Pointer_QTree_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_initBufi_d ;
  logic \call_map''_map''_Bool_Bool_Bool_initBufi_r ;
  C5_t go_6_goMux_choice_d;
  logic go_6_goMux_choice_r;
  Go_t go_6_goMux_data_d;
  logic go_6_goMux_data_r;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork1_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork1_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork2_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork3_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork3_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork4_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork4_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork5_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork5_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork6_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork6_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_initBuf_d ;
  logic \call_map''_map''_Bool_Bool_Bool_initBuf_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_goMux1_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux1_r ;
  MyDTBool_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux2_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux2_r ;
  MyDTBool_Bool_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux3_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux3_r ;
  MyBool_t \call_map''_map''_Bool_Bool_Bool_goMux4_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux4_r ;
  Pointer_QTree_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux5_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux5_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_Bool_goMux6_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux6_r ;
  Go_t es_0_1_1MyFalse_d;
  logic es_0_1_1MyFalse_r;
  Go_t es_0_1_1MyTrue_d;
  logic es_0_1_1MyTrue_r;
  Go_t es_0_1_1MyFalse_1_argbuf_d;
  logic es_0_1_1MyFalse_1_argbuf_r;
  Go_t es_0_1_1MyTrue_1_d;
  logic es_0_1_1MyTrue_1_r;
  Go_t es_0_1_1MyTrue_2_d;
  logic es_0_1_1MyTrue_2_r;
  QTree_Bool_t es_0_1_1MyTrue_1QNone_Bool_d;
  logic es_0_1_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t es_0_1_1MyTrue_2_argbuf_d;
  logic es_0_1_1MyTrue_2_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyFalse_d;
  logic es_0_1_2MyFalse_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyTrue_d;
  logic es_0_1_2MyTrue_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyFalse_1_argbuf_d;
  logic es_0_1_2MyFalse_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyTrue_1_argbuf_d;
  logic es_0_1_2MyTrue_1_argbuf_r;
  MyBool_t es_0_1_3MyFalse_d;
  logic es_0_1_3MyFalse_r;
  MyBool_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  QTree_Bool_t es_0_1_3MyFalse_1QVal_Bool_d;
  logic es_0_1_3MyFalse_1QVal_Bool_r;
  QTree_Bool_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  MyDTBool_Bool_Bool_t gacB_2_2_argbuf_d;
  logic gacB_2_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacB_2_1_d;
  logic gacB_2_1_r;
  MyDTBool_Bool_Bool_t gacB_2_2_d;
  logic gacB_2_2_r;
  MyDTBool_Bool_Bool_t gacB_3_2_argbuf_d;
  logic gacB_3_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacB_3_1_d;
  logic gacB_3_1_r;
  MyDTBool_Bool_Bool_t gacB_3_2_d;
  logic gacB_3_2_r;
  MyDTBool_Bool_Bool_t gacB_4_1_argbuf_d;
  logic gacB_4_1_argbuf_r;
  MyDTBool_Bool_Bool_t gacK_2_2_argbuf_d;
  logic gacK_2_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacK_2_1_d;
  logic gacK_2_1_r;
  MyDTBool_Bool_Bool_t gacK_2_2_d;
  logic gacK_2_2_r;
  MyDTBool_Bool_Bool_t gacK_3_2_argbuf_d;
  logic gacK_3_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacK_3_1_d;
  logic gacK_3_1_r;
  MyDTBool_Bool_Bool_t gacK_3_2_d;
  logic gacK_3_2_r;
  MyDTBool_Bool_Bool_t gacK_4_1_argbuf_d;
  logic gacK_4_1_argbuf_r;
  MyDTBool_Bool_Bool_t \go_1Dcon_&&_d ;
  logic \go_1Dcon_&&_r ;
  C4_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C4_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C6_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C6_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C5_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C5_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  MyDTBool_Bool_Bool_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  MyDTBool_Bool_t go_2Dcon_main1_d;
  logic go_2Dcon_main1_r;
  MyDTBool_Bool_t es_2_1_argbuf_d;
  logic es_2_1_argbuf_r;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r;
  Go_t go_4_argbuf_d;
  logic go_4_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r;
  C5_t go_4_goMux_choice_1_d;
  logic go_4_goMux_choice_1_r;
  C5_t go_4_goMux_choice_2_d;
  logic go_4_goMux_choice_2_r;
  C5_t go_4_goMux_choice_3_d;
  logic go_4_goMux_choice_3_r;
  C5_t go_4_goMux_choice_4_d;
  logic go_4_goMux_choice_4_r;
  C5_t go_4_goMux_choice_5_d;
  logic go_4_goMux_choice_5_r;
  MyDTBool_Bool_t isZacJ_goMux_mux_d;
  logic isZacJ_goMux_mux_r;
  MyDTBool_Bool_Bool_t gacK_goMux_mux_d;
  logic gacK_goMux_mux_r;
  Pointer_QTree_Bool_t m1acL_goMux_mux_d;
  logic m1acL_goMux_mux_r;
  Pointer_QTree_Bool_t m2acM_goMux_mux_d;
  logic m2acM_goMux_mux_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_5_goMux_choice_1_d;
  logic go_5_goMux_choice_1_r;
  C5_t go_5_goMux_choice_2_d;
  logic go_5_goMux_choice_2_r;
  C5_t go_5_goMux_choice_3_d;
  logic go_5_goMux_choice_3_r;
  Pointer_QTree_Bool_t maci_goMux_mux_d;
  logic maci_goMux_mux_r;
  Pointer_MaskQTree_t mskacj_goMux_mux_d;
  logic mskacj_goMux_mux_r;
  Pointer_CTmain_mask_Bool_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_6_goMux_choice_1_d;
  logic go_6_goMux_choice_1_r;
  C5_t go_6_goMux_choice_2_d;
  logic go_6_goMux_choice_2_r;
  C5_t go_6_goMux_choice_3_d;
  logic go_6_goMux_choice_3_r;
  C5_t go_6_goMux_choice_4_d;
  logic go_6_goMux_choice_4_r;
  C5_t go_6_goMux_choice_5_d;
  logic go_6_goMux_choice_5_r;
  MyDTBool_Bool_t isZacA_goMux_mux_d;
  logic isZacA_goMux_mux_r;
  MyDTBool_Bool_Bool_t gacB_goMux_mux_d;
  logic gacB_goMux_mux_r;
  MyBool_t \v'acC_goMux_mux_d ;
  logic \v'acC_goMux_mux_r ;
  Pointer_QTree_Bool_t macD_goMux_mux_d;
  logic macD_goMux_mux_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  CTkron_kron_Bool_Bool_Bool_t go_7_1Lkron_kron_Bool_Bool_Boolsbos_d;
  logic go_7_1Lkron_kron_Bool_Bool_Boolsbos_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t go_7_2_argbuf_d;
  logic go_7_2_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r;
  CTmain_mask_Bool_t go_8_1Lmain_mask_Boolsbos_d;
  logic go_8_1Lmain_mask_Boolsbos_r;
  CTmain_mask_Bool_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t go_8_2_argbuf_d;
  logic go_8_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_d ;
  logic \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Go_t go_9_2_argbuf_d;
  logic go_9_2_argbuf_r;
  \TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r ;
  MyDTBool_Bool_t isZacA_2_2_argbuf_d;
  logic isZacA_2_2_argbuf_r;
  MyDTBool_Bool_t isZacA_2_1_d;
  logic isZacA_2_1_r;
  MyDTBool_Bool_t isZacA_2_2_d;
  logic isZacA_2_2_r;
  MyDTBool_Bool_t isZacA_3_2_argbuf_d;
  logic isZacA_3_2_argbuf_r;
  MyDTBool_Bool_t isZacA_3_1_d;
  logic isZacA_3_1_r;
  MyDTBool_Bool_t isZacA_3_2_d;
  logic isZacA_3_2_r;
  MyDTBool_Bool_t isZacA_4_1_argbuf_d;
  logic isZacA_4_1_argbuf_r;
  MyDTBool_Bool_t isZacJ_2_2_argbuf_d;
  logic isZacJ_2_2_argbuf_r;
  MyDTBool_Bool_t isZacJ_2_1_d;
  logic isZacJ_2_1_r;
  MyDTBool_Bool_t isZacJ_2_2_d;
  logic isZacJ_2_2_r;
  MyDTBool_Bool_t isZacJ_3_2_argbuf_d;
  logic isZacJ_3_2_argbuf_r;
  MyDTBool_Bool_t isZacJ_3_1_d;
  logic isZacJ_3_1_r;
  MyDTBool_Bool_t isZacJ_3_2_d;
  logic isZacJ_3_2_r;
  MyDTBool_Bool_t isZacJ_4_1_argbuf_d;
  logic isZacJ_4_1_argbuf_r;
  Go_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_r;
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_r;
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_r;
  MyDTBool_Bool_Bool_t gacK_1_1_argbuf_d;
  logic gacK_1_1_argbuf_r;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  MyDTBool_Bool_t isZacJ_1_1_argbuf_d;
  logic isZacJ_1_1_argbuf_r;
  Pointer_QTree_Bool_t m1acL_1_1_argbuf_d;
  logic m1acL_1_1_argbuf_r;
  Pointer_QTree_Bool_t m2acM_1_1_argbuf_d;
  logic m2acM_1_1_argbuf_r;
  Pointer_QTree_Bool_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  Pointer_QTree_Bool_t q1acO_destruct_d;
  logic q1acO_destruct_r;
  Pointer_QTree_Bool_t q2acP_destruct_d;
  logic q2acP_destruct_r;
  Pointer_QTree_Bool_t q3acQ_destruct_d;
  logic q3acQ_destruct_r;
  Pointer_QTree_Bool_t q4acR_destruct_d;
  logic q4acR_destruct_r;
  MyBool_t vacN_destruct_d;
  logic vacN_destruct_r;
  QTree_Bool_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  QTree_Bool_t lizzieLet0_1QVal_Bool_d;
  logic lizzieLet0_1QVal_Bool_r;
  QTree_Bool_t lizzieLet0_1QNode_Bool_d;
  logic lizzieLet0_1QNode_Bool_r;
  QTree_Bool_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  MyDTBool_Bool_Bool_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet0_3QVal_Bool_d;
  logic lizzieLet0_3QVal_Bool_r;
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_d;
  logic lizzieLet0_3QNode_Bool_r;
  MyDTBool_Bool_Bool_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_1_d;
  logic lizzieLet0_3QNode_Bool_1_r;
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_2_d;
  logic lizzieLet0_3QNode_Bool_2_r;
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_2_argbuf_d;
  logic lizzieLet0_3QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_Bool_t lizzieLet0_3QVal_Bool_1_argbuf_d;
  logic lizzieLet0_3QVal_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_r;
  Go_t lizzieLet0_4QVal_Bool_d;
  logic lizzieLet0_4QVal_Bool_r;
  Go_t lizzieLet0_4QNode_Bool_d;
  logic lizzieLet0_4QNode_Bool_r;
  Go_t lizzieLet0_4QError_Bool_d;
  logic lizzieLet0_4QError_Bool_r;
  Go_t lizzieLet0_4QError_Bool_1_d;
  logic lizzieLet0_4QError_Bool_1_r;
  Go_t lizzieLet0_4QError_Bool_2_d;
  logic lizzieLet0_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QError_Bool_1QError_Bool_d;
  logic lizzieLet0_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet3_1_argbuf_d;
  logic lizzieLet3_1_argbuf_r;
  Go_t lizzieLet0_4QError_Bool_2_argbuf_d;
  logic lizzieLet0_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet0_4QNode_Bool_1_argbuf_d;
  logic lizzieLet0_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_1_d;
  logic lizzieLet0_4QNone_Bool_1_r;
  Go_t lizzieLet0_4QNone_Bool_2_d;
  logic lizzieLet0_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet0_4QNone_Bool_1QNone_Bool_d;
  logic lizzieLet0_4QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet1_1_argbuf_d;
  logic lizzieLet1_1_argbuf_r;
  Go_t lizzieLet0_4QNone_Bool_2_argbuf_d;
  logic lizzieLet0_4QNone_Bool_2_argbuf_r;
  C4_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t lizzieLet0_4QVal_Bool_1_d;
  logic lizzieLet0_4QVal_Bool_1_r;
  Go_t lizzieLet0_4QVal_Bool_2_d;
  logic lizzieLet0_4QVal_Bool_2_r;
  Go_t lizzieLet0_4QVal_Bool_1_argbuf_d;
  logic lizzieLet0_4QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r ;
  Go_t lizzieLet0_4QVal_Bool_2_argbuf_d;
  logic lizzieLet0_4QVal_Bool_2_argbuf_r;
  MyDTBool_Bool_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  MyDTBool_Bool_t lizzieLet0_5QVal_Bool_d;
  logic lizzieLet0_5QVal_Bool_r;
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_d;
  logic lizzieLet0_5QNode_Bool_r;
  MyDTBool_Bool_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_1_d;
  logic lizzieLet0_5QNode_Bool_1_r;
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_2_d;
  logic lizzieLet0_5QNode_Bool_2_r;
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_2_argbuf_d;
  logic lizzieLet0_5QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_t lizzieLet0_5QVal_Bool_1_argbuf_d;
  logic lizzieLet0_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_6QVal_Bool_d;
  logic lizzieLet0_6QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_d;
  logic lizzieLet0_6QNode_Bool_r;
  Pointer_QTree_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_1_d;
  logic lizzieLet0_6QNode_Bool_1_r;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_2_d;
  logic lizzieLet0_6QNode_Bool_2_r;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_2_argbuf_d;
  logic lizzieLet0_6QNode_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet0_6QVal_Bool_1_argbuf_d;
  logic lizzieLet0_6QVal_Bool_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNone_Bool_d;
  logic lizzieLet0_7QNone_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QVal_Bool_d;
  logic lizzieLet0_7QVal_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNode_Bool_d;
  logic lizzieLet0_7QNode_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QError_Bool_d;
  logic lizzieLet0_7QError_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QError_Bool_1_argbuf_d;
  logic lizzieLet0_7QError_Bool_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNone_Bool_1_argbuf_d;
  logic lizzieLet0_7QNone_Bool_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QVal_Bool_1_argbuf_d;
  logic lizzieLet0_7QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t q1acF_destruct_d;
  logic q1acF_destruct_r;
  Pointer_QTree_Bool_t q2acG_destruct_d;
  logic q2acG_destruct_r;
  Pointer_QTree_Bool_t q3acH_destruct_d;
  logic q3acH_destruct_r;
  Pointer_QTree_Bool_t q4acI_destruct_d;
  logic q4acI_destruct_r;
  MyBool_t vacE_destruct_d;
  logic vacE_destruct_r;
  QTree_Bool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  QTree_Bool_t lizzieLet11_1_1QVal_Bool_d;
  logic lizzieLet11_1_1QVal_Bool_r;
  QTree_Bool_t lizzieLet11_1_1QNode_Bool_d;
  logic lizzieLet11_1_1QNode_Bool_r;
  QTree_Bool_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  MyDTBool_Bool_Bool_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QVal_Bool_d;
  logic lizzieLet11_1_3QVal_Bool_r;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_d;
  logic lizzieLet11_1_3QNode_Bool_r;
  MyDTBool_Bool_Bool_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_1_d;
  logic lizzieLet11_1_3QNode_Bool_1_r;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_2_d;
  logic lizzieLet11_1_3QNode_Bool_2_r;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_2_argbuf_d;
  logic lizzieLet11_1_3QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QVal_Bool_1_argbuf_d;
  logic lizzieLet11_1_3QVal_Bool_1_argbuf_r;
  Go_t lizzieLet11_1_4QNone_Bool_d;
  logic lizzieLet11_1_4QNone_Bool_r;
  Go_t lizzieLet11_1_4QVal_Bool_d;
  logic lizzieLet11_1_4QVal_Bool_r;
  Go_t lizzieLet11_1_4QNode_Bool_d;
  logic lizzieLet11_1_4QNode_Bool_r;
  Go_t lizzieLet11_1_4QError_Bool_d;
  logic lizzieLet11_1_4QError_Bool_r;
  Go_t lizzieLet11_1_4QError_Bool_1_d;
  logic lizzieLet11_1_4QError_Bool_1_r;
  Go_t lizzieLet11_1_4QError_Bool_2_d;
  logic lizzieLet11_1_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet11_1_4QError_Bool_1QError_Bool_d;
  logic lizzieLet11_1_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t lizzieLet11_1_4QError_Bool_2_argbuf_d;
  logic lizzieLet11_1_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet11_1_4QNode_Bool_1_argbuf_d;
  logic lizzieLet11_1_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet11_1_4QNone_Bool_1_d;
  logic lizzieLet11_1_4QNone_Bool_1_r;
  Go_t lizzieLet11_1_4QNone_Bool_2_d;
  logic lizzieLet11_1_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet11_1_4QNone_Bool_1QNone_Bool_d;
  logic lizzieLet11_1_4QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Go_t lizzieLet11_1_4QNone_Bool_2_argbuf_d;
  logic lizzieLet11_1_4QNone_Bool_2_argbuf_r;
  C5_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t lizzieLet11_1_4QVal_Bool_1_d;
  logic lizzieLet11_1_4QVal_Bool_1_r;
  Go_t lizzieLet11_1_4QVal_Bool_2_d;
  logic lizzieLet11_1_4QVal_Bool_2_r;
  Go_t lizzieLet11_1_4QVal_Bool_3_d;
  logic lizzieLet11_1_4QVal_Bool_3_r;
  Go_t lizzieLet11_1_4QVal_Bool_1_argbuf_d;
  logic lizzieLet11_1_4QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r;
  Go_t lizzieLet11_1_4QVal_Bool_2_argbuf_d;
  logic lizzieLet11_1_4QVal_Bool_2_argbuf_r;
  TupGo___MyDTBool_Bool___MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r;
  MyDTBool_Bool_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTBool_Bool_t lizzieLet11_1_5QVal_Bool_d;
  logic lizzieLet11_1_5QVal_Bool_r;
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_d;
  logic lizzieLet11_1_5QNode_Bool_r;
  MyDTBool_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_1_d;
  logic lizzieLet11_1_5QNode_Bool_1_r;
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_2_d;
  logic lizzieLet11_1_5QNode_Bool_2_r;
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_2_argbuf_d;
  logic lizzieLet11_1_5QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_t lizzieLet11_1_5QVal_Bool_1_argbuf_d;
  logic lizzieLet11_1_5QVal_Bool_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QNone_Bool_d;
  logic lizzieLet11_1_6QNone_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QVal_Bool_d;
  logic lizzieLet11_1_6QVal_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QNode_Bool_d;
  logic lizzieLet11_1_6QNode_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QError_Bool_d;
  logic lizzieLet11_1_6QError_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QError_Bool_1_argbuf_d;
  logic lizzieLet11_1_6QError_Bool_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QNone_Bool_1_argbuf_d;
  logic lizzieLet11_1_6QNone_Bool_1_argbuf_r;
  MyBool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyBool_t lizzieLet11_1_7QVal_Bool_d;
  logic lizzieLet11_1_7QVal_Bool_r;
  MyBool_t lizzieLet11_1_7QNode_Bool_d;
  logic lizzieLet11_1_7QNode_Bool_r;
  MyBool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  MyBool_t lizzieLet11_1_7QNode_Bool_1_d;
  logic lizzieLet11_1_7QNode_Bool_1_r;
  MyBool_t lizzieLet11_1_7QNode_Bool_2_d;
  logic lizzieLet11_1_7QNode_Bool_2_r;
  MyBool_t lizzieLet11_1_7QNode_Bool_2_argbuf_d;
  logic lizzieLet11_1_7QNode_Bool_2_argbuf_r;
  MyBool_t lizzieLet11_1_7QVal_Bool_1_argbuf_d;
  logic lizzieLet11_1_7QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t es_1_destruct_d;
  logic es_1_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  MyDTBool_Bool_t isZacJ_4_destruct_d;
  logic isZacJ_4_destruct_r;
  MyDTBool_Bool_Bool_t gacK_4_destruct_d;
  logic gacK_4_destruct_r;
  Pointer_QTree_Bool_t q1acO_3_destruct_d;
  logic q1acO_3_destruct_r;
  Pointer_QTree_Bool_t m2acM_4_destruct_d;
  logic m2acM_4_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  MyDTBool_Bool_t isZacJ_3_destruct_d;
  logic isZacJ_3_destruct_r;
  MyDTBool_Bool_Bool_t gacK_3_destruct_d;
  logic gacK_3_destruct_r;
  Pointer_QTree_Bool_t q1acO_2_destruct_d;
  logic q1acO_2_destruct_r;
  Pointer_QTree_Bool_t m2acM_3_destruct_d;
  logic m2acM_3_destruct_r;
  Pointer_QTree_Bool_t q2acP_2_destruct_d;
  logic q2acP_2_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  MyDTBool_Bool_t isZacJ_2_destruct_d;
  logic isZacJ_2_destruct_r;
  MyDTBool_Bool_Bool_t gacK_2_destruct_d;
  logic gacK_2_destruct_r;
  Pointer_QTree_Bool_t q1acO_1_destruct_d;
  logic q1acO_1_destruct_r;
  Pointer_QTree_Bool_t m2acM_2_destruct_d;
  logic m2acM_2_destruct_r;
  Pointer_QTree_Bool_t q2acP_1_destruct_d;
  logic q2acP_1_destruct_r;
  Pointer_QTree_Bool_t q3acQ_1_destruct_d;
  logic q3acQ_1_destruct_r;
  CTkron_kron_Bool_Bool_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_r;
  Go_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d;
  logic lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_r;
  QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_r;
  QTree_Bool_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d;
  logic lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d;
  logic lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r;
  Go_t call_kron_kron_Bool_Bool_Bool_goConst_d;
  logic call_kron_kron_Bool_Bool_Bool_goConst_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_d;
  logic kron_kron_Bool_Bool_Bool_resbuf_r;
  Pointer_QTree_Bool_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Bool_t es_2_4_destruct_d;
  logic es_2_4_destruct_r;
  Pointer_QTree_Bool_t es_3_6_destruct_d;
  logic es_3_6_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Bool_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Bool_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Bool_t t1acp_3_destruct_d;
  logic t1acp_3_destruct_r;
  Pointer_MaskQTree_t q1ack_3_destruct_d;
  logic q1ack_3_destruct_r;
  Pointer_QTree_Bool_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Bool_t t1acp_2_destruct_d;
  logic t1acp_2_destruct_r;
  Pointer_MaskQTree_t q1ack_2_destruct_d;
  logic q1ack_2_destruct_r;
  Pointer_QTree_Bool_t t2acq_2_destruct_d;
  logic t2acq_2_destruct_r;
  Pointer_MaskQTree_t q2acl_2_destruct_d;
  logic q2acl_2_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Bool_t t1acp_1_destruct_d;
  logic t1acp_1_destruct_r;
  Pointer_MaskQTree_t q1ack_1_destruct_d;
  logic q1ack_1_destruct_r;
  Pointer_QTree_Bool_t t2acq_1_destruct_d;
  logic t2acq_1_destruct_r;
  Pointer_MaskQTree_t q2acl_1_destruct_d;
  logic q2acl_1_destruct_r;
  Pointer_QTree_Bool_t t3acr_1_destruct_d;
  logic t3acr_1_destruct_r;
  Pointer_MaskQTree_t q3acm_1_destruct_d;
  logic q3acm_1_destruct_r;
  CTmain_mask_Bool_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  CTmain_mask_Bool_t lizzieLet25_1Lcall_main_mask_Bool3_d;
  logic lizzieLet25_1Lcall_main_mask_Bool3_r;
  CTmain_mask_Bool_t lizzieLet25_1Lcall_main_mask_Bool2_d;
  logic lizzieLet25_1Lcall_main_mask_Bool2_r;
  CTmain_mask_Bool_t lizzieLet25_1Lcall_main_mask_Bool1_d;
  logic lizzieLet25_1Lcall_main_mask_Bool1_r;
  CTmain_mask_Bool_t lizzieLet25_1Lcall_main_mask_Bool0_d;
  logic lizzieLet25_1Lcall_main_mask_Bool0_r;
  Go_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Go_t lizzieLet25_3Lcall_main_mask_Bool3_d;
  logic lizzieLet25_3Lcall_main_mask_Bool3_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool2_d;
  logic lizzieLet25_3Lcall_main_mask_Bool2_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool1_d;
  logic lizzieLet25_3Lcall_main_mask_Bool1_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool0_d;
  logic lizzieLet25_3Lcall_main_mask_Bool0_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_d;
  logic lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_d;
  logic lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_d;
  logic lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_r;
  Go_t lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_d;
  logic lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lmain_mask_Boolsbos_d;
  logic lizzieLet25_4Lmain_mask_Boolsbos_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool3_d;
  logic lizzieLet25_4Lcall_main_mask_Bool3_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool2_d;
  logic lizzieLet25_4Lcall_main_mask_Bool2_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool1_d;
  logic lizzieLet25_4Lcall_main_mask_Bool1_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool0_d;
  logic lizzieLet25_4Lcall_main_mask_Bool0_r;
  QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_d;
  logic lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_r;
  QTree_Bool_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_d;
  logic lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_r;
  CTmain_mask_Bool_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_d;
  logic lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_r;
  CTmain_mask_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_d;
  logic lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_r;
  CTmain_mask_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d;
  logic lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d;
  logic lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r;
  Go_t call_main_mask_Bool_goConst_d;
  logic call_main_mask_Bool_goConst_r;
  Pointer_QTree_Bool_t main_mask_Bool_resbuf_d;
  logic main_mask_Bool_resbuf_r;
  Pointer_QTree_Bool_t es_2_5_destruct_d;
  logic es_2_5_destruct_r;
  Pointer_QTree_Bool_t es_3_8_destruct_d;
  logic es_3_8_destruct_r;
  Pointer_QTree_Bool_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Bool_t es_3_7_destruct_d;
  logic es_3_7_destruct_r;
  Pointer_QTree_Bool_t es_4_1_destruct_d;
  logic es_4_1_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  MyDTBool_Bool_t isZacA_4_destruct_d;
  logic isZacA_4_destruct_r;
  MyDTBool_Bool_Bool_t gacB_4_destruct_d;
  logic gacB_4_destruct_r;
  MyBool_t \v'acC_4_destruct_d ;
  logic \v'acC_4_destruct_r ;
  Pointer_QTree_Bool_t q1acF_3_destruct_d;
  logic q1acF_3_destruct_r;
  Pointer_QTree_Bool_t es_4_destruct_d;
  logic es_4_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  MyDTBool_Bool_t isZacA_3_destruct_d;
  logic isZacA_3_destruct_r;
  MyDTBool_Bool_Bool_t gacB_3_destruct_d;
  logic gacB_3_destruct_r;
  MyBool_t \v'acC_3_destruct_d ;
  logic \v'acC_3_destruct_r ;
  Pointer_QTree_Bool_t q1acF_2_destruct_d;
  logic q1acF_2_destruct_r;
  Pointer_QTree_Bool_t q2acG_2_destruct_d;
  logic q2acG_2_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  MyDTBool_Bool_t isZacA_2_destruct_d;
  logic isZacA_2_destruct_r;
  MyDTBool_Bool_Bool_t gacB_2_destruct_d;
  logic gacB_2_destruct_r;
  MyBool_t \v'acC_2_destruct_d ;
  logic \v'acC_2_destruct_r ;
  Pointer_QTree_Bool_t q1acF_1_destruct_d;
  logic q1acF_1_destruct_r;
  Pointer_QTree_Bool_t q2acG_1_destruct_d;
  logic q2acG_1_destruct_r;
  Pointer_QTree_Bool_t q3acH_1_destruct_d;
  logic q3acH_1_destruct_r;
  \CTmap''_map''_Bool_Bool_Bool_t  _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_r ;
  Go_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d ;
  logic \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_r ;
  QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_goConst_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goConst_r ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_d ;
  logic \map''_map''_Bool_Bool_Bool_resbuf_r ;
  Pointer_MaskQTree_t q1ack_destruct_d;
  logic q1ack_destruct_r;
  Pointer_MaskQTree_t q2acl_destruct_d;
  logic q2acl_destruct_r;
  Pointer_MaskQTree_t q3acm_destruct_d;
  logic q3acm_destruct_r;
  Pointer_MaskQTree_t q4acn_destruct_d;
  logic q4acn_destruct_r;
  MaskQTree_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  MaskQTree_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  MaskQTree_t lizzieLet4_1MQNode_d;
  logic lizzieLet4_1MQNode_r;
  Go_t lizzieLet4_3MQNone_d;
  logic lizzieLet4_3MQNone_r;
  Go_t lizzieLet4_3MQVal_d;
  logic lizzieLet4_3MQVal_r;
  Go_t lizzieLet4_3MQNode_d;
  logic lizzieLet4_3MQNode_r;
  Go_t lizzieLet4_3MQNone_1_d;
  logic lizzieLet4_3MQNone_1_r;
  Go_t lizzieLet4_3MQNone_2_d;
  logic lizzieLet4_3MQNone_2_r;
  QTree_Bool_t lizzieLet4_3MQNone_1QNone_Bool_d;
  logic lizzieLet4_3MQNone_1QNone_Bool_r;
  QTree_Bool_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Go_t lizzieLet4_3MQNone_2_argbuf_d;
  logic lizzieLet4_3MQNone_2_argbuf_r;
  C6_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t lizzieLet4_3MQVal_1_argbuf_d;
  logic lizzieLet4_3MQVal_1_argbuf_r;
  QTree_Bool_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  QTree_Bool_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  QTree_Bool_t lizzieLet4_4MQNode_d;
  logic lizzieLet4_4MQNode_r;
  QTree_Bool_t lizzieLet4_4MQNode_1_d;
  logic lizzieLet4_4MQNode_1_r;
  QTree_Bool_t lizzieLet4_4MQNode_2_d;
  logic lizzieLet4_4MQNode_2_r;
  QTree_Bool_t lizzieLet4_4MQNode_3_d;
  logic lizzieLet4_4MQNode_3_r;
  QTree_Bool_t lizzieLet4_4MQNode_4_d;
  logic lizzieLet4_4MQNode_4_r;
  QTree_Bool_t lizzieLet4_4MQNode_5_d;
  logic lizzieLet4_4MQNode_5_r;
  QTree_Bool_t lizzieLet4_4MQNode_6_d;
  logic lizzieLet4_4MQNode_6_r;
  QTree_Bool_t lizzieLet4_4MQNode_7_d;
  logic lizzieLet4_4MQNode_7_r;
  QTree_Bool_t lizzieLet4_4MQNode_8_d;
  logic lizzieLet4_4MQNode_8_r;
  Pointer_QTree_Bool_t t1acp_destruct_d;
  logic t1acp_destruct_r;
  Pointer_QTree_Bool_t t2acq_destruct_d;
  logic t2acq_destruct_r;
  Pointer_QTree_Bool_t t3acr_destruct_d;
  logic t3acr_destruct_r;
  Pointer_QTree_Bool_t t4acs_destruct_d;
  logic t4acs_destruct_r;
  QTree_Bool_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  QTree_Bool_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  QTree_Bool_t lizzieLet4_4MQNode_1QNode_Bool_d;
  logic lizzieLet4_4MQNode_1QNode_Bool_r;
  QTree_Bool_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  Go_t lizzieLet4_4MQNode_3QNone_Bool_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_r;
  Go_t lizzieLet4_4MQNode_3QVal_Bool_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_r;
  Go_t lizzieLet4_4MQNode_3QNode_Bool_d;
  logic lizzieLet4_4MQNode_3QNode_Bool_r;
  Go_t lizzieLet4_4MQNode_3QError_Bool_d;
  logic lizzieLet4_4MQNode_3QError_Bool_r;
  Go_t lizzieLet4_4MQNode_3QError_Bool_1_d;
  logic lizzieLet4_4MQNode_3QError_Bool_1_r;
  Go_t lizzieLet4_4MQNode_3QError_Bool_2_d;
  logic lizzieLet4_4MQNode_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_d;
  logic lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QError_Bool_2_argbuf_d;
  logic lizzieLet4_4MQNode_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_d;
  logic lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QNone_Bool_1_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_1_r;
  Go_t lizzieLet4_4MQNode_3QNone_Bool_2_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_2_r;
  QTree_Bool_t lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QVal_Bool_1_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_1_r;
  Go_t lizzieLet4_4MQNode_3QVal_Bool_2_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Go_t lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNone_Bool_d;
  logic lizzieLet4_4MQNode_4QNone_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QVal_Bool_d;
  logic lizzieLet4_4MQNode_4QVal_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNode_Bool_d;
  logic lizzieLet4_4MQNode_4QNode_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QError_Bool_d;
  logic lizzieLet4_4MQNode_4QError_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QError_Bool_1_argbuf_d;
  logic lizzieLet4_4MQNode_4QError_Bool_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d;
  logic lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r;
  CTmain_mask_Bool_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_d;
  logic lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_d;
  logic lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Pointer_MaskQTree_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_5QNode_Bool_d;
  logic lizzieLet4_4MQNode_5QNode_Bool_r;
  Pointer_MaskQTree_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Pointer_MaskQTree_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  Pointer_MaskQTree_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_6QNode_Bool_d;
  logic lizzieLet4_4MQNode_6QNode_Bool_r;
  Pointer_MaskQTree_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_MaskQTree_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Pointer_MaskQTree_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_7QNode_Bool_d;
  logic lizzieLet4_4MQNode_7QNode_Bool_r;
  Pointer_MaskQTree_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_MaskQTree_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_MaskQTree_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_8QNode_Bool_d;
  logic lizzieLet4_4MQNode_8QNode_Bool_r;
  Pointer_MaskQTree_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_d;
  logic lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet4_5MQVal_d;
  logic lizzieLet4_5MQVal_r;
  Pointer_QTree_Bool_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet4_5MQVal_1_argbuf_d;
  logic lizzieLet4_5MQVal_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQNone_d;
  logic lizzieLet4_6MQNone_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQVal_d;
  logic lizzieLet4_6MQVal_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQNode_d;
  logic lizzieLet4_6MQNode_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQNone_1_argbuf_d;
  logic lizzieLet4_6MQNone_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQVal_1_argbuf_d;
  logic lizzieLet4_6MQVal_1_argbuf_r;
  Pointer_QTree_Bool_t m1acL_1_argbuf_d;
  logic m1acL_1_argbuf_r;
  Pointer_QTree_Bool_t m2acM_2_2_argbuf_d;
  logic m2acM_2_2_argbuf_r;
  Pointer_QTree_Bool_t m2acM_2_1_d;
  logic m2acM_2_1_r;
  Pointer_QTree_Bool_t m2acM_2_2_d;
  logic m2acM_2_2_r;
  Pointer_QTree_Bool_t m2acM_3_2_argbuf_d;
  logic m2acM_3_2_argbuf_r;
  Pointer_QTree_Bool_t m2acM_3_1_d;
  logic m2acM_3_1_r;
  Pointer_QTree_Bool_t m2acM_3_2_d;
  logic m2acM_3_2_r;
  Pointer_QTree_Bool_t m2acM_4_1_argbuf_d;
  logic m2acM_4_1_argbuf_r;
  Pointer_QTree_Bool_t macD_1_argbuf_d;
  logic macD_1_argbuf_r;
  Pointer_QTree_Bool_t maci_1_argbuf_d;
  logic maci_1_argbuf_r;
  Pointer_QTree_Bool_t maci_1_d;
  logic maci_1_r;
  Pointer_QTree_Bool_t maci_2_d;
  logic maci_2_r;
  Go_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_r;
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_r;
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_r;
  Go_t go_8_1_d;
  logic go_8_1_r;
  Go_t go_8_2_d;
  logic go_8_2_r;
  Pointer_QTree_Bool_t maci_1_1_argbuf_d;
  logic maci_1_1_argbuf_r;
  Pointer_MaskQTree_t mskacj_1_1_argbuf_d;
  logic mskacj_1_1_argbuf_r;
  Go_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_r ;
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_r ;
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_r ;
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_r ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_r ;
  MyDTBool_Bool_Bool_t gacB_1_1_argbuf_d;
  logic gacB_1_1_argbuf_r;
  Go_t go_9_1_d;
  logic go_9_1_r;
  Go_t go_9_2_d;
  logic go_9_2_r;
  MyDTBool_Bool_t isZacA_1_1_argbuf_d;
  logic isZacA_1_1_argbuf_r;
  Pointer_QTree_Bool_t macD_1_1_argbuf_d;
  logic macD_1_1_argbuf_r;
  MyBool_t \v'acC_1_1_argbuf_d ;
  logic \v'acC_1_1_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_MaskQTree_t mskacj_1_argbuf_d;
  logic mskacj_1_argbuf_r;
  Pointer_QTree_Bool_t q1acF_3_1_argbuf_d;
  logic q1acF_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1acO_3_1_argbuf_d;
  logic q1acO_3_1_argbuf_r;
  Pointer_MaskQTree_t q1ack_3_1_argbuf_d;
  logic q1ack_3_1_argbuf_r;
  Pointer_QTree_Bool_t q2acG_2_1_argbuf_d;
  logic q2acG_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2acP_2_1_argbuf_d;
  logic q2acP_2_1_argbuf_r;
  Pointer_MaskQTree_t q2acl_2_1_argbuf_d;
  logic q2acl_2_1_argbuf_r;
  Pointer_QTree_Bool_t q3acH_1_1_argbuf_d;
  logic q3acH_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3acQ_1_1_argbuf_d;
  logic q3acQ_1_1_argbuf_r;
  Pointer_MaskQTree_t q3acm_1_1_argbuf_d;
  logic q3acm_1_1_argbuf_r;
  Pointer_QTree_Bool_t q4acI_1_argbuf_d;
  logic q4acI_1_argbuf_r;
  Pointer_QTree_Bool_t q4acR_1_argbuf_d;
  logic q4acR_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_1_d;
  logic lizzieLet20_1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_2_d;
  logic lizzieLet20_2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_3_d;
  logic lizzieLet20_3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4_d;
  logic lizzieLet20_4_r;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r;
  CTmain_mask_Bool_t lizzieLet25_1_d;
  logic lizzieLet25_1_r;
  CTmain_mask_Bool_t lizzieLet25_2_d;
  logic lizzieLet25_2_r;
  CTmain_mask_Bool_t lizzieLet25_3_d;
  logic lizzieLet25_3_r;
  CTmain_mask_Bool_t lizzieLet25_4_d;
  logic lizzieLet25_4_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet30_1_d;
  logic lizzieLet30_1_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet30_2_d;
  logic lizzieLet30_2_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet30_3_d;
  logic lizzieLet30_3_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet30_4_d;
  logic lizzieLet30_4_r;
  MaskQTree_t readPointer_MaskQTreemskacj_1_argbuf_rwb_d;
  logic readPointer_MaskQTreemskacj_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  MaskQTree_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  MaskQTree_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  MaskQTree_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  MaskQTree_t lizzieLet4_5_d;
  logic lizzieLet4_5_r;
  MaskQTree_t lizzieLet4_6_d;
  logic lizzieLet4_6_r;
  QTree_Bool_t readPointer_QTree_Boolm1acL_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm1acL_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet0_1_d;
  logic lizzieLet0_1_r;
  QTree_Bool_t lizzieLet0_2_d;
  logic lizzieLet0_2_r;
  QTree_Bool_t lizzieLet0_3_d;
  logic lizzieLet0_3_r;
  QTree_Bool_t lizzieLet0_4_d;
  logic lizzieLet0_4_r;
  QTree_Bool_t lizzieLet0_5_d;
  logic lizzieLet0_5_r;
  QTree_Bool_t lizzieLet0_6_d;
  logic lizzieLet0_6_r;
  QTree_Bool_t lizzieLet0_7_d;
  logic lizzieLet0_7_r;
  QTree_Bool_t readPointer_QTree_BoolmacD_1_argbuf_rwb_d;
  logic readPointer_QTree_BoolmacD_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet11_1_1_d;
  logic lizzieLet11_1_1_r;
  QTree_Bool_t lizzieLet11_1_2_d;
  logic lizzieLet11_1_2_r;
  QTree_Bool_t lizzieLet11_1_3_d;
  logic lizzieLet11_1_3_r;
  QTree_Bool_t lizzieLet11_1_4_d;
  logic lizzieLet11_1_4_r;
  QTree_Bool_t lizzieLet11_1_5_d;
  logic lizzieLet11_1_5_r;
  QTree_Bool_t lizzieLet11_1_6_d;
  logic lizzieLet11_1_6_r;
  QTree_Bool_t lizzieLet11_1_7_d;
  logic lizzieLet11_1_7_r;
  QTree_Bool_t readPointer_QTree_Boolmaci_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolmaci_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Bool_t t1acp_3_1_argbuf_d;
  logic t1acp_3_1_argbuf_r;
  Pointer_QTree_Bool_t t2acq_2_1_argbuf_d;
  logic t2acq_2_1_argbuf_r;
  Pointer_QTree_Bool_t t3acr_1_1_argbuf_d;
  logic t3acr_1_1_argbuf_r;
  Pointer_QTree_Bool_t t4acs_1_argbuf_d;
  logic t4acs_1_argbuf_r;
  MyBool_t \v'acC_2_2_argbuf_d ;
  logic \v'acC_2_2_argbuf_r ;
  MyBool_t \v'acC_2_1_d ;
  logic \v'acC_2_1_r ;
  MyBool_t \v'acC_2_2_d ;
  logic \v'acC_2_2_r ;
  MyBool_t \v'acC_3_2_argbuf_d ;
  logic \v'acC_3_2_argbuf_r ;
  MyBool_t \v'acC_3_1_d ;
  logic \v'acC_3_1_r ;
  MyBool_t \v'acC_3_2_d ;
  logic \v'acC_3_2_r ;
  MyBool_t \v'acC_4_1_argbuf_d ;
  logic \v'acC_4_1_argbuf_r ;
  MyBool_t vacE_1_argbuf_d;
  logic vacE_1_argbuf_r;
  MyBool_t vacN_1_argbuf_d;
  logic vacN_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet13_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet16_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet8_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  MyBool_t xabY_1_argbuf_d;
  logic xabY_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go)] */
  logic [9:0] sourceGo_emitted;
  logic [9:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign sourceGo_done = (sourceGo_emitted | ({go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 10'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 10'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Bool,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0,
                                go_1_dummy_write_QTree_Bool_d[0]};
  assign go_1_dummy_write_QTree_Bool_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Bool,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go_2_dummy_write_QTree_Bool_d[0])
          incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go_2_dummy_write_QTree_Bool_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go_2_dummy_write_QTree_Bool_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                                            2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Bool_snk,Word16#) > */
  assign {forkHP1_QTree_Bool_snk_r,
          forkHP1_QTree_Bool_snk_dout} = {forkHP1_QTree_Bool_snk_rout,
                                          forkHP1_QTree_Bool_snk_d};
  
  /* source (Ty Go) : > (\QTree_Bool_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Bool_src,Go) > [(go_1_dummy_write_QTree_Bool,Go),
                                       (go_2_dummy_write_QTree_Bool,Go)] */
  logic [1:0] \\QTree_Bool_src_emitted ;
  logic [1:0] \\QTree_Bool_src_done ;
  assign go_1_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [0]));
  assign go_2_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [1]));
  assign \\QTree_Bool_src_done  = (\\QTree_Bool_src_emitted  | ({go_2_dummy_write_QTree_Bool_d[0],
                                                                 go_1_dummy_write_QTree_Bool_d[0]} & {go_2_dummy_write_QTree_Bool_r,
                                                                                                      go_1_dummy_write_QTree_Bool_r}));
  assign \\QTree_Bool_src_r  = (& \\QTree_Bool_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Bool_src_emitted  <= 2'd0;
    else
      \\QTree_Bool_src_emitted  <= (\\QTree_Bool_src_r  ? 2'd0 :
                                    \\QTree_Bool_src_done );
  
  /* source (Ty QTree_Bool) : > (dummy_write_QTree_Bool,QTree_Bool) */
  
  /* sink (Ty Pointer_QTree_Bool) : (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool) > */
  assign {dummy_write_QTree_Bool_sink_r,
          dummy_write_QTree_Bool_sink_dout} = {dummy_write_QTree_Bool_sink_rout,
                                               dummy_write_QTree_Bool_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Bool_snk,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#),
                                                        (forkHP1_QTree_Boo4,Word16#)] */
  logic [3:0] mergeHP_QTree_Bool_buf_emitted;
  logic [3:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Bool_snk_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                     (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign forkHP1_QTree_Boo4_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[3]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo4_d[0],
                                                                           forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Bool_snk_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo4_r,
                                                                                                       forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Bool_snk_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 4'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Bool) : [(m1acL_1_argbuf,Pointer_QTree_Bool),
                                     (macD_1_argbuf,Pointer_QTree_Bool),
                                     (maci_1_argbuf,Pointer_QTree_Bool)] > (readMerge_choice_QTree_Bool,C3) (readMerge_data_QTree_Bool,Pointer_QTree_Bool) */
  logic [2:0] m1acL_1_argbuf_select_d;
  assign m1acL_1_argbuf_select_d = ((| m1acL_1_argbuf_select_q) ? m1acL_1_argbuf_select_q :
                                    (m1acL_1_argbuf_d[0] ? 3'd1 :
                                     (macD_1_argbuf_d[0] ? 3'd2 :
                                      (maci_1_argbuf_d[0] ? 3'd4 :
                                       3'd0))));
  logic [2:0] m1acL_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acL_1_argbuf_select_q <= 3'd0;
    else
      m1acL_1_argbuf_select_q <= (m1acL_1_argbuf_done ? 3'd0 :
                                  m1acL_1_argbuf_select_d);
  logic [1:0] m1acL_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acL_1_argbuf_emit_q <= 2'd0;
    else
      m1acL_1_argbuf_emit_q <= (m1acL_1_argbuf_done ? 2'd0 :
                                m1acL_1_argbuf_emit_d);
  logic [1:0] m1acL_1_argbuf_emit_d;
  assign m1acL_1_argbuf_emit_d = (m1acL_1_argbuf_emit_q | ({readMerge_choice_QTree_Bool_d[0],
                                                            readMerge_data_QTree_Bool_d[0]} & {readMerge_choice_QTree_Bool_r,
                                                                                               readMerge_data_QTree_Bool_r}));
  logic m1acL_1_argbuf_done;
  assign m1acL_1_argbuf_done = (& m1acL_1_argbuf_emit_d);
  assign {maci_1_argbuf_r,
          macD_1_argbuf_r,
          m1acL_1_argbuf_r} = (m1acL_1_argbuf_done ? m1acL_1_argbuf_select_d :
                               3'd0);
  assign readMerge_data_QTree_Bool_d = ((m1acL_1_argbuf_select_d[0] && (! m1acL_1_argbuf_emit_q[0])) ? m1acL_1_argbuf_d :
                                        ((m1acL_1_argbuf_select_d[1] && (! m1acL_1_argbuf_emit_q[0])) ? macD_1_argbuf_d :
                                         ((m1acL_1_argbuf_select_d[2] && (! m1acL_1_argbuf_emit_q[0])) ? maci_1_argbuf_d :
                                          {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Bool_d = ((m1acL_1_argbuf_select_d[0] && (! m1acL_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((m1acL_1_argbuf_select_d[1] && (! m1acL_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((m1acL_1_argbuf_select_d[2] && (! m1acL_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Bool) : (readMerge_choice_QTree_Bool,C3) (destructReadOut_QTree_Bool,QTree_Bool) > [(readPointer_QTree_Boolm1acL_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_BoolmacD_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolmaci_1_argbuf,QTree_Bool)] */
  logic [2:0] destructReadOut_QTree_Bool_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Bool_d[0] && destructReadOut_QTree_Bool_d[0]))
      unique case (readMerge_choice_QTree_Bool_d[2:1])
        2'd0: destructReadOut_QTree_Bool_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Bool_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Bool_onehotd = 3'd4;
        default: destructReadOut_QTree_Bool_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Bool_onehotd = 3'd0;
  assign readPointer_QTree_Boolm1acL_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[0]};
  assign readPointer_QTree_BoolmacD_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                  destructReadOut_QTree_Bool_onehotd[1]};
  assign readPointer_QTree_Boolmaci_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                  destructReadOut_QTree_Bool_onehotd[2]};
  assign destructReadOut_QTree_Bool_r = (| (destructReadOut_QTree_Bool_onehotd & {readPointer_QTree_Boolmaci_1_argbuf_r,
                                                                                  readPointer_QTree_BoolmacD_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm1acL_1_argbuf_r}));
  assign readMerge_choice_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (readMerge_data_QTree_Bool,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {readMerge_data_QTree_Bool_d[16:1],
                                        readMerge_data_QTree_Bool_d[0]};
  assign readMerge_data_QTree_Bool_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(destructReadOut_QTree_Bool,QTree_Bool)] */
  assign destructReadOut_QTree_Bool_d = {memReadOut_QTree_Bool_d[67:2],
                                         memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* mergectrl (Ty C14,
           Ty QTree_Bool) : [(lizzieLet10_1_1_argbuf,QTree_Bool),
                             (lizzieLet12_1_1_argbuf,QTree_Bool),
                             (lizzieLet13_1_argbuf,QTree_Bool),
                             (lizzieLet14_1_argbuf,QTree_Bool),
                             (lizzieLet16_1_argbuf,QTree_Bool),
                             (lizzieLet1_1_argbuf,QTree_Bool),
                             (lizzieLet24_1_argbuf,QTree_Bool),
                             (lizzieLet29_1_argbuf,QTree_Bool),
                             (lizzieLet34_1_argbuf,QTree_Bool),
                             (lizzieLet3_1_argbuf,QTree_Bool),
                             (lizzieLet5_1_argbuf,QTree_Bool),
                             (lizzieLet7_1_argbuf,QTree_Bool),
                             (lizzieLet8_1_argbuf,QTree_Bool),
                             (dummy_write_QTree_Bool,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C14) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [13:0] lizzieLet10_1_1_argbuf_select_d;
  assign lizzieLet10_1_1_argbuf_select_d = ((| lizzieLet10_1_1_argbuf_select_q) ? lizzieLet10_1_1_argbuf_select_q :
                                            (lizzieLet10_1_1_argbuf_d[0] ? 14'd1 :
                                             (lizzieLet12_1_1_argbuf_d[0] ? 14'd2 :
                                              (lizzieLet13_1_argbuf_d[0] ? 14'd4 :
                                               (lizzieLet14_1_argbuf_d[0] ? 14'd8 :
                                                (lizzieLet16_1_argbuf_d[0] ? 14'd16 :
                                                 (lizzieLet1_1_argbuf_d[0] ? 14'd32 :
                                                  (lizzieLet24_1_argbuf_d[0] ? 14'd64 :
                                                   (lizzieLet29_1_argbuf_d[0] ? 14'd128 :
                                                    (lizzieLet34_1_argbuf_d[0] ? 14'd256 :
                                                     (lizzieLet3_1_argbuf_d[0] ? 14'd512 :
                                                      (lizzieLet5_1_argbuf_d[0] ? 14'd1024 :
                                                       (lizzieLet7_1_argbuf_d[0] ? 14'd2048 :
                                                        (lizzieLet8_1_argbuf_d[0] ? 14'd4096 :
                                                         (dummy_write_QTree_Bool_d[0] ? 14'd8192 :
                                                          14'd0)))))))))))))));
  logic [13:0] lizzieLet10_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_select_q <= 14'd0;
    else
      lizzieLet10_1_1_argbuf_select_q <= (lizzieLet10_1_1_argbuf_done ? 14'd0 :
                                          lizzieLet10_1_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_1_argbuf_emit_q <= (lizzieLet10_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet10_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_d;
  assign lizzieLet10_1_1_argbuf_emit_d = (lizzieLet10_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                            writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                                writeMerge_data_QTree_Bool_r}));
  logic lizzieLet10_1_1_argbuf_done;
  assign lizzieLet10_1_1_argbuf_done = (& lizzieLet10_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Bool_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet3_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet1_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet13_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = (lizzieLet10_1_1_argbuf_done ? lizzieLet10_1_1_argbuf_select_d :
                                       14'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet10_1_1_argbuf_d :
                                         ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet12_1_1_argbuf_d :
                                          ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_argbuf_d :
                                           ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                            ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                             ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet1_1_argbuf_d :
                                              ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                               ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                                ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                 ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet3_1_argbuf_d :
                                                  ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                                   ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                    ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                                     ((lizzieLet10_1_1_argbuf_select_d[13] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Bool_d :
                                                      {66'd0, 1'd0}))))))))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C1_14_dc(1'd1) :
                                           ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C2_14_dc(1'd1) :
                                            ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C3_14_dc(1'd1) :
                                             ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C4_14_dc(1'd1) :
                                              ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C5_14_dc(1'd1) :
                                               ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C6_14_dc(1'd1) :
                                                ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C7_14_dc(1'd1) :
                                                 ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C8_14_dc(1'd1) :
                                                  ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C9_14_dc(1'd1) :
                                                   ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C10_14_dc(1'd1) :
                                                    ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C11_14_dc(1'd1) :
                                                     ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C12_14_dc(1'd1) :
                                                      ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C13_14_dc(1'd1) :
                                                       ((lizzieLet10_1_1_argbuf_select_d[13] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C14_14_dc(1'd1) :
                                                        {4'd0, 1'd0}))))))))))))));
  
  /* demux (Ty C14,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C14) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet12_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet13_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet16_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet24_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet29_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet8_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool)] */
  logic [13:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[4:1])
        4'd0: demuxWriteResult_QTree_Bool_onehotd = 14'd1;
        4'd1: demuxWriteResult_QTree_Bool_onehotd = 14'd2;
        4'd2: demuxWriteResult_QTree_Bool_onehotd = 14'd4;
        4'd3: demuxWriteResult_QTree_Bool_onehotd = 14'd8;
        4'd4: demuxWriteResult_QTree_Bool_onehotd = 14'd16;
        4'd5: demuxWriteResult_QTree_Bool_onehotd = 14'd32;
        4'd6: demuxWriteResult_QTree_Bool_onehotd = 14'd64;
        4'd7: demuxWriteResult_QTree_Bool_onehotd = 14'd128;
        4'd8: demuxWriteResult_QTree_Bool_onehotd = 14'd256;
        4'd9: demuxWriteResult_QTree_Bool_onehotd = 14'd512;
        4'd10: demuxWriteResult_QTree_Bool_onehotd = 14'd1024;
        4'd11: demuxWriteResult_QTree_Bool_onehotd = 14'd2048;
        4'd12: demuxWriteResult_QTree_Bool_onehotd = 14'd4096;
        4'd13: demuxWriteResult_QTree_Bool_onehotd = 14'd8192;
        default: demuxWriteResult_QTree_Bool_onehotd = 14'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 14'd0;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet12_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet13_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet16_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet24_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet29_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[7]};
  assign writeQTree_BoollizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[8]};
  assign writeQTree_BoollizzieLet3_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[9]};
  assign writeQTree_BoollizzieLet5_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[10]};
  assign writeQTree_BoollizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[11]};
  assign writeQTree_BoollizzieLet8_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[12]};
  assign dummy_write_QTree_Bool_sink_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                          demuxWriteResult_QTree_Bool_onehotd[13]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {dummy_write_QTree_Bool_sink_r,
                                                                                    writeQTree_BoollizzieLet8_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet7_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet5_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet3_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet34_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet29_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet24_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet16_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet14_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet13_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet12_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet10_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo3_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo3_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo4,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo4_d[0]}), forkHP1_QTree_Boo4_d);
  assign {forkHP1_QTree_Boo4_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_50,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _50_d = {dconPtr_QTree_Bool_d[16:1],
                  dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _50_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__5,Go) > (initHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \initHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd0,
                                                    go__5_d[0]};
  assign go__5_r = \initHP_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmap''_map''_Bool_Bool_Bool1,Go) > (incrHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd1,
                                                    \incrHP_CTmap''_map''_Bool_Bool_Bool1_d [0]};
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool1_r  = \incrHP_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* merge (Ty Go) : [(go__6,Go),
                 (incrHP_CTmap''_map''_Bool_Bool_Bool2,Go)] > (incrHP_mergeCTmap''_map''_Bool_Bool_Bool,Go) */
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ;
  always_comb
    begin
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  = 2'd0;
      if ((| \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  = \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ;
      else
        if (go__6_d[0])
          \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [0] = 1'd1;
        else if (\incrHP_CTmap''_map''_Bool_Bool_Bool2_d [0])
          \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select  <= (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  ? 2'd0 :
                                                            \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected );
  always_comb
    if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [0])
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = go__6_d;
    else if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [1])
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = \incrHP_CTmap''_map''_Bool_Bool_Bool2_d ;
    else \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = 1'd0;
  assign {\incrHP_CTmap''_map''_Bool_Bool_Bool2_r ,
          go__6_r} = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  ? \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf,Go) > [(incrHP_CTmap''_map''_Bool_Bool_Bool1,Go),
                                                                    (incrHP_CTmap''_map''_Bool_Bool_Bool2,Go)] */
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done ;
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool1_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted [0]));
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool2_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted [1]));
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  | ({\incrHP_CTmap''_map''_Bool_Bool_Bool2_d [0],
                                                                                                                           \incrHP_CTmap''_map''_Bool_Bool_Bool1_d [0]} & {\incrHP_CTmap''_map''_Bool_Bool_Bool2_r ,
                                                                                                                                                                           \incrHP_CTmap''_map''_Bool_Bool_Bool1_r }));
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  = (& \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  <= (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  ? 2'd0 :
                                                                 \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmap''_map''_Bool_Bool_Bool,Word16#) (forkHP1_CTmap''_map''_Bool_Bool_Bool,Word16#) > (addHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \addHP_CTmap''_map''_Bool_Bool_Bool_d  = {(\incrHP_CTmap''_map''_Bool_Bool_Bool_d [16:1] + \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [16:1]),
                                                   (\incrHP_CTmap''_map''_Bool_Bool_Bool_d [0] && \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [0])};
  assign {\incrHP_CTmap''_map''_Bool_Bool_Bool_r ,
          \forkHP1_CTmap''_map''_Bool_Bool_Bool_r } = {2 {(\addHP_CTmap''_map''_Bool_Bool_Bool_r  && \addHP_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmap''_map''_Bool_Bool_Bool,Word16#),
                      (addHP_CTmap''_map''_Bool_Bool_Bool,Word16#)] > (mergeHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  logic [1:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected ;
  logic [1:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ;
  always_comb
    begin
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  = 2'd0;
      if ((| \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  = \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ;
      else
        if (\initHP_CTmap''_map''_Bool_Bool_Bool_d [0])
          \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [0] = 1'd1;
        else if (\addHP_CTmap''_map''_Bool_Bool_Bool_d [0])
          \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_select  <= 2'd0;
    else
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_select  <= (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r  ? 2'd0 :
                                                        \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected );
  always_comb
    if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [0])
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = \initHP_CTmap''_map''_Bool_Bool_Bool_d ;
    else if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [1])
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = \addHP_CTmap''_map''_Bool_Bool_Bool_d ;
    else \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd0, 1'd0};
  assign {\addHP_CTmap''_map''_Bool_Bool_Bool_r ,
          \initHP_CTmap''_map''_Bool_Bool_Bool_r } = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r  ? \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  :
                                                      2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmap''_map''_Bool_Bool_Bool,Go) > (incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf,Go) */
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r ;
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  = ((! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d [0]) || \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r )
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d  <= \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf ;
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r  = (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]);
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0] ? \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  :
                                                             \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  && \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r ) && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0])))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmap''_map''_Bool_Bool_Bool,Word16#) > (mergeHP_CTmap''_map''_Bool_Bool_Bool_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r ;
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_r  = ((! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d [0]) || \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r )
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d  <= \mergeHP_CTmap''_map''_Bool_Bool_Bool_d ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf ;
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r  = (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]);
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d  = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0] ? \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  :
                                                         \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  && \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r ) && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0])))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmap''_map''_Bool_Bool_Bool_buf,Word16#) > [(forkHP1_CTmap''_map''_Bool_Bool_Bool,Word16#),
                                                                          (forkHP1_CTmap''_map''_Bool_Bool_Boo2,Word16#),
                                                                          (forkHP1_CTmap''_map''_Bool_Bool_Boo3,Word16#)] */
  logic [2:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted ;
  logic [2:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done ;
  assign \forkHP1_CTmap''_map''_Bool_Bool_Bool_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [0]))};
  assign \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [1]))};
  assign \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [2]))};
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done  = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  | ({\forkHP1_CTmap''_map''_Bool_Bool_Boo3_d [0],
                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d [0],
                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_r ,
                                                                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ,
                                                                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Bool_r }));
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  = (& \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  <= (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  ? 3'd0 :
                                                             \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : [(dconReadIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool),
                                                     (dconWriteIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool)] > (memMergeChoice_CTmap''_map''_Bool_Bool_Bool,C2) (memMergeIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d  = ((| \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q ) ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  :
                                                               (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_d [0] ? 2'd1 :
                                                                (\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d [0] ? 2'd2 :
                                                                 2'd0)));
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  <= (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? 2'd0 :
                                                             \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  <= (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? 2'd0 :
                                                           \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d  = (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  | ({\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [0],
                                                                                                                  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                                                                     \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r }));
  logic \dconReadIn_CTmap''_map''_Bool_Bool_Bool_done ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  = (& \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d );
  assign {\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r ,
          \dconReadIn_CTmap''_map''_Bool_Bool_Bool_r } = (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d  :
                                                          2'd0);
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d  = ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [0] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [0])) ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d  :
                                                        ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [1] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [0])) ? \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d  :
                                                         {85'd0, 1'd0}));
  assign \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d  = ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [0] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [1])) ? C1_2_dc(1'd1) :
                                                            ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [1] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [1])) ? C2_2_dc(1'd1) :
                                                             {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  logic [67:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ;
  logic [67:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
  logic [67:0] \memOut_CTmap''_map''_Bool_Bool_Bool_q ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_valid ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_we ;
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din  = \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [85:18];
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address  = \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [17:2];
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we  = (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [1:1] && \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmap''_map''_Bool_Bool_Bool_we  <= 1'd0;
        \memOut_CTmap''_map''_Bool_Bool_Bool_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmap''_map''_Bool_Bool_Bool_we  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we ;
        \memOut_CTmap''_map''_Bool_Bool_Bool_valid  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0];
        if (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we )
          begin
            \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ] <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
            \memOut_CTmap''_map''_Bool_Bool_Bool_q  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
          end
        else
          \memOut_CTmap''_map''_Bool_Bool_Bool_q  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ];
      end
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_q ,
                                                    \memOut_CTmap''_map''_Bool_Bool_Bool_we ,
                                                    \memOut_CTmap''_map''_Bool_Bool_Bool_valid };
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r  = ((! \memOut_CTmap''_map''_Bool_Bool_Bool_valid ) || \memOut_CTmap''_map''_Bool_Bool_Bool_r );
  logic [31:0] \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read ;
  logic [31:0] \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  <= 0;
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  <= 0;
      end
    else
      if ((\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we  == 1'd1))
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  <= (\profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  + 1);
      else
        if ((\memOut_CTmap''_map''_Bool_Bool_Bool_valid  == 1'd1))
          \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  <= (\profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memMergeChoice_CTmap''_map''_Bool_Bool_Bool,C2) (memOut_CTmap''_map''_Bool_Bool_Bool_dbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) > [(memReadOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                    (memWriteOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [0] && \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]))
      unique case (\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [1:1])
        1'd0: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [69:1],
                                                        \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd [0]};
  assign \memWriteOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [69:1],
                                                         \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd [1]};
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r  = (| (\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  & {\memWriteOut_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                  \memReadOut_CTmap''_map''_Bool_Bool_Bool_r }));
  assign \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r  = \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r  = ((! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]) || \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= {85'd0, 1'd0};
    else
      if (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r )
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf ;
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r  = (! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0]);
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d  = (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0] ? \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  :
                                                             \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= {85'd0, 1'd0};
    else
      if ((\memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r  && \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0]))
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= {85'd0, 1'd0};
      else if (((! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r ) && (! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0])))
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d ;
  
  /* dbuf (Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memOut_CTmap''_map''_Bool_Bool_Bool_rbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool_dbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r  = ((! \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]) || \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= {69'd0, 1'd0};
    else
      if (\memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r )
        \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool_rbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_buf ;
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_r  = (! \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0]);
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d  = (\memOut_CTmap''_map''_Bool_Bool_Bool_buf [0] ? \memOut_CTmap''_map''_Bool_Bool_Bool_buf  :
                                                         \memOut_CTmap''_map''_Bool_Bool_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= {69'd0, 1'd0};
    else
      if ((\memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r  && \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0]))
        \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= {69'd0, 1'd0};
      else if (((! \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r ) && (! \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0])))
        \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= \memOut_CTmap''_map''_Bool_Bool_Bool_d ;
  
  /* destruct (Ty Pointer_CTmap''_map''_Bool_Bool_Bool,
          Dcon Pointer_CTmap''_map''_Bool_Bool_Bool) : (scfarg_0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(destructReadIn_CTmap''_map''_Bool_Bool_Bool,Word16#)] */
  assign \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                                            scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Dcon ReadIn_CTmap''_map''_Bool_Bool_Bool) : [(destructReadIn_CTmap''_map''_Bool_Bool_Bool,Word16#)] > (dconReadIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d  = \ReadIn_CTmap''_map''_Bool_Bool_Bool_dc ((& {\destructReadIn_CTmap''_map''_Bool_Bool_Bool_d [0]}), \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d );
  assign {\destructReadIn_CTmap''_map''_Bool_Bool_Bool_r } = {1 {(\dconReadIn_CTmap''_map''_Bool_Bool_Bool_r  && \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* destruct (Ty MemOut_CTmap''_map''_Bool_Bool_Bool,
          Dcon ReadOut_CTmap''_map''_Bool_Bool_Bool) : (memReadOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) > [(readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf,CTmap''_map''_Bool_Bool_Bool)] */
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d  = {\memReadOut_CTmap''_map''_Bool_Bool_Bool_d [69:2],
                                                                            \memReadOut_CTmap''_map''_Bool_Bool_Bool_d [0]};
  assign \memReadOut_CTmap''_map''_Bool_Bool_Bool_r  = \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmap''_map''_Bool_Bool_Bool) : [(lizzieLet15_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet19_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet31_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet32_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet33_1_argbuf,CTmap''_map''_Bool_Bool_Bool)] > (writeMerge_choice_CTmap''_map''_Bool_Bool_Bool,C5) (writeMerge_data_CTmap''_map''_Bool_Bool_Bool,CTmap''_map''_Bool_Bool_Bool) */
  logic [4:0] lizzieLet15_1_argbuf_select_d;
  assign lizzieLet15_1_argbuf_select_d = ((| lizzieLet15_1_argbuf_select_q) ? lizzieLet15_1_argbuf_select_q :
                                          (lizzieLet15_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet19_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet31_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet32_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet33_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet15_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet15_1_argbuf_select_q <= (lizzieLet15_1_argbuf_done ? 5'd0 :
                                        lizzieLet15_1_argbuf_select_d);
  logic [1:0] lizzieLet15_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet15_1_argbuf_emit_q <= (lizzieLet15_1_argbuf_done ? 2'd0 :
                                      lizzieLet15_1_argbuf_emit_d);
  logic [1:0] lizzieLet15_1_argbuf_emit_d;
  assign lizzieLet15_1_argbuf_emit_d = (lizzieLet15_1_argbuf_emit_q | ({\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [0],
                                                                        \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                                \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r }));
  logic lizzieLet15_1_argbuf_done;
  assign lizzieLet15_1_argbuf_done = (& lizzieLet15_1_argbuf_emit_d);
  assign {lizzieLet33_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet15_1_argbuf_r} = (lizzieLet15_1_argbuf_done ? lizzieLet15_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d  = ((lizzieLet15_1_argbuf_select_d[0] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                                             ((lizzieLet15_1_argbuf_select_d[1] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                                              ((lizzieLet15_1_argbuf_select_d[2] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                               ((lizzieLet15_1_argbuf_select_d[3] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                                ((lizzieLet15_1_argbuf_select_d[4] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                                 {68'd0, 1'd0})))));
  assign \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d  = ((lizzieLet15_1_argbuf_select_d[0] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                               ((lizzieLet15_1_argbuf_select_d[1] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                                ((lizzieLet15_1_argbuf_select_d[2] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                 ((lizzieLet15_1_argbuf_select_d[3] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                  ((lizzieLet15_1_argbuf_select_d[4] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                   {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeMerge_choice_CTmap''_map''_Bool_Bool_Bool,C5) (demuxWriteResult_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [4:0] \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [0] && \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [0]))
      unique case (\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [3:1])
        3'd0:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd0;
      endcase
    else
      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd0;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [0]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [1]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [2]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [3]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [4]};
  assign \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r  = (| (\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  & {\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_r }));
  assign \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r  = \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Dcon WriteIn_CTmap''_map''_Bool_Bool_Bool) : [(forkHP1_CTmap''_map''_Bool_Bool_Boo2,Word16#),
                                                    (writeMerge_data_CTmap''_map''_Bool_Bool_Bool,CTmap''_map''_Bool_Bool_Bool)] > (dconWriteIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d  = \WriteIn_CTmap''_map''_Bool_Bool_Bool_dc ((& {\forkHP1_CTmap''_map''_Bool_Bool_Boo2_d [0],
                                                                                                      \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d [0]}), \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d , \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d );
  assign {\forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ,
          \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r } = {2 {(\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r  && \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* dcon (Ty Pointer_CTmap''_map''_Bool_Bool_Bool,
      Dcon Pointer_CTmap''_map''_Bool_Bool_Bool) : [(forkHP1_CTmap''_map''_Bool_Bool_Boo3,Word16#)] > (dconPtr_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconPtr_CTmap''_map''_Bool_Bool_Bool_d  = \Pointer_CTmap''_map''_Bool_Bool_Bool_dc ((& {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_d [0]}), \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d );
  assign {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_r } = {1 {(\dconPtr_CTmap''_map''_Bool_Bool_Bool_r  && \dconPtr_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* demux (Ty MemOut_CTmap''_map''_Bool_Bool_Bool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (memWriteOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) (dconPtr_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(_49,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                                                (demuxWriteResult_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd ;
  always_comb
    if ((\memWriteOut_CTmap''_map''_Bool_Bool_Bool_d [0] && \dconPtr_CTmap''_map''_Bool_Bool_Bool_d [0]))
      unique case (\memWriteOut_CTmap''_map''_Bool_Bool_Bool_d [1:1])
        1'd0: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd2;
        default: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd0;
  assign _49_d = {\dconPtr_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                  \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd [0]};
  assign \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d  = {\dconPtr_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                              \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd [1]};
  assign \dconPtr_CTmap''_map''_Bool_Bool_Bool_r  = (| (\dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  & {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                          _49_r}));
  assign \memWriteOut_CTmap''_map''_Bool_Bool_Bool_r  = \dconPtr_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go__7,Go) > (initHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign initHP_CTkron_kron_Bool_Bool_Bool_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_CTkron_kron_Bool_Bool_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTkron_kron_Bool_Bool_Bool1,Go) > (incrHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign incrHP_CTkron_kron_Bool_Bool_Bool_d = {16'd1,
                                                incrHP_CTkron_kron_Bool_Bool_Bool1_d[0]};
  assign incrHP_CTkron_kron_Bool_Bool_Bool1_r = incrHP_CTkron_kron_Bool_Bool_Bool_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CTkron_kron_Bool_Bool_Bool2,Go)] > (incrHP_mergeCTkron_kron_Bool_Bool_Bool,Go) */
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected;
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_select;
  always_comb
    begin
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected = 2'd0;
      if ((| incrHP_mergeCTkron_kron_Bool_Bool_Bool_select))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected = incrHP_mergeCTkron_kron_Bool_Bool_Bool_select;
      else
        if (go__8_d[0])
          incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[0] = 1'd1;
        else if (incrHP_CTkron_kron_Bool_Bool_Bool2_d[0])
          incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_select <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_select <= (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r ? 2'd0 :
                                                        incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected);
  always_comb
    if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[0])
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = go__8_d;
    else if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[1])
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = incrHP_CTkron_kron_Bool_Bool_Bool2_d;
    else incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = 1'd0;
  assign {incrHP_CTkron_kron_Bool_Bool_Bool2_r,
          go__8_r} = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r ? incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf,Go) > [(incrHP_CTkron_kron_Bool_Bool_Bool1,Go),
                                                                  (incrHP_CTkron_kron_Bool_Bool_Bool2,Go)] */
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted;
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done;
  assign incrHP_CTkron_kron_Bool_Bool_Bool1_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d[0] && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted[0]));
  assign incrHP_CTkron_kron_Bool_Bool_Bool2_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d[0] && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted[1]));
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted | ({incrHP_CTkron_kron_Bool_Bool_Bool2_d[0],
                                                                                                                   incrHP_CTkron_kron_Bool_Bool_Bool1_d[0]} & {incrHP_CTkron_kron_Bool_Bool_Bool2_r,
                                                                                                                                                               incrHP_CTkron_kron_Bool_Bool_Bool1_r}));
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r = (& incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted <= (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r ? 2'd0 :
                                                             incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTkron_kron_Bool_Bool_Bool,Word16#) (forkHP1_CTkron_kron_Bool_Bool_Bool,Word16#) > (addHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign addHP_CTkron_kron_Bool_Bool_Bool_d = {(incrHP_CTkron_kron_Bool_Bool_Bool_d[16:1] + forkHP1_CTkron_kron_Bool_Bool_Bool_d[16:1]),
                                               (incrHP_CTkron_kron_Bool_Bool_Bool_d[0] && forkHP1_CTkron_kron_Bool_Bool_Bool_d[0])};
  assign {incrHP_CTkron_kron_Bool_Bool_Bool_r,
          forkHP1_CTkron_kron_Bool_Bool_Bool_r} = {2 {(addHP_CTkron_kron_Bool_Bool_Bool_r && addHP_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTkron_kron_Bool_Bool_Bool,Word16#),
                      (addHP_CTkron_kron_Bool_Bool_Bool,Word16#)] > (mergeHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  logic [1:0] mergeHP_CTkron_kron_Bool_Bool_Bool_selected;
  logic [1:0] mergeHP_CTkron_kron_Bool_Bool_Bool_select;
  always_comb
    begin
      mergeHP_CTkron_kron_Bool_Bool_Bool_selected = 2'd0;
      if ((| mergeHP_CTkron_kron_Bool_Bool_Bool_select))
        mergeHP_CTkron_kron_Bool_Bool_Bool_selected = mergeHP_CTkron_kron_Bool_Bool_Bool_select;
      else
        if (initHP_CTkron_kron_Bool_Bool_Bool_d[0])
          mergeHP_CTkron_kron_Bool_Bool_Bool_selected[0] = 1'd1;
        else if (addHP_CTkron_kron_Bool_Bool_Bool_d[0])
          mergeHP_CTkron_kron_Bool_Bool_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_select <= 2'd0;
    else
      mergeHP_CTkron_kron_Bool_Bool_Bool_select <= (mergeHP_CTkron_kron_Bool_Bool_Bool_r ? 2'd0 :
                                                    mergeHP_CTkron_kron_Bool_Bool_Bool_selected);
  always_comb
    if (mergeHP_CTkron_kron_Bool_Bool_Bool_selected[0])
      mergeHP_CTkron_kron_Bool_Bool_Bool_d = initHP_CTkron_kron_Bool_Bool_Bool_d;
    else if (mergeHP_CTkron_kron_Bool_Bool_Bool_selected[1])
      mergeHP_CTkron_kron_Bool_Bool_Bool_d = addHP_CTkron_kron_Bool_Bool_Bool_d;
    else mergeHP_CTkron_kron_Bool_Bool_Bool_d = {16'd0, 1'd0};
  assign {addHP_CTkron_kron_Bool_Bool_Bool_r,
          initHP_CTkron_kron_Bool_Bool_Bool_r} = (mergeHP_CTkron_kron_Bool_Bool_Bool_r ? mergeHP_CTkron_kron_Bool_Bool_Bool_selected :
                                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTkron_kron_Bool_Bool_Bool,Go) > (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf,Go) */
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r;
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_r = ((! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d[0]) || incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r)
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d <= incrHP_mergeCTkron_kron_Bool_Bool_Bool_d;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf;
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r = (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0]);
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0] ? incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf :
                                                         incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r && incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0]))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r) && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0])))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTkron_kron_Bool_Bool_Bool,Word16#) > (mergeHP_CTkron_kron_Bool_Bool_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r;
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_r = ((! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d[0]) || mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTkron_kron_Bool_Bool_Bool_r)
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d <= mergeHP_CTkron_kron_Bool_Bool_Bool_d;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf;
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r = (! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0]);
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d = (mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0] ? mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf :
                                                     mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r && mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0]))
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r) && (! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0])))
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTkron_kron_Bool_Bool_Bool_buf,Word16#) > [(forkHP1_CTkron_kron_Bool_Bool_Bool,Word16#),
                                                                        (forkHP1_CTkron_kron_Bool_Bool_Boo2,Word16#),
                                                                        (forkHP1_CTkron_kron_Bool_Bool_Boo3,Word16#)] */
  logic [2:0] mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted;
  logic [2:0] mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done;
  assign forkHP1_CTkron_kron_Bool_Bool_Bool_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[0]))};
  assign forkHP1_CTkron_kron_Bool_Bool_Boo2_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[1]))};
  assign forkHP1_CTkron_kron_Bool_Bool_Boo3_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[2]))};
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done = (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted | ({forkHP1_CTkron_kron_Bool_Bool_Boo3_d[0],
                                                                                                           forkHP1_CTkron_kron_Bool_Bool_Boo2_d[0],
                                                                                                           forkHP1_CTkron_kron_Bool_Bool_Bool_d[0]} & {forkHP1_CTkron_kron_Bool_Bool_Boo3_r,
                                                                                                                                                       forkHP1_CTkron_kron_Bool_Bool_Boo2_r,
                                                                                                                                                       forkHP1_CTkron_kron_Bool_Bool_Bool_r}));
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r = (& mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted <= (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r ? 3'd0 :
                                                         mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTkron_kron_Bool_Bool_Bool) : [(dconReadIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool),
                                                   (dconWriteIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool)] > (memMergeChoice_CTkron_kron_Bool_Bool_Bool,C2) (memMergeIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d = ((| dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q) ? dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q :
                                                           (dconReadIn_CTkron_kron_Bool_Bool_Bool_d[0] ? 2'd1 :
                                                            (dconWriteIn_CTkron_kron_Bool_Bool_Bool_d[0] ? 2'd2 :
                                                             2'd0)));
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q <= (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? 2'd0 :
                                                         dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d);
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q <= (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? 2'd0 :
                                                       dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d);
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d = (dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q | ({memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[0],
                                                                                                          memMergeIn_CTkron_kron_Bool_Bool_Bool_d[0]} & {memMergeChoice_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                                                                         memMergeIn_CTkron_kron_Bool_Bool_Bool_r}));
  logic dconReadIn_CTkron_kron_Bool_Bool_Bool_done;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_done = (& dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d);
  assign {dconWriteIn_CTkron_kron_Bool_Bool_Bool_r,
          dconReadIn_CTkron_kron_Bool_Bool_Bool_r} = (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d :
                                                      2'd0);
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_d = ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[0] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[0])) ? dconReadIn_CTkron_kron_Bool_Bool_Bool_d :
                                                    ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[1] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[0])) ? dconWriteIn_CTkron_kron_Bool_Bool_Bool_d :
                                                     {100'd0, 1'd0}));
  assign memMergeChoice_CTkron_kron_Bool_Bool_Bool_d = ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[0] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                                        ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[1] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf,MemIn_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) */
  logic [82:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address;
  logic [82:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
  logic [82:0] memOut_CTkron_kron_Bool_Bool_Bool_q;
  logic memOut_CTkron_kron_Bool_Bool_Bool_valid;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we;
  logic memOut_CTkron_kron_Bool_Bool_Bool_we;
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din = memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[100:18];
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address = memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[17:2];
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we = (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[1:1] && memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTkron_kron_Bool_Bool_Bool_we <= 1'd0;
        memOut_CTkron_kron_Bool_Bool_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_CTkron_kron_Bool_Bool_Bool_we <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we;
        memOut_CTkron_kron_Bool_Bool_Bool_valid <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0];
        if (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we)
          begin
            memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address] <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
            memOut_CTkron_kron_Bool_Bool_Bool_q <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
          end
        else
          memOut_CTkron_kron_Bool_Bool_Bool_q <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address];
      end
  assign memOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_q,
                                                memOut_CTkron_kron_Bool_Bool_Bool_we,
                                                memOut_CTkron_kron_Bool_Bool_Bool_valid};
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r = ((! memOut_CTkron_kron_Bool_Bool_Bool_valid) || memOut_CTkron_kron_Bool_Bool_Bool_r);
  logic [31:0] profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read;
  logic [31:0] profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write <= 0;
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read <= 0;
      end
    else
      if ((memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we == 1'd1))
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write <= (profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write + 1);
      else
        if ((memOut_CTkron_kron_Bool_Bool_Bool_valid == 1'd1))
          profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read <= (profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memMergeChoice_CTkron_kron_Bool_Bool_Bool,C2) (memOut_CTkron_kron_Bool_Bool_Bool_dbuf,MemOut_CTkron_kron_Bool_Bool_Bool) > [(memReadOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                            (memWriteOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool)] */
  logic [1:0] memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[0] && memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]))
      unique case (memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[1:1])
        1'd0: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd2;
        default: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[84:1],
                                                    memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd[0]};
  assign memWriteOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[84:1],
                                                     memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd[1]};
  assign memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r = (| (memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd & {memWriteOut_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                          memReadOut_CTkron_kron_Bool_Bool_Bool_r}));
  assign memMergeChoice_CTkron_kron_Bool_Bool_Bool_r = memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf,MemIn_CTkron_kron_Bool_Bool_Bool) > (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r = ((! memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]) || memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d <= {100'd0, 1'd0};
    else
      if (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r)
        memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d <= memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) > (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf,MemIn_CTkron_kron_Bool_Bool_Bool) */
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_buf;
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_r = (! memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0]);
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d = (memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0] ? memMergeIn_CTkron_kron_Bool_Bool_Bool_buf :
                                                         memMergeIn_CTkron_kron_Bool_Bool_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= {100'd0, 1'd0};
    else
      if ((memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r && memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0]))
        memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= {100'd0, 1'd0};
      else if (((! memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r) && (! memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0])))
        memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= memMergeIn_CTkron_kron_Bool_Bool_Bool_d;
  
  /* dbuf (Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memOut_CTkron_kron_Bool_Bool_Bool_rbuf,MemOut_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool_dbuf,MemOut_CTkron_kron_Bool_Bool_Bool) */
  assign memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r = ((! memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]) || memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d <= {84'd0, 1'd0};
    else
      if (memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r)
        memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d <= memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool_rbuf,MemOut_CTkron_kron_Bool_Bool_Bool) */
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_buf;
  assign memOut_CTkron_kron_Bool_Bool_Bool_r = (! memOut_CTkron_kron_Bool_Bool_Bool_buf[0]);
  assign memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d = (memOut_CTkron_kron_Bool_Bool_Bool_buf[0] ? memOut_CTkron_kron_Bool_Bool_Bool_buf :
                                                     memOut_CTkron_kron_Bool_Bool_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Bool_Bool_Bool_buf <= {84'd0, 1'd0};
    else
      if ((memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r && memOut_CTkron_kron_Bool_Bool_Bool_buf[0]))
        memOut_CTkron_kron_Bool_Bool_Bool_buf <= {84'd0, 1'd0};
      else if (((! memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r) && (! memOut_CTkron_kron_Bool_Bool_Bool_buf[0])))
        memOut_CTkron_kron_Bool_Bool_Bool_buf <= memOut_CTkron_kron_Bool_Bool_Bool_d;
  
  /* destruct (Ty Pointer_CTkron_kron_Bool_Bool_Bool,
          Dcon Pointer_CTkron_kron_Bool_Bool_Bool) : (scfarg_0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > [(destructReadIn_CTkron_kron_Bool_Bool_Bool,Word16#)] */
  assign destructReadIn_CTkron_kron_Bool_Bool_Bool_d = {scfarg_0_1_argbuf_d[16:1],
                                                        scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CTkron_kron_Bool_Bool_Bool_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Dcon ReadIn_CTkron_kron_Bool_Bool_Bool) : [(destructReadIn_CTkron_kron_Bool_Bool_Bool,Word16#)] > (dconReadIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_d = ReadIn_CTkron_kron_Bool_Bool_Bool_dc((& {destructReadIn_CTkron_kron_Bool_Bool_Bool_d[0]}), destructReadIn_CTkron_kron_Bool_Bool_Bool_d);
  assign {destructReadIn_CTkron_kron_Bool_Bool_Bool_r} = {1 {(dconReadIn_CTkron_kron_Bool_Bool_Bool_r && dconReadIn_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* destruct (Ty MemOut_CTkron_kron_Bool_Bool_Bool,
          Dcon ReadOut_CTkron_kron_Bool_Bool_Bool) : (memReadOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) > [(readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf,CTkron_kron_Bool_Bool_Bool)] */
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d = {memReadOut_CTkron_kron_Bool_Bool_Bool_d[84:2],
                                                                      memReadOut_CTkron_kron_Bool_Bool_Bool_d[0]};
  assign memReadOut_CTkron_kron_Bool_Bool_Bool_r = readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTkron_kron_Bool_Bool_Bool) : [(lizzieLet17_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet21_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet22_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet23_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet2_1_argbuf,CTkron_kron_Bool_Bool_Bool)] > (writeMerge_choice_CTkron_kron_Bool_Bool_Bool,C5) (writeMerge_data_CTkron_kron_Bool_Bool_Bool,CTkron_kron_Bool_Bool_Bool) */
  logic [4:0] lizzieLet17_1_argbuf_select_d;
  assign lizzieLet17_1_argbuf_select_d = ((| lizzieLet17_1_argbuf_select_q) ? lizzieLet17_1_argbuf_select_q :
                                          (lizzieLet17_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet21_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet22_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet23_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet2_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet17_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet17_1_argbuf_select_q <= (lizzieLet17_1_argbuf_done ? 5'd0 :
                                        lizzieLet17_1_argbuf_select_d);
  logic [1:0] lizzieLet17_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet17_1_argbuf_emit_q <= (lizzieLet17_1_argbuf_done ? 2'd0 :
                                      lizzieLet17_1_argbuf_emit_d);
  logic [1:0] lizzieLet17_1_argbuf_emit_d;
  assign lizzieLet17_1_argbuf_emit_d = (lizzieLet17_1_argbuf_emit_q | ({writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[0],
                                                                        writeMerge_data_CTkron_kron_Bool_Bool_Bool_d[0]} & {writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                                            writeMerge_data_CTkron_kron_Bool_Bool_Bool_r}));
  logic lizzieLet17_1_argbuf_done;
  assign lizzieLet17_1_argbuf_done = (& lizzieLet17_1_argbuf_emit_d);
  assign {lizzieLet2_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet17_1_argbuf_r} = (lizzieLet17_1_argbuf_done ? lizzieLet17_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTkron_kron_Bool_Bool_Bool_d = ((lizzieLet17_1_argbuf_select_d[0] && (! lizzieLet17_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                                         ((lizzieLet17_1_argbuf_select_d[1] && (! lizzieLet17_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                                          ((lizzieLet17_1_argbuf_select_d[2] && (! lizzieLet17_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                                           ((lizzieLet17_1_argbuf_select_d[3] && (! lizzieLet17_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                            ((lizzieLet17_1_argbuf_select_d[4] && (! lizzieLet17_1_argbuf_emit_q[0])) ? lizzieLet2_1_argbuf_d :
                                                             {83'd0, 1'd0})))));
  assign writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d = ((lizzieLet17_1_argbuf_select_d[0] && (! lizzieLet17_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                           ((lizzieLet17_1_argbuf_select_d[1] && (! lizzieLet17_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                            ((lizzieLet17_1_argbuf_select_d[2] && (! lizzieLet17_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                             ((lizzieLet17_1_argbuf_select_d[3] && (! lizzieLet17_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                              ((lizzieLet17_1_argbuf_select_d[4] && (! lizzieLet17_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                               {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeMerge_choice_CTkron_kron_Bool_Bool_Bool,C5) (demuxWriteResult_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > [(writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [4:0] demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[0] && demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[0]))
      unique case (writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[3:1])
        3'd0: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd16;
        default:
          demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd0;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[0]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[1]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[2]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[3]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                 demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[4]};
  assign demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r = (| (demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd & {writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_r}));
  assign writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r = demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Dcon WriteIn_CTkron_kron_Bool_Bool_Bool) : [(forkHP1_CTkron_kron_Bool_Bool_Boo2,Word16#),
                                                  (writeMerge_data_CTkron_kron_Bool_Bool_Bool,CTkron_kron_Bool_Bool_Bool)] > (dconWriteIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign dconWriteIn_CTkron_kron_Bool_Bool_Bool_d = WriteIn_CTkron_kron_Bool_Bool_Bool_dc((& {forkHP1_CTkron_kron_Bool_Bool_Boo2_d[0],
                                                                                              writeMerge_data_CTkron_kron_Bool_Bool_Bool_d[0]}), forkHP1_CTkron_kron_Bool_Bool_Boo2_d, writeMerge_data_CTkron_kron_Bool_Bool_Bool_d);
  assign {forkHP1_CTkron_kron_Bool_Bool_Boo2_r,
          writeMerge_data_CTkron_kron_Bool_Bool_Bool_r} = {2 {(dconWriteIn_CTkron_kron_Bool_Bool_Bool_r && dconWriteIn_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* dcon (Ty Pointer_CTkron_kron_Bool_Bool_Bool,
      Dcon Pointer_CTkron_kron_Bool_Bool_Bool) : [(forkHP1_CTkron_kron_Bool_Bool_Boo3,Word16#)] > (dconPtr_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign dconPtr_CTkron_kron_Bool_Bool_Bool_d = Pointer_CTkron_kron_Bool_Bool_Bool_dc((& {forkHP1_CTkron_kron_Bool_Bool_Boo3_d[0]}), forkHP1_CTkron_kron_Bool_Bool_Boo3_d);
  assign {forkHP1_CTkron_kron_Bool_Bool_Boo3_r} = {1 {(dconPtr_CTkron_kron_Bool_Bool_Bool_r && dconPtr_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* demux (Ty MemOut_CTkron_kron_Bool_Bool_Bool,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (memWriteOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) (dconPtr_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > [(_48,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                                      (demuxWriteResult_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [1:0] dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd;
  always_comb
    if ((memWriteOut_CTkron_kron_Bool_Bool_Bool_d[0] && dconPtr_CTkron_kron_Bool_Bool_Bool_d[0]))
      unique case (memWriteOut_CTkron_kron_Bool_Bool_Bool_d[1:1])
        1'd0: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd1;
        1'd1: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd2;
        default: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd0;
  assign _48_d = {dconPtr_CTkron_kron_Bool_Bool_Bool_d[16:1],
                  dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd[0]};
  assign demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d = {dconPtr_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                          dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd[1]};
  assign dconPtr_CTkron_kron_Bool_Bool_Bool_r = (| (dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd & {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                  _48_r}));
  assign memWriteOut_CTkron_kron_Bool_Bool_Bool_r = dconPtr_CTkron_kron_Bool_Bool_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTmain_mask_Bool,Word16#) */
  assign initHP_CTmain_mask_Bool_d = {16'd0, go__9_d[0]};
  assign go__9_r = initHP_CTmain_mask_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_mask_Bool1,Go) > (incrHP_CTmain_mask_Bool,Word16#) */
  assign incrHP_CTmain_mask_Bool_d = {16'd1,
                                      incrHP_CTmain_mask_Bool1_d[0]};
  assign incrHP_CTmain_mask_Bool1_r = incrHP_CTmain_mask_Bool_r;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTmain_mask_Bool2,Go)] > (incrHP_mergeCTmain_mask_Bool,Go) */
  logic [1:0] incrHP_mergeCTmain_mask_Bool_selected;
  logic [1:0] incrHP_mergeCTmain_mask_Bool_select;
  always_comb
    begin
      incrHP_mergeCTmain_mask_Bool_selected = 2'd0;
      if ((| incrHP_mergeCTmain_mask_Bool_select))
        incrHP_mergeCTmain_mask_Bool_selected = incrHP_mergeCTmain_mask_Bool_select;
      else
        if (go__10_d[0]) incrHP_mergeCTmain_mask_Bool_selected[0] = 1'd1;
        else if (incrHP_CTmain_mask_Bool2_d[0])
          incrHP_mergeCTmain_mask_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Bool_select <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Bool_select <= (incrHP_mergeCTmain_mask_Bool_r ? 2'd0 :
                                              incrHP_mergeCTmain_mask_Bool_selected);
  always_comb
    if (incrHP_mergeCTmain_mask_Bool_selected[0])
      incrHP_mergeCTmain_mask_Bool_d = go__10_d;
    else if (incrHP_mergeCTmain_mask_Bool_selected[1])
      incrHP_mergeCTmain_mask_Bool_d = incrHP_CTmain_mask_Bool2_d;
    else incrHP_mergeCTmain_mask_Bool_d = 1'd0;
  assign {incrHP_CTmain_mask_Bool2_r,
          go__10_r} = (incrHP_mergeCTmain_mask_Bool_r ? incrHP_mergeCTmain_mask_Bool_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_mask_Bool_buf,Go) > [(incrHP_CTmain_mask_Bool1,Go),
                                                        (incrHP_CTmain_mask_Bool2,Go)] */
  logic [1:0] incrHP_mergeCTmain_mask_Bool_buf_emitted;
  logic [1:0] incrHP_mergeCTmain_mask_Bool_buf_done;
  assign incrHP_CTmain_mask_Bool1_d = (incrHP_mergeCTmain_mask_Bool_buf_d[0] && (! incrHP_mergeCTmain_mask_Bool_buf_emitted[0]));
  assign incrHP_CTmain_mask_Bool2_d = (incrHP_mergeCTmain_mask_Bool_buf_d[0] && (! incrHP_mergeCTmain_mask_Bool_buf_emitted[1]));
  assign incrHP_mergeCTmain_mask_Bool_buf_done = (incrHP_mergeCTmain_mask_Bool_buf_emitted | ({incrHP_CTmain_mask_Bool2_d[0],
                                                                                               incrHP_CTmain_mask_Bool1_d[0]} & {incrHP_CTmain_mask_Bool2_r,
                                                                                                                                 incrHP_CTmain_mask_Bool1_r}));
  assign incrHP_mergeCTmain_mask_Bool_buf_r = (& incrHP_mergeCTmain_mask_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Bool_buf_emitted <= (incrHP_mergeCTmain_mask_Bool_buf_r ? 2'd0 :
                                                   incrHP_mergeCTmain_mask_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_mask_Bool,Word16#) (forkHP1_CTmain_mask_Bool,Word16#) > (addHP_CTmain_mask_Bool,Word16#) */
  assign addHP_CTmain_mask_Bool_d = {(incrHP_CTmain_mask_Bool_d[16:1] + forkHP1_CTmain_mask_Bool_d[16:1]),
                                     (incrHP_CTmain_mask_Bool_d[0] && forkHP1_CTmain_mask_Bool_d[0])};
  assign {incrHP_CTmain_mask_Bool_r,
          forkHP1_CTmain_mask_Bool_r} = {2 {(addHP_CTmain_mask_Bool_r && addHP_CTmain_mask_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_mask_Bool,Word16#),
                      (addHP_CTmain_mask_Bool,Word16#)] > (mergeHP_CTmain_mask_Bool,Word16#) */
  logic [1:0] mergeHP_CTmain_mask_Bool_selected;
  logic [1:0] mergeHP_CTmain_mask_Bool_select;
  always_comb
    begin
      mergeHP_CTmain_mask_Bool_selected = 2'd0;
      if ((| mergeHP_CTmain_mask_Bool_select))
        mergeHP_CTmain_mask_Bool_selected = mergeHP_CTmain_mask_Bool_select;
      else
        if (initHP_CTmain_mask_Bool_d[0])
          mergeHP_CTmain_mask_Bool_selected[0] = 1'd1;
        else if (addHP_CTmain_mask_Bool_d[0])
          mergeHP_CTmain_mask_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Bool_select <= 2'd0;
    else
      mergeHP_CTmain_mask_Bool_select <= (mergeHP_CTmain_mask_Bool_r ? 2'd0 :
                                          mergeHP_CTmain_mask_Bool_selected);
  always_comb
    if (mergeHP_CTmain_mask_Bool_selected[0])
      mergeHP_CTmain_mask_Bool_d = initHP_CTmain_mask_Bool_d;
    else if (mergeHP_CTmain_mask_Bool_selected[1])
      mergeHP_CTmain_mask_Bool_d = addHP_CTmain_mask_Bool_d;
    else mergeHP_CTmain_mask_Bool_d = {16'd0, 1'd0};
  assign {addHP_CTmain_mask_Bool_r,
          initHP_CTmain_mask_Bool_r} = (mergeHP_CTmain_mask_Bool_r ? mergeHP_CTmain_mask_Bool_selected :
                                        2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_mask_Bool,Go) > (incrHP_mergeCTmain_mask_Bool_buf,Go) */
  Go_t incrHP_mergeCTmain_mask_Bool_bufchan_d;
  logic incrHP_mergeCTmain_mask_Bool_bufchan_r;
  assign incrHP_mergeCTmain_mask_Bool_r = ((! incrHP_mergeCTmain_mask_Bool_bufchan_d[0]) || incrHP_mergeCTmain_mask_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTmain_mask_Bool_r)
        incrHP_mergeCTmain_mask_Bool_bufchan_d <= incrHP_mergeCTmain_mask_Bool_d;
  Go_t incrHP_mergeCTmain_mask_Bool_bufchan_buf;
  assign incrHP_mergeCTmain_mask_Bool_bufchan_r = (! incrHP_mergeCTmain_mask_Bool_bufchan_buf[0]);
  assign incrHP_mergeCTmain_mask_Bool_buf_d = (incrHP_mergeCTmain_mask_Bool_bufchan_buf[0] ? incrHP_mergeCTmain_mask_Bool_bufchan_buf :
                                               incrHP_mergeCTmain_mask_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTmain_mask_Bool_buf_r && incrHP_mergeCTmain_mask_Bool_bufchan_buf[0]))
        incrHP_mergeCTmain_mask_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTmain_mask_Bool_buf_r) && (! incrHP_mergeCTmain_mask_Bool_bufchan_buf[0])))
        incrHP_mergeCTmain_mask_Bool_bufchan_buf <= incrHP_mergeCTmain_mask_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_mask_Bool,Word16#) > (mergeHP_CTmain_mask_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_CTmain_mask_Bool_bufchan_d;
  logic mergeHP_CTmain_mask_Bool_bufchan_r;
  assign mergeHP_CTmain_mask_Bool_r = ((! mergeHP_CTmain_mask_Bool_bufchan_d[0]) || mergeHP_CTmain_mask_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTmain_mask_Bool_r)
        mergeHP_CTmain_mask_Bool_bufchan_d <= mergeHP_CTmain_mask_Bool_d;
  \Word16#_t  mergeHP_CTmain_mask_Bool_bufchan_buf;
  assign mergeHP_CTmain_mask_Bool_bufchan_r = (! mergeHP_CTmain_mask_Bool_bufchan_buf[0]);
  assign mergeHP_CTmain_mask_Bool_buf_d = (mergeHP_CTmain_mask_Bool_bufchan_buf[0] ? mergeHP_CTmain_mask_Bool_bufchan_buf :
                                           mergeHP_CTmain_mask_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTmain_mask_Bool_buf_r && mergeHP_CTmain_mask_Bool_bufchan_buf[0]))
        mergeHP_CTmain_mask_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTmain_mask_Bool_buf_r) && (! mergeHP_CTmain_mask_Bool_bufchan_buf[0])))
        mergeHP_CTmain_mask_Bool_bufchan_buf <= mergeHP_CTmain_mask_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_mask_Bool_buf,Word16#) > [(forkHP1_CTmain_mask_Bool,Word16#),
                                                              (forkHP1_CTmain_mask_Boo2,Word16#),
                                                              (forkHP1_CTmain_mask_Boo3,Word16#)] */
  logic [2:0] mergeHP_CTmain_mask_Bool_buf_emitted;
  logic [2:0] mergeHP_CTmain_mask_Bool_buf_done;
  assign forkHP1_CTmain_mask_Bool_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[0]))};
  assign forkHP1_CTmain_mask_Boo2_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[1]))};
  assign forkHP1_CTmain_mask_Boo3_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[2]))};
  assign mergeHP_CTmain_mask_Bool_buf_done = (mergeHP_CTmain_mask_Bool_buf_emitted | ({forkHP1_CTmain_mask_Boo3_d[0],
                                                                                       forkHP1_CTmain_mask_Boo2_d[0],
                                                                                       forkHP1_CTmain_mask_Bool_d[0]} & {forkHP1_CTmain_mask_Boo3_r,
                                                                                                                         forkHP1_CTmain_mask_Boo2_r,
                                                                                                                         forkHP1_CTmain_mask_Bool_r}));
  assign mergeHP_CTmain_mask_Bool_buf_r = (& mergeHP_CTmain_mask_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_CTmain_mask_Bool_buf_emitted <= (mergeHP_CTmain_mask_Bool_buf_r ? 3'd0 :
                                               mergeHP_CTmain_mask_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_mask_Bool) : [(dconReadIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool),
                                         (dconWriteIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool)] > (memMergeChoice_CTmain_mask_Bool,C2) (memMergeIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  logic [1:0] dconReadIn_CTmain_mask_Bool_select_d;
  assign dconReadIn_CTmain_mask_Bool_select_d = ((| dconReadIn_CTmain_mask_Bool_select_q) ? dconReadIn_CTmain_mask_Bool_select_q :
                                                 (dconReadIn_CTmain_mask_Bool_d[0] ? 2'd1 :
                                                  (dconWriteIn_CTmain_mask_Bool_d[0] ? 2'd2 :
                                                   2'd0)));
  logic [1:0] dconReadIn_CTmain_mask_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Bool_select_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Bool_select_q <= (dconReadIn_CTmain_mask_Bool_done ? 2'd0 :
                                               dconReadIn_CTmain_mask_Bool_select_d);
  logic [1:0] dconReadIn_CTmain_mask_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Bool_emit_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Bool_emit_q <= (dconReadIn_CTmain_mask_Bool_done ? 2'd0 :
                                             dconReadIn_CTmain_mask_Bool_emit_d);
  logic [1:0] dconReadIn_CTmain_mask_Bool_emit_d;
  assign dconReadIn_CTmain_mask_Bool_emit_d = (dconReadIn_CTmain_mask_Bool_emit_q | ({memMergeChoice_CTmain_mask_Bool_d[0],
                                                                                      memMergeIn_CTmain_mask_Bool_d[0]} & {memMergeChoice_CTmain_mask_Bool_r,
                                                                                                                           memMergeIn_CTmain_mask_Bool_r}));
  logic dconReadIn_CTmain_mask_Bool_done;
  assign dconReadIn_CTmain_mask_Bool_done = (& dconReadIn_CTmain_mask_Bool_emit_d);
  assign {dconWriteIn_CTmain_mask_Bool_r,
          dconReadIn_CTmain_mask_Bool_r} = (dconReadIn_CTmain_mask_Bool_done ? dconReadIn_CTmain_mask_Bool_select_d :
                                            2'd0);
  assign memMergeIn_CTmain_mask_Bool_d = ((dconReadIn_CTmain_mask_Bool_select_d[0] && (! dconReadIn_CTmain_mask_Bool_emit_q[0])) ? dconReadIn_CTmain_mask_Bool_d :
                                          ((dconReadIn_CTmain_mask_Bool_select_d[1] && (! dconReadIn_CTmain_mask_Bool_emit_q[0])) ? dconWriteIn_CTmain_mask_Bool_d :
                                           {132'd0, 1'd0}));
  assign memMergeChoice_CTmain_mask_Bool_d = ((dconReadIn_CTmain_mask_Bool_select_d[0] && (! dconReadIn_CTmain_mask_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                              ((dconReadIn_CTmain_mask_Bool_select_d[1] && (! dconReadIn_CTmain_mask_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                               {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_mask_Bool,
      Ty MemOut_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool_dbuf,MemIn_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) */
  logic [114:0] memMergeIn_CTmain_mask_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTmain_mask_Bool_dbuf_address;
  logic [114:0] memMergeIn_CTmain_mask_Bool_dbuf_din;
  logic [114:0] memOut_CTmain_mask_Bool_q;
  logic memOut_CTmain_mask_Bool_valid;
  logic memMergeIn_CTmain_mask_Bool_dbuf_we;
  logic memOut_CTmain_mask_Bool_we;
  assign memMergeIn_CTmain_mask_Bool_dbuf_din = memMergeIn_CTmain_mask_Bool_dbuf_d[132:18];
  assign memMergeIn_CTmain_mask_Bool_dbuf_address = memMergeIn_CTmain_mask_Bool_dbuf_d[17:2];
  assign memMergeIn_CTmain_mask_Bool_dbuf_we = (memMergeIn_CTmain_mask_Bool_dbuf_d[1:1] && memMergeIn_CTmain_mask_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTmain_mask_Bool_we <= 1'd0;
        memOut_CTmain_mask_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_CTmain_mask_Bool_we <= memMergeIn_CTmain_mask_Bool_dbuf_we;
        memOut_CTmain_mask_Bool_valid <= memMergeIn_CTmain_mask_Bool_dbuf_d[0];
        if (memMergeIn_CTmain_mask_Bool_dbuf_we)
          begin
            memMergeIn_CTmain_mask_Bool_dbuf_mem[memMergeIn_CTmain_mask_Bool_dbuf_address] <= memMergeIn_CTmain_mask_Bool_dbuf_din;
            memOut_CTmain_mask_Bool_q <= memMergeIn_CTmain_mask_Bool_dbuf_din;
          end
        else
          memOut_CTmain_mask_Bool_q <= memMergeIn_CTmain_mask_Bool_dbuf_mem[memMergeIn_CTmain_mask_Bool_dbuf_address];
      end
  assign memOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_q,
                                      memOut_CTmain_mask_Bool_we,
                                      memOut_CTmain_mask_Bool_valid};
  assign memMergeIn_CTmain_mask_Bool_dbuf_r = ((! memOut_CTmain_mask_Bool_valid) || memOut_CTmain_mask_Bool_r);
  logic [31:0] profiling_MemIn_CTmain_mask_Bool_read;
  logic [31:0] profiling_MemIn_CTmain_mask_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTmain_mask_Bool_write <= 0;
        profiling_MemIn_CTmain_mask_Bool_read <= 0;
      end
    else
      if ((memMergeIn_CTmain_mask_Bool_dbuf_we == 1'd1))
        profiling_MemIn_CTmain_mask_Bool_write <= (profiling_MemIn_CTmain_mask_Bool_write + 1);
      else
        if ((memOut_CTmain_mask_Bool_valid == 1'd1))
          profiling_MemIn_CTmain_mask_Bool_read <= (profiling_MemIn_CTmain_mask_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_mask_Bool) : (memMergeChoice_CTmain_mask_Bool,C2) (memOut_CTmain_mask_Bool_dbuf,MemOut_CTmain_mask_Bool) > [(memReadOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool),
                                                                                                                                    (memWriteOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool)] */
  logic [1:0] memOut_CTmain_mask_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTmain_mask_Bool_d[0] && memOut_CTmain_mask_Bool_dbuf_d[0]))
      unique case (memMergeChoice_CTmain_mask_Bool_d[1:1])
        1'd0: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd2;
        default: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_dbuf_d[116:1],
                                          memOut_CTmain_mask_Bool_dbuf_onehotd[0]};
  assign memWriteOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_dbuf_d[116:1],
                                           memOut_CTmain_mask_Bool_dbuf_onehotd[1]};
  assign memOut_CTmain_mask_Bool_dbuf_r = (| (memOut_CTmain_mask_Bool_dbuf_onehotd & {memWriteOut_CTmain_mask_Bool_r,
                                                                                      memReadOut_CTmain_mask_Bool_r}));
  assign memMergeChoice_CTmain_mask_Bool_r = memOut_CTmain_mask_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool_rbuf,MemIn_CTmain_mask_Bool) > (memMergeIn_CTmain_mask_Bool_dbuf,MemIn_CTmain_mask_Bool) */
  assign memMergeIn_CTmain_mask_Bool_rbuf_r = ((! memMergeIn_CTmain_mask_Bool_dbuf_d[0]) || memMergeIn_CTmain_mask_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Bool_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTmain_mask_Bool_rbuf_r)
        memMergeIn_CTmain_mask_Bool_dbuf_d <= memMergeIn_CTmain_mask_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) > (memMergeIn_CTmain_mask_Bool_rbuf,MemIn_CTmain_mask_Bool) */
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_buf;
  assign memMergeIn_CTmain_mask_Bool_r = (! memMergeIn_CTmain_mask_Bool_buf[0]);
  assign memMergeIn_CTmain_mask_Bool_rbuf_d = (memMergeIn_CTmain_mask_Bool_buf[0] ? memMergeIn_CTmain_mask_Bool_buf :
                                               memMergeIn_CTmain_mask_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Bool_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTmain_mask_Bool_rbuf_r && memMergeIn_CTmain_mask_Bool_buf[0]))
        memMergeIn_CTmain_mask_Bool_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTmain_mask_Bool_rbuf_r) && (! memMergeIn_CTmain_mask_Bool_buf[0])))
        memMergeIn_CTmain_mask_Bool_buf <= memMergeIn_CTmain_mask_Bool_d;
  
  /* dbuf (Ty MemOut_CTmain_mask_Bool) : (memOut_CTmain_mask_Bool_rbuf,MemOut_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool_dbuf,MemOut_CTmain_mask_Bool) */
  assign memOut_CTmain_mask_Bool_rbuf_r = ((! memOut_CTmain_mask_Bool_dbuf_d[0]) || memOut_CTmain_mask_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTmain_mask_Bool_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTmain_mask_Bool_rbuf_r)
        memOut_CTmain_mask_Bool_dbuf_d <= memOut_CTmain_mask_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_CTmain_mask_Bool) : (memOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool_rbuf,MemOut_CTmain_mask_Bool) */
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_buf;
  assign memOut_CTmain_mask_Bool_r = (! memOut_CTmain_mask_Bool_buf[0]);
  assign memOut_CTmain_mask_Bool_rbuf_d = (memOut_CTmain_mask_Bool_buf[0] ? memOut_CTmain_mask_Bool_buf :
                                           memOut_CTmain_mask_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTmain_mask_Bool_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTmain_mask_Bool_rbuf_r && memOut_CTmain_mask_Bool_buf[0]))
        memOut_CTmain_mask_Bool_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTmain_mask_Bool_rbuf_r) && (! memOut_CTmain_mask_Bool_buf[0])))
        memOut_CTmain_mask_Bool_buf <= memOut_CTmain_mask_Bool_d;
  
  /* destruct (Ty Pointer_CTmain_mask_Bool,
          Dcon Pointer_CTmain_mask_Bool) : (scfarg_0_1_1_argbuf,Pointer_CTmain_mask_Bool) > [(destructReadIn_CTmain_mask_Bool,Word16#)] */
  assign destructReadIn_CTmain_mask_Bool_d = {scfarg_0_1_1_argbuf_d[16:1],
                                              scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CTmain_mask_Bool_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Bool,
      Dcon ReadIn_CTmain_mask_Bool) : [(destructReadIn_CTmain_mask_Bool,Word16#)] > (dconReadIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  assign dconReadIn_CTmain_mask_Bool_d = ReadIn_CTmain_mask_Bool_dc((& {destructReadIn_CTmain_mask_Bool_d[0]}), destructReadIn_CTmain_mask_Bool_d);
  assign {destructReadIn_CTmain_mask_Bool_r} = {1 {(dconReadIn_CTmain_mask_Bool_r && dconReadIn_CTmain_mask_Bool_d[0])}};
  
  /* destruct (Ty MemOut_CTmain_mask_Bool,
          Dcon ReadOut_CTmain_mask_Bool) : (memReadOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) > [(readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf,CTmain_mask_Bool)] */
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d = {memReadOut_CTmain_mask_Bool_d[116:2],
                                                              memReadOut_CTmain_mask_Bool_d[0]};
  assign memReadOut_CTmain_mask_Bool_r = readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTmain_mask_Bool) : [(lizzieLet18_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet26_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet27_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet28_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet9_1_argbuf,CTmain_mask_Bool)] > (writeMerge_choice_CTmain_mask_Bool,C5) (writeMerge_data_CTmain_mask_Bool,CTmain_mask_Bool) */
  logic [4:0] lizzieLet18_1_argbuf_select_d;
  assign lizzieLet18_1_argbuf_select_d = ((| lizzieLet18_1_argbuf_select_q) ? lizzieLet18_1_argbuf_select_q :
                                          (lizzieLet18_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet26_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet27_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet28_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet9_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet18_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet18_1_argbuf_select_q <= (lizzieLet18_1_argbuf_done ? 5'd0 :
                                        lizzieLet18_1_argbuf_select_d);
  logic [1:0] lizzieLet18_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet18_1_argbuf_emit_q <= (lizzieLet18_1_argbuf_done ? 2'd0 :
                                      lizzieLet18_1_argbuf_emit_d);
  logic [1:0] lizzieLet18_1_argbuf_emit_d;
  assign lizzieLet18_1_argbuf_emit_d = (lizzieLet18_1_argbuf_emit_q | ({writeMerge_choice_CTmain_mask_Bool_d[0],
                                                                        writeMerge_data_CTmain_mask_Bool_d[0]} & {writeMerge_choice_CTmain_mask_Bool_r,
                                                                                                                  writeMerge_data_CTmain_mask_Bool_r}));
  logic lizzieLet18_1_argbuf_done;
  assign lizzieLet18_1_argbuf_done = (& lizzieLet18_1_argbuf_emit_d);
  assign {lizzieLet9_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet18_1_argbuf_r} = (lizzieLet18_1_argbuf_done ? lizzieLet18_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTmain_mask_Bool_d = ((lizzieLet18_1_argbuf_select_d[0] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                               ((lizzieLet18_1_argbuf_select_d[1] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                ((lizzieLet18_1_argbuf_select_d[2] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                                 ((lizzieLet18_1_argbuf_select_d[3] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                                  ((lizzieLet18_1_argbuf_select_d[4] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                   {115'd0, 1'd0})))));
  assign writeMerge_choice_CTmain_mask_Bool_d = ((lizzieLet18_1_argbuf_select_d[0] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                 ((lizzieLet18_1_argbuf_select_d[1] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                  ((lizzieLet18_1_argbuf_select_d[2] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                   ((lizzieLet18_1_argbuf_select_d[3] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                    ((lizzieLet18_1_argbuf_select_d[4] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                     {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_mask_Bool) : (writeMerge_choice_CTmain_mask_Bool,C5) (demuxWriteResult_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) > [(writeCTmain_mask_BoollizzieLet18_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet26_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet27_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet28_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet9_1_argbuf,Pointer_CTmain_mask_Bool)] */
  logic [4:0] demuxWriteResult_CTmain_mask_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_CTmain_mask_Bool_d[0] && demuxWriteResult_CTmain_mask_Bool_d[0]))
      unique case (writeMerge_choice_CTmain_mask_Bool_d[3:1])
        3'd0: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd16;
        default: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd0;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[0]};
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[1]};
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[2]};
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[3]};
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Bool_onehotd[4]};
  assign demuxWriteResult_CTmain_mask_Bool_r = (| (demuxWriteResult_CTmain_mask_Bool_onehotd & {writeCTmain_mask_BoollizzieLet9_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet28_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet27_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet26_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet18_1_argbuf_r}));
  assign writeMerge_choice_CTmain_mask_Bool_r = demuxWriteResult_CTmain_mask_Bool_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Bool,
      Dcon WriteIn_CTmain_mask_Bool) : [(forkHP1_CTmain_mask_Boo2,Word16#),
                                        (writeMerge_data_CTmain_mask_Bool,CTmain_mask_Bool)] > (dconWriteIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  assign dconWriteIn_CTmain_mask_Bool_d = WriteIn_CTmain_mask_Bool_dc((& {forkHP1_CTmain_mask_Boo2_d[0],
                                                                          writeMerge_data_CTmain_mask_Bool_d[0]}), forkHP1_CTmain_mask_Boo2_d, writeMerge_data_CTmain_mask_Bool_d);
  assign {forkHP1_CTmain_mask_Boo2_r,
          writeMerge_data_CTmain_mask_Bool_r} = {2 {(dconWriteIn_CTmain_mask_Bool_r && dconWriteIn_CTmain_mask_Bool_d[0])}};
  
  /* dcon (Ty Pointer_CTmain_mask_Bool,
      Dcon Pointer_CTmain_mask_Bool) : [(forkHP1_CTmain_mask_Boo3,Word16#)] > (dconPtr_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) */
  assign dconPtr_CTmain_mask_Bool_d = Pointer_CTmain_mask_Bool_dc((& {forkHP1_CTmain_mask_Boo3_d[0]}), forkHP1_CTmain_mask_Boo3_d);
  assign {forkHP1_CTmain_mask_Boo3_r} = {1 {(dconPtr_CTmain_mask_Bool_r && dconPtr_CTmain_mask_Bool_d[0])}};
  
  /* demux (Ty MemOut_CTmain_mask_Bool,
       Ty Pointer_CTmain_mask_Bool) : (memWriteOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) (dconPtr_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) > [(_47,Pointer_CTmain_mask_Bool),
                                                                                                                                                    (demuxWriteResult_CTmain_mask_Bool,Pointer_CTmain_mask_Bool)] */
  logic [1:0] dconPtr_CTmain_mask_Bool_onehotd;
  always_comb
    if ((memWriteOut_CTmain_mask_Bool_d[0] && dconPtr_CTmain_mask_Bool_d[0]))
      unique case (memWriteOut_CTmain_mask_Bool_d[1:1])
        1'd0: dconPtr_CTmain_mask_Bool_onehotd = 2'd1;
        1'd1: dconPtr_CTmain_mask_Bool_onehotd = 2'd2;
        default: dconPtr_CTmain_mask_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_CTmain_mask_Bool_onehotd = 2'd0;
  assign _47_d = {dconPtr_CTmain_mask_Bool_d[16:1],
                  dconPtr_CTmain_mask_Bool_onehotd[0]};
  assign demuxWriteResult_CTmain_mask_Bool_d = {dconPtr_CTmain_mask_Bool_d[16:1],
                                                dconPtr_CTmain_mask_Bool_onehotd[1]};
  assign dconPtr_CTmain_mask_Bool_r = (| (dconPtr_CTmain_mask_Bool_onehotd & {demuxWriteResult_CTmain_mask_Bool_r,
                                                                              _47_r}));
  assign memWriteOut_CTmain_mask_Bool_r = dconPtr_CTmain_mask_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  logic [31:0] profiling_MemIn_MaskQTree_read;
  logic [31:0] profiling_MemIn_MaskQTree_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_MaskQTree_write <= 0;
        profiling_MemIn_MaskQTree_read <= 0;
      end
    else
      if ((memMergeIn_MaskQTree_dbuf_we == 1'd1))
        profiling_MemIn_MaskQTree_write <= (profiling_MemIn_MaskQTree_write + 1);
      else
        if ((memOut_MaskQTree_valid == 1'd1))
          profiling_MemIn_MaskQTree_read <= (profiling_MemIn_MaskQTree_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (mskacj_1_argbuf,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {mskacj_1_argbuf_d[16:1],
                                       mskacj_1_argbuf_d[0]};
  assign mskacj_1_argbuf_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(readPointer_MaskQTreemskacj_1_argbuf,MaskQTree)] */
  assign readPointer_MaskQTreemskacj_1_argbuf_d = {memReadOut_MaskQTree_d[67:2],
                                                   memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = readPointer_MaskQTreemskacj_1_argbuf_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_46,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _46_d = {dconPtr_MaskQTree_d[16:1],
                  dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _46_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1acS_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m2acT_1,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m3acU_2,Pointer_QTree_Bool) */
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyBool,
          Dcon TupGo___MyDTBool_Bool___MyBool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) > [(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2,Go),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done;
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[1:1],
                                                                   (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted | ({applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]} & {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r ? 3'd0 :
                                                                     applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool) > [(arg0_1,MyDTBool_Bool),
                                                                                                  (arg0_2,MyDTBool_Bool),
                                                                                                  (arg0_3,MyDTBool_Bool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done;
  assign arg0_1_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[0]));
  assign arg0_2_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[1]));
  assign arg0_3_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[2]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted | ({arg0_3_d[0],
                                                                                                                                       arg0_2_d[0],
                                                                                                                                       arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                                       arg0_2_r,
                                                                                                                                                       arg0_1_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r ? 3'd0 :
                                                                       applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  
  /* fork (Ty MyBool) : (applyfnBool_Bool_5_resbuf,MyBool) > [(es_0_1_1,MyBool),
                                                         (es_0_1_2,MyBool),
                                                         (es_0_1_3,MyBool)] */
  logic [2:0] applyfnBool_Bool_5_resbuf_emitted;
  logic [2:0] applyfnBool_Bool_5_resbuf_done;
  assign es_0_1_1_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[0]))};
  assign es_0_1_2_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[1]))};
  assign es_0_1_3_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[2]))};
  assign applyfnBool_Bool_5_resbuf_done = (applyfnBool_Bool_5_resbuf_emitted | ({es_0_1_3_d[0],
                                                                                 es_0_1_2_d[0],
                                                                                 es_0_1_1_d[0]} & {es_0_1_3_r,
                                                                                                   es_0_1_2_r,
                                                                                                   es_0_1_1_r}));
  assign applyfnBool_Bool_5_resbuf_r = (& applyfnBool_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnBool_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnBool_Bool_5_resbuf_emitted <= (applyfnBool_Bool_5_resbuf_r ? 3'd0 :
                                            applyfnBool_Bool_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
          Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) > [(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2,MyDTBool_Bool_Bool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1,MyBool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done;
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[1:1],
                                                                                      (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[2:2],
                                                                                        (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[3]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted | ({applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]} & {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r ? 4'd0 :
                                                                                        applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool_Bool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2,MyDTBool_Bool_Bool) > [(arg0_2_1,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_2_2,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_2_3,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_2_4,MyDTBool_Bool_Bool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_done;
  assign arg0_2_1_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted[2]));
  assign arg0_2_4_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted[3]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted | ({arg0_2_4_d[0],
                                                                                                                                                                                 arg0_2_3_d[0],
                                                                                                                                                                                 arg0_2_2_d[0],
                                                                                                                                                                                 arg0_2_1_d[0]} & {arg0_2_4_r,
                                                                                                                                                                                                   arg0_2_3_r,
                                                                                                                                                                                                   arg0_2_2_r,
                                                                                                                                                                                                   arg0_2_1_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_r ? 4'd0 :
                                                                                            applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_2_done);
  
  /* fork (Ty MyBool) : (applyfnBool_Bool_Bool_5_resbuf,MyBool) > [(xabY_1,MyBool),
                                                              (xabY_2,MyBool)] */
  logic [1:0] applyfnBool_Bool_Bool_5_resbuf_emitted;
  logic [1:0] applyfnBool_Bool_Bool_5_resbuf_done;
  assign xabY_1_d = {applyfnBool_Bool_Bool_5_resbuf_d[1:1],
                     (applyfnBool_Bool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_Bool_5_resbuf_emitted[0]))};
  assign xabY_2_d = {applyfnBool_Bool_Bool_5_resbuf_d[1:1],
                     (applyfnBool_Bool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_Bool_5_resbuf_emitted[1]))};
  assign applyfnBool_Bool_Bool_5_resbuf_done = (applyfnBool_Bool_Bool_5_resbuf_emitted | ({xabY_2_d[0],
                                                                                           xabY_1_d[0]} & {xabY_2_r,
                                                                                                           xabY_1_r}));
  assign applyfnBool_Bool_Bool_5_resbuf_r = (& applyfnBool_Bool_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5_resbuf_emitted <= 2'd0;
    else
      applyfnBool_Bool_Bool_5_resbuf_emitted <= (applyfnBool_Bool_Bool_5_resbuf_r ? 2'd0 :
                                                 applyfnBool_Bool_Bool_5_resbuf_done);
  
  /* demux (Ty MyDTBool_Bool,
       Ty MyBool) : (arg0_1,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool) > [(arg0_1Dcon_main1,MyBool)] */
  assign arg0_1Dcon_main1_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[1:1],
                               (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0])};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  
  /* fork (Ty MyBool) : (arg0_1Dcon_main1,MyBool) > [(arg0_1Dcon_main1_1,MyBool),
                                                (arg0_1Dcon_main1_2,MyBool)] */
  logic [1:0] arg0_1Dcon_main1_emitted;
  logic [1:0] arg0_1Dcon_main1_done;
  assign arg0_1Dcon_main1_1_d = {arg0_1Dcon_main1_d[1:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[0]))};
  assign arg0_1Dcon_main1_2_d = {arg0_1Dcon_main1_d[1:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[1]))};
  assign arg0_1Dcon_main1_done = (arg0_1Dcon_main1_emitted | ({arg0_1Dcon_main1_2_d[0],
                                                               arg0_1Dcon_main1_1_d[0]} & {arg0_1Dcon_main1_2_r,
                                                                                           arg0_1Dcon_main1_1_r}));
  assign arg0_1Dcon_main1_r = (& arg0_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_main1_emitted <= 2'd0;
    else
      arg0_1Dcon_main1_emitted <= (arg0_1Dcon_main1_r ? 2'd0 :
                                   arg0_1Dcon_main1_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_1Dcon_main1_1,MyBool) (arg0_2Dcon_main1,Go) > [(arg0_1Dcon_main1_1MyFalse,Go),
                                                                     (arg0_1Dcon_main1_1MyTrue,Go)] */
  logic [1:0] arg0_2Dcon_main1_onehotd;
  always_comb
    if ((arg0_1Dcon_main1_1_d[0] && arg0_2Dcon_main1_d[0]))
      unique case (arg0_1Dcon_main1_1_d[1:1])
        1'd0: arg0_2Dcon_main1_onehotd = 2'd1;
        1'd1: arg0_2Dcon_main1_onehotd = 2'd2;
        default: arg0_2Dcon_main1_onehotd = 2'd0;
      endcase
    else arg0_2Dcon_main1_onehotd = 2'd0;
  assign arg0_1Dcon_main1_1MyFalse_d = arg0_2Dcon_main1_onehotd[0];
  assign arg0_1Dcon_main1_1MyTrue_d = arg0_2Dcon_main1_onehotd[1];
  assign arg0_2Dcon_main1_r = (| (arg0_2Dcon_main1_onehotd & {arg0_1Dcon_main1_1MyTrue_r,
                                                              arg0_1Dcon_main1_1MyFalse_r}));
  assign arg0_1Dcon_main1_1_r = arg0_2Dcon_main1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(arg0_1Dcon_main1_1MyFalse,Go)] > (arg0_1Dcon_main1_1MyFalse_1MyTrue,MyBool) */
  assign arg0_1Dcon_main1_1MyFalse_1MyTrue_d = MyTrue_dc((& {arg0_1Dcon_main1_1MyFalse_d[0]}), arg0_1Dcon_main1_1MyFalse_d);
  assign {arg0_1Dcon_main1_1MyFalse_r} = {1 {(arg0_1Dcon_main1_1MyFalse_1MyTrue_r && arg0_1Dcon_main1_1MyFalse_1MyTrue_d[0])}};
  
  /* buf (Ty MyBool) : (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux,MyBool) > (applyfnBool_Bool_5_resbuf,MyBool) */
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r;
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r = ((! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d[0]) || arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d <= {1'd0,
                                                                                               1'd0};
    else
      if (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r)
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d <= arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf;
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r = (! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]);
  assign applyfnBool_Bool_5_resbuf_d = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0] ? arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf :
                                        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                 1'd0};
    else
      if ((applyfnBool_Bool_5_resbuf_r && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]))
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                   1'd0};
      else if (((! applyfnBool_Bool_5_resbuf_r) && (! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0])))
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(arg0_1Dcon_main1_1MyTrue,Go)] > (arg0_1Dcon_main1_1MyTrue_1MyFalse,MyBool) */
  assign arg0_1Dcon_main1_1MyTrue_1MyFalse_d = MyFalse_dc((& {arg0_1Dcon_main1_1MyTrue_d[0]}), arg0_1Dcon_main1_1MyTrue_d);
  assign {arg0_1Dcon_main1_1MyTrue_r} = {1 {(arg0_1Dcon_main1_1MyTrue_1MyFalse_r && arg0_1Dcon_main1_1MyTrue_1MyFalse_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_1Dcon_main1_2,MyBool) [(arg0_1Dcon_main1_1MyFalse_1MyTrue,MyBool),
                                               (arg0_1Dcon_main1_1MyTrue_1MyFalse,MyBool)] > (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux,MyBool) */
  logic [1:0] arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux;
  logic [1:0] arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot;
  always_comb
    unique case (arg0_1Dcon_main1_2_d[1:1])
      1'd0:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd1,
                                                                                        arg0_1Dcon_main1_1MyFalse_1MyTrue_d};
      1'd1:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd2,
                                                                                        arg0_1Dcon_main1_1MyTrue_1MyFalse_d};
      default:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd0,
                                                                                        {1'd0,
                                                                                         1'd0}};
    endcase
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d = {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux[1:1],
                                                                                     (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux[0] && arg0_1Dcon_main1_2_d[0])};
  assign arg0_1Dcon_main1_2_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r);
  assign {arg0_1Dcon_main1_1MyTrue_1MyFalse_r,
          arg0_1Dcon_main1_1MyFalse_1MyTrue_r} = (arg0_1Dcon_main1_2_r ? arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot :
                                                  2'd0);
  
  /* demux (Ty MyDTBool_Bool,
       Ty Go) : (arg0_2,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2,Go) > [(arg0_2Dcon_main1,Go)] */
  assign arg0_2Dcon_main1_d = (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]);
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]));
  assign arg0_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]));
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_2_1,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1,MyBool) > [(arg0_2_1Dcon_&&,MyBool)] */
  assign \arg0_2_1Dcon_&&_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d[1:1],
                                (arg0_2_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_r = (\arg0_2_1Dcon_&&_r  && (arg0_2_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d[0]));
  assign arg0_2_1_r = (\arg0_2_1Dcon_&&_r  && (arg0_2_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_1_d[0]));
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_2_2,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool) > [(arg0_2_2Dcon_&&,MyBool)] */
  assign \arg0_2_2Dcon_&&_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[1:1],
                                (arg0_2_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r = (\arg0_2_2Dcon_&&_r  && (arg0_2_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  assign arg0_2_2_r = (\arg0_2_2Dcon_&&_r  && (arg0_2_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  
  /* fork (Ty MyBool) : (arg0_2_2Dcon_&&,MyBool) > [(arg0_2_2Dcon_&&_1,MyBool),
                                               (arg0_2_2Dcon_&&_2,MyBool),
                                               (arg0_2_2Dcon_&&_3,MyBool)] */
  logic [2:0] \arg0_2_2Dcon_&&_emitted ;
  logic [2:0] \arg0_2_2Dcon_&&_done ;
  assign \arg0_2_2Dcon_&&_1_d  = {\arg0_2_2Dcon_&&_d [1:1],
                                  (\arg0_2_2Dcon_&&_d [0] && (! \arg0_2_2Dcon_&&_emitted [0]))};
  assign \arg0_2_2Dcon_&&_2_d  = {\arg0_2_2Dcon_&&_d [1:1],
                                  (\arg0_2_2Dcon_&&_d [0] && (! \arg0_2_2Dcon_&&_emitted [1]))};
  assign \arg0_2_2Dcon_&&_3_d  = {\arg0_2_2Dcon_&&_d [1:1],
                                  (\arg0_2_2Dcon_&&_d [0] && (! \arg0_2_2Dcon_&&_emitted [2]))};
  assign \arg0_2_2Dcon_&&_done  = (\arg0_2_2Dcon_&&_emitted  | ({\arg0_2_2Dcon_&&_3_d [0],
                                                                 \arg0_2_2Dcon_&&_2_d [0],
                                                                 \arg0_2_2Dcon_&&_1_d [0]} & {\arg0_2_2Dcon_&&_3_r ,
                                                                                              \arg0_2_2Dcon_&&_2_r ,
                                                                                              \arg0_2_2Dcon_&&_1_r }));
  assign \arg0_2_2Dcon_&&_r  = (& \arg0_2_2Dcon_&&_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_2Dcon_&&_emitted  <= 3'd0;
    else
      \arg0_2_2Dcon_&&_emitted  <= (\arg0_2_2Dcon_&&_r  ? 3'd0 :
                                    \arg0_2_2Dcon_&&_done );
  
  /* demux (Ty MyBool,
       Ty MyBool) : (arg0_2_2Dcon_&&_1,MyBool) (arg0_2_1Dcon_&&,MyBool) > [(_45,MyBool),
                                                                           (arg0_2_2Dcon_&&_1MyTrue,MyBool)] */
  logic [1:0] \arg0_2_1Dcon_&&_onehotd ;
  always_comb
    if ((\arg0_2_2Dcon_&&_1_d [0] && \arg0_2_1Dcon_&&_d [0]))
      unique case (\arg0_2_2Dcon_&&_1_d [1:1])
        1'd0: \arg0_2_1Dcon_&&_onehotd  = 2'd1;
        1'd1: \arg0_2_1Dcon_&&_onehotd  = 2'd2;
        default: \arg0_2_1Dcon_&&_onehotd  = 2'd0;
      endcase
    else \arg0_2_1Dcon_&&_onehotd  = 2'd0;
  assign _45_d = {\arg0_2_1Dcon_&&_d [1:1],
                  \arg0_2_1Dcon_&&_onehotd [0]};
  assign \arg0_2_2Dcon_&&_1MyTrue_d  = {\arg0_2_1Dcon_&&_d [1:1],
                                        \arg0_2_1Dcon_&&_onehotd [1]};
  assign \arg0_2_1Dcon_&&_r  = (| (\arg0_2_1Dcon_&&_onehotd  & {\arg0_2_2Dcon_&&_1MyTrue_r ,
                                                                _45_r}));
  assign \arg0_2_2Dcon_&&_1_r  = \arg0_2_1Dcon_&&_r ;
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_2_2Dcon_&&_2,MyBool) (arg0_2_3Dcon_&&,Go) > [(arg0_2_2Dcon_&&_2MyFalse,Go),
                                                                   (_44,Go)] */
  logic [1:0] \arg0_2_3Dcon_&&_onehotd ;
  always_comb
    if ((\arg0_2_2Dcon_&&_2_d [0] && \arg0_2_3Dcon_&&_d [0]))
      unique case (\arg0_2_2Dcon_&&_2_d [1:1])
        1'd0: \arg0_2_3Dcon_&&_onehotd  = 2'd1;
        1'd1: \arg0_2_3Dcon_&&_onehotd  = 2'd2;
        default: \arg0_2_3Dcon_&&_onehotd  = 2'd0;
      endcase
    else \arg0_2_3Dcon_&&_onehotd  = 2'd0;
  assign \arg0_2_2Dcon_&&_2MyFalse_d  = \arg0_2_3Dcon_&&_onehotd [0];
  assign _44_d = \arg0_2_3Dcon_&&_onehotd [1];
  assign \arg0_2_3Dcon_&&_r  = (| (\arg0_2_3Dcon_&&_onehotd  & {_44_r,
                                                                \arg0_2_2Dcon_&&_2MyFalse_r }));
  assign \arg0_2_2Dcon_&&_2_r  = \arg0_2_3Dcon_&&_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(arg0_2_2Dcon_&&_2MyFalse,Go)] > (arg0_2_2Dcon_&&_2MyFalse_1MyFalse,MyBool) */
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_d  = MyFalse_dc((& {\arg0_2_2Dcon_&&_2MyFalse_d [0]}), \arg0_2_2Dcon_&&_2MyFalse_d );
  assign {\arg0_2_2Dcon_&&_2MyFalse_r } = {1 {(\arg0_2_2Dcon_&&_2MyFalse_1MyFalse_r  && \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_d [0])}};
  
  /* buf (Ty MyBool) : (arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux,MyBool) > (applyfnBool_Bool_Bool_5_resbuf,MyBool) */
  MyBool_t \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d ;
  logic \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r ;
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_r  = ((! \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d [0]) || \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d  <= {1'd0,
                                                                                         1'd0};
    else
      if (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_r )
        \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d  <= \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_d ;
  MyBool_t \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf ;
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r  = (! \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0]);
  assign applyfnBool_Bool_Bool_5_resbuf_d = (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0] ? \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  :
                                             \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= {1'd0,
                                                                                           1'd0};
    else
      if ((applyfnBool_Bool_Bool_5_resbuf_r && \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0]))
        \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= {1'd0,
                                                                                             1'd0};
      else if (((! applyfnBool_Bool_Bool_5_resbuf_r) && (! \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0])))
        \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d ;
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_2_2Dcon_&&_3,MyBool) [(arg0_2_2Dcon_&&_2MyFalse_1MyFalse,MyBool),
                                              (arg0_2_2Dcon_&&_1MyTrue,MyBool)] > (arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux,MyBool) */
  logic [1:0] \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux ;
  logic [1:0] \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_onehot ;
  always_comb
    unique case (\arg0_2_2Dcon_&&_3_d [1:1])
      1'd0:
        {\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd1,
                                                                                  \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_d };
      1'd1:
        {\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd2,
                                                                                  \arg0_2_2Dcon_&&_1MyTrue_d };
      default:
        {\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd0,
                                                                                  {1'd0, 1'd0}};
    endcase
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d  = {\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux [1:1],
                                                                               (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux [0] && \arg0_2_2Dcon_&&_3_d [0])};
  assign \arg0_2_2Dcon_&&_3_r  = (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d [0] && \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_r );
  assign {\arg0_2_2Dcon_&&_1MyTrue_r ,
          \arg0_2_2Dcon_&&_2MyFalse_1MyFalse_r } = (\arg0_2_2Dcon_&&_3_r  ? \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_onehot  :
                                                    2'd0);
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty Go) : (arg0_2_3,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go) > [(arg0_2_3Dcon_&&,Go)] */
  assign \arg0_2_3Dcon_&&_d  = (arg0_2_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]);
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r = (\arg0_2_3Dcon_&&_r  && (arg0_2_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  assign arg0_2_3_r = (\arg0_2_3Dcon_&&_r  && (arg0_2_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  
  /* mux (Ty MyDTBool_Bool_Bool,
     Ty MyBool) : (arg0_2_4,MyDTBool_Bool_Bool) [(arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux,MyBool)] > (arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux,MyBool) */
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_d  = {\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d [1:1],
                                                                                   (arg0_2_4_d[0] && \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d [0])};
  assign \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_r  = (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_r  && (arg0_2_4_d[0] && \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d [0]));
  assign arg0_2_4_r = (\arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_mux_r  && (arg0_2_4_d[0] && \arg0_2_2Dcon_&&_2MyFalse_1MyFalsearg0_2_2Dcon_&&_1MyTrue_1_mux_d [0]));
  
  /* mux (Ty MyDTBool_Bool,
     Ty MyBool) : (arg0_3,MyDTBool_Bool) [(arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux,MyBool)] > (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux,MyBool) */
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d = {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[1:1],
                                                                                         (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0])};
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0]));
  assign arg0_3_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) : (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) > [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [5:0] call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted;
  logic [5:0] call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done;
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[0]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[1]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[2]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[16:1],
                                                                                                                                                                          (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[3]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[32:17],
                                                                                                                                                                          (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[4]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[48:33],
                                                                                                                                                                         (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[5]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted | ({call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d[0]} & {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_r}));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r = (& call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted <= 6'd0;
    else
      call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted <= (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r ? 6'd0 :
                                                                                                                                                                           call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done);
  
  /* rbuf (Ty Go) : (call_kron_kron_Bool_Bool_Bool_goConst,Go) > (call_kron_kron_Bool_Bool_Bool_initBufi,Go) */
  Go_t call_kron_kron_Bool_Bool_Bool_goConst_buf;
  assign call_kron_kron_Bool_Bool_Bool_goConst_r = (! call_kron_kron_Bool_Bool_Bool_goConst_buf[0]);
  assign call_kron_kron_Bool_Bool_Bool_initBufi_d = (call_kron_kron_Bool_Bool_Bool_goConst_buf[0] ? call_kron_kron_Bool_Bool_Bool_goConst_buf :
                                                     call_kron_kron_Bool_Bool_Bool_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goConst_buf <= 1'd0;
    else
      if ((call_kron_kron_Bool_Bool_Bool_initBufi_r && call_kron_kron_Bool_Bool_Bool_goConst_buf[0]))
        call_kron_kron_Bool_Bool_Bool_goConst_buf <= 1'd0;
      else if (((! call_kron_kron_Bool_Bool_Bool_initBufi_r) && (! call_kron_kron_Bool_Bool_Bool_goConst_buf[0])))
        call_kron_kron_Bool_Bool_Bool_goConst_buf <= call_kron_kron_Bool_Bool_Bool_goConst_d;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_kron_kron_Bool_Bool_Bool_goMux1,Go),
                     (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf,Go),
                     (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf,Go),
                     (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf,Go),
                     (lizzieLet0_4QNode_Bool_1_argbuf,Go)] > (go_4_goMux_choice,C5) (go_4_goMux_data,Go) */
  logic [4:0] call_kron_kron_Bool_Bool_Bool_goMux1_select_d;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_select_d = ((| call_kron_kron_Bool_Bool_Bool_goMux1_select_q) ? call_kron_kron_Bool_Bool_Bool_goMux1_select_q :
                                                          (call_kron_kron_Bool_Bool_Bool_goMux1_d[0] ? 5'd1 :
                                                           (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d[0] ? 5'd2 :
                                                            (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d[0] ? 5'd4 :
                                                             (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d[0] ? 5'd8 :
                                                              (lizzieLet0_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                               5'd0))))));
  logic [4:0] call_kron_kron_Bool_Bool_Bool_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goMux1_select_q <= 5'd0;
    else
      call_kron_kron_Bool_Bool_Bool_goMux1_select_q <= (call_kron_kron_Bool_Bool_Bool_goMux1_done ? 5'd0 :
                                                        call_kron_kron_Bool_Bool_Bool_goMux1_select_d);
  logic [1:0] call_kron_kron_Bool_Bool_Bool_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goMux1_emit_q <= 2'd0;
    else
      call_kron_kron_Bool_Bool_Bool_goMux1_emit_q <= (call_kron_kron_Bool_Bool_Bool_goMux1_done ? 2'd0 :
                                                      call_kron_kron_Bool_Bool_Bool_goMux1_emit_d);
  logic [1:0] call_kron_kron_Bool_Bool_Bool_goMux1_emit_d;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_emit_d = (call_kron_kron_Bool_Bool_Bool_goMux1_emit_q | ({go_4_goMux_choice_d[0],
                                                                                                        go_4_goMux_data_d[0]} & {go_4_goMux_choice_r,
                                                                                                                                 go_4_goMux_data_r}));
  logic call_kron_kron_Bool_Bool_Bool_goMux1_done;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_done = (& call_kron_kron_Bool_Bool_Bool_goMux1_emit_d);
  assign {lizzieLet0_4QNode_Bool_1_argbuf_r,
          lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r,
          lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r,
          lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux1_r} = (call_kron_kron_Bool_Bool_Bool_goMux1_done ? call_kron_kron_Bool_Bool_Bool_goMux1_select_d :
                                                     5'd0);
  assign go_4_goMux_data_d = ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[0] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? call_kron_kron_Bool_Bool_Bool_goMux1_d :
                              ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[1] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d :
                               ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[2] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d :
                                ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[3] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d :
                                 ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[4] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet0_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_4_goMux_choice_d = ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[0] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[1] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[2] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[3] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[4] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_kron_kron_Bool_Bool_Bool_initBuf,Go) > [(call_kron_kron_Bool_Bool_Bool_unlockFork1,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork2,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork3,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork4,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork5,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork6,Go)] */
  logic [5:0] call_kron_kron_Bool_Bool_Bool_initBuf_emitted;
  logic [5:0] call_kron_kron_Bool_Bool_Bool_initBuf_done;
  assign call_kron_kron_Bool_Bool_Bool_unlockFork1_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork2_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[1]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork3_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[2]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork4_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[3]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork5_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[4]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork6_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[5]));
  assign call_kron_kron_Bool_Bool_Bool_initBuf_done = (call_kron_kron_Bool_Bool_Bool_initBuf_emitted | ({call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0]} & {call_kron_kron_Bool_Bool_Bool_unlockFork6_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork5_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork4_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork3_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork2_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork1_r}));
  assign call_kron_kron_Bool_Bool_Bool_initBuf_r = (& call_kron_kron_Bool_Bool_Bool_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_initBuf_emitted <= 6'd0;
    else
      call_kron_kron_Bool_Bool_Bool_initBuf_emitted <= (call_kron_kron_Bool_Bool_Bool_initBuf_r ? 6'd0 :
                                                        call_kron_kron_Bool_Bool_Bool_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_kron_kron_Bool_Bool_Bool_initBufi,Go) > (call_kron_kron_Bool_Bool_Bool_initBuf,Go) */
  assign call_kron_kron_Bool_Bool_Bool_initBufi_r = ((! call_kron_kron_Bool_Bool_Bool_initBuf_d[0]) || call_kron_kron_Bool_Bool_Bool_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_initBuf_d <= Go_dc(1'd1);
    else
      if (call_kron_kron_Bool_Bool_Bool_initBufi_r)
        call_kron_kron_Bool_Bool_Bool_initBuf_d <= call_kron_kron_Bool_Bool_Bool_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_kron_kron_Bool_Bool_Bool_unlockFork1,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4,Go)] > (call_kron_kron_Bool_Bool_Bool_goMux1,Go) */
  assign call_kron_kron_Bool_Bool_Bool_goMux1_d = (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_r = (call_kron_kron_Bool_Bool_Bool_goMux1_r && (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork1_r = (call_kron_kron_Bool_Bool_Bool_goMux1_r && (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_4_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork2,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ,MyDTBool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux2,MyDTBool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux2_d = (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_r = (call_kron_kron_Bool_Bool_Bool_goMux2_r && (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork2_r = (call_kron_kron_Bool_Bool_Bool_goMux2_r && (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZacJ_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork3,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK,MyDTBool_Bool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux3_d = (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_r = (call_kron_kron_Bool_Bool_Bool_goMux3_r && (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork3_r = (call_kron_kron_Bool_Bool_Bool_goMux3_r && (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolgacK_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork4,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL,Pointer_QTree_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux4,Pointer_QTree_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux4_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_r = (call_kron_kron_Bool_Bool_Bool_goMux4_r && (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork4_r = (call_kron_kron_Bool_Bool_Bool_goMux4_r && (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1acL_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork5,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM,Pointer_QTree_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux5_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_r = (call_kron_kron_Bool_Bool_Bool_goMux5_r && (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork5_r = (call_kron_kron_Bool_Bool_Bool_goMux5_r && (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2acM_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork6,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0,Pointer_CTkron_kron_Bool_Bool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux6,Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux6_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r = (call_kron_kron_Bool_Bool_Bool_goMux6_r && (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork6_r = (call_kron_kron_Bool_Bool_Bool_goMux6_r && (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) : (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) > [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5,Go),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1,Pointer_CTmain_mask_Bool)] */
  logic [3:0] call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted;
  logic [3:0] call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done;
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d = (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[0]));
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[16:1],
                                                                                                               (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[1]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[32:17],
                                                                                                                 (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[2]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[48:33],
                                                                                                                 (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[3]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done = (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted | ({call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]} & {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r}));
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r = (& call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted <= 4'd0;
    else
      call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted <= (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r ? 4'd0 :
                                                                                                                 call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done);
  
  /* rbuf (Ty Go) : (call_main_mask_Bool_goConst,Go) > (call_main_mask_Bool_initBufi,Go) */
  Go_t call_main_mask_Bool_goConst_buf;
  assign call_main_mask_Bool_goConst_r = (! call_main_mask_Bool_goConst_buf[0]);
  assign call_main_mask_Bool_initBufi_d = (call_main_mask_Bool_goConst_buf[0] ? call_main_mask_Bool_goConst_buf :
                                           call_main_mask_Bool_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goConst_buf <= 1'd0;
    else
      if ((call_main_mask_Bool_initBufi_r && call_main_mask_Bool_goConst_buf[0]))
        call_main_mask_Bool_goConst_buf <= 1'd0;
      else if (((! call_main_mask_Bool_initBufi_r) && (! call_main_mask_Bool_goConst_buf[0])))
        call_main_mask_Bool_goConst_buf <= call_main_mask_Bool_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_mask_Bool_goMux1,Go),
                           (lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf,Go),
                           (lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf,Go),
                           (lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf,Go),
                           (lizzieLet4_4MQNode_3QNode_Bool_1_argbuf,Go)] > (go_5_goMux_choice,C5) (go_5_goMux_data,Go) */
  logic [4:0] call_main_mask_Bool_goMux1_select_d;
  assign call_main_mask_Bool_goMux1_select_d = ((| call_main_mask_Bool_goMux1_select_q) ? call_main_mask_Bool_goMux1_select_q :
                                                (call_main_mask_Bool_goMux1_d[0] ? 5'd1 :
                                                 (lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_d[0] ? 5'd2 :
                                                  (lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_d[0] ? 5'd4 :
                                                   (lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_d[0] ? 5'd8 :
                                                    (lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                     5'd0))))));
  logic [4:0] call_main_mask_Bool_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goMux1_select_q <= 5'd0;
    else
      call_main_mask_Bool_goMux1_select_q <= (call_main_mask_Bool_goMux1_done ? 5'd0 :
                                              call_main_mask_Bool_goMux1_select_d);
  logic [1:0] call_main_mask_Bool_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goMux1_emit_q <= 2'd0;
    else
      call_main_mask_Bool_goMux1_emit_q <= (call_main_mask_Bool_goMux1_done ? 2'd0 :
                                            call_main_mask_Bool_goMux1_emit_d);
  logic [1:0] call_main_mask_Bool_goMux1_emit_d;
  assign call_main_mask_Bool_goMux1_emit_d = (call_main_mask_Bool_goMux1_emit_q | ({go_5_goMux_choice_d[0],
                                                                                    go_5_goMux_data_d[0]} & {go_5_goMux_choice_r,
                                                                                                             go_5_goMux_data_r}));
  logic call_main_mask_Bool_goMux1_done;
  assign call_main_mask_Bool_goMux1_done = (& call_main_mask_Bool_goMux1_emit_d);
  assign {lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_r,
          lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_r,
          lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_r,
          lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_r,
          call_main_mask_Bool_goMux1_r} = (call_main_mask_Bool_goMux1_done ? call_main_mask_Bool_goMux1_select_d :
                                           5'd0);
  assign go_5_goMux_data_d = ((call_main_mask_Bool_goMux1_select_d[0] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? call_main_mask_Bool_goMux1_d :
                              ((call_main_mask_Bool_goMux1_select_d[1] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_d :
                               ((call_main_mask_Bool_goMux1_select_d[2] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_d :
                                ((call_main_mask_Bool_goMux1_select_d[3] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_d :
                                 ((call_main_mask_Bool_goMux1_select_d[4] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_5_goMux_choice_d = ((call_main_mask_Bool_goMux1_select_d[0] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_main_mask_Bool_goMux1_select_d[1] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_main_mask_Bool_goMux1_select_d[2] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_main_mask_Bool_goMux1_select_d[3] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_main_mask_Bool_goMux1_select_d[4] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_mask_Bool_initBuf,Go) > [(call_main_mask_Bool_unlockFork1,Go),
                                                   (call_main_mask_Bool_unlockFork2,Go),
                                                   (call_main_mask_Bool_unlockFork3,Go),
                                                   (call_main_mask_Bool_unlockFork4,Go)] */
  logic [3:0] call_main_mask_Bool_initBuf_emitted;
  logic [3:0] call_main_mask_Bool_initBuf_done;
  assign call_main_mask_Bool_unlockFork1_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[0]));
  assign call_main_mask_Bool_unlockFork2_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[1]));
  assign call_main_mask_Bool_unlockFork3_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[2]));
  assign call_main_mask_Bool_unlockFork4_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[3]));
  assign call_main_mask_Bool_initBuf_done = (call_main_mask_Bool_initBuf_emitted | ({call_main_mask_Bool_unlockFork4_d[0],
                                                                                     call_main_mask_Bool_unlockFork3_d[0],
                                                                                     call_main_mask_Bool_unlockFork2_d[0],
                                                                                     call_main_mask_Bool_unlockFork1_d[0]} & {call_main_mask_Bool_unlockFork4_r,
                                                                                                                              call_main_mask_Bool_unlockFork3_r,
                                                                                                                              call_main_mask_Bool_unlockFork2_r,
                                                                                                                              call_main_mask_Bool_unlockFork1_r}));
  assign call_main_mask_Bool_initBuf_r = (& call_main_mask_Bool_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_initBuf_emitted <= 4'd0;
    else
      call_main_mask_Bool_initBuf_emitted <= (call_main_mask_Bool_initBuf_r ? 4'd0 :
                                              call_main_mask_Bool_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_mask_Bool_initBufi,Go) > (call_main_mask_Bool_initBuf,Go) */
  assign call_main_mask_Bool_initBufi_r = ((! call_main_mask_Bool_initBuf_d[0]) || call_main_mask_Bool_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_initBuf_d <= Go_dc(1'd1);
    else
      if (call_main_mask_Bool_initBufi_r)
        call_main_mask_Bool_initBuf_d <= call_main_mask_Bool_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_mask_Bool_unlockFork1,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5,Go)] > (call_main_mask_Bool_goMux1,Go) */
  assign call_main_mask_Bool_goMux1_d = (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]);
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r = (call_main_mask_Bool_goMux1_r && (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]));
  assign call_main_mask_Bool_unlockFork1_r = (call_main_mask_Bool_goMux1_r && (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_main_mask_Bool_unlockFork2,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci,Pointer_QTree_Bool)] > (call_main_mask_Bool_goMux2,Pointer_QTree_Bool) */
  assign call_main_mask_Bool_goMux2_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d[16:1],
                                         (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_r = (call_main_mask_Bool_goMux2_r && (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d[0]));
  assign call_main_mask_Bool_unlockFork2_r = (call_main_mask_Bool_goMux2_r && (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmaci_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_main_mask_Bool_unlockFork3,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj,Pointer_MaskQTree)] > (call_main_mask_Bool_goMux3,Pointer_MaskQTree) */
  assign call_main_mask_Bool_goMux3_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d[16:1],
                                         (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_r = (call_main_mask_Bool_goMux3_r && (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d[0]));
  assign call_main_mask_Bool_unlockFork3_r = (call_main_mask_Bool_goMux3_r && (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmskacj_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_mask_Bool) : (call_main_mask_Bool_unlockFork4,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1,Pointer_CTmain_mask_Bool)] > (call_main_mask_Bool_goMux4,Pointer_CTmain_mask_Bool) */
  assign call_main_mask_Bool_goMux4_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[16:1],
                                         (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r = (call_main_mask_Bool_goMux4_r && (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0]));
  assign call_main_mask_Bool_unlockFork4_r = (call_main_mask_Bool_goMux4_r && (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) : (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) > [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6,Go),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC,MyBool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [5:0] \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted ;
  logic [5:0] \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done ;
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [0]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [1]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [2]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [1:1],
                                                                                                                                                                    (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [3]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [17:2],
                                                                                                                                                                   (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [4]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [33:18],
                                                                                                                                                                     (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [5]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  | ({\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d [0]} & {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_r }));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  = (& \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  <= 6'd0;
    else
      \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  <= (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  ? 6'd0 :
                                                                                                                                                                     \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done );
  
  /* rbuf (Ty Go) : (call_map''_map''_Bool_Bool_Bool_goConst,Go) > (call_map''_map''_Bool_Bool_Bool_initBufi,Go) */
  Go_t \call_map''_map''_Bool_Bool_Bool_goConst_buf ;
  assign \call_map''_map''_Bool_Bool_Bool_goConst_r  = (! \call_map''_map''_Bool_Bool_Bool_goConst_buf [0]);
  assign \call_map''_map''_Bool_Bool_Bool_initBufi_d  = (\call_map''_map''_Bool_Bool_Bool_goConst_buf [0] ? \call_map''_map''_Bool_Bool_Bool_goConst_buf  :
                                                         \call_map''_map''_Bool_Bool_Bool_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= 1'd0;
    else
      if ((\call_map''_map''_Bool_Bool_Bool_initBufi_r  && \call_map''_map''_Bool_Bool_Bool_goConst_buf [0]))
        \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= 1'd0;
      else if (((! \call_map''_map''_Bool_Bool_Bool_initBufi_r ) && (! \call_map''_map''_Bool_Bool_Bool_goConst_buf [0])))
        \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= \call_map''_map''_Bool_Bool_Bool_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_map''_map''_Bool_Bool_Bool_goMux1,Go),
                     (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf,Go),
                     (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf,Go),
                     (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf,Go),
                     (lizzieLet11_1_4QNode_Bool_1_argbuf,Go)] > (go_6_goMux_choice,C5) (go_6_goMux_data,Go) */
  logic [4:0] \call_map''_map''_Bool_Bool_Bool_goMux1_select_d ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_select_d  = ((| \call_map''_map''_Bool_Bool_Bool_goMux1_select_q ) ? \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  :
                                                              (\call_map''_map''_Bool_Bool_Bool_goMux1_d [0] ? 5'd1 :
                                                               (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d [0] ? 5'd2 :
                                                                (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d [0] ? 5'd4 :
                                                                 (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d [0] ? 5'd8 :
                                                                  (lizzieLet11_1_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                                   5'd0))))));
  logic [4:0] \call_map''_map''_Bool_Bool_Bool_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  <= 5'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  <= (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? 5'd0 :
                                                            \call_map''_map''_Bool_Bool_Bool_goMux1_select_d );
  logic [1:0] \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  <= 2'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  <= (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? 2'd0 :
                                                          \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d );
  logic [1:0] \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d  = (\call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  | ({go_6_goMux_choice_d[0],
                                                                                                                go_6_goMux_data_d[0]} & {go_6_goMux_choice_r,
                                                                                                                                         go_6_goMux_data_r}));
  logic \call_map''_map''_Bool_Bool_Bool_goMux1_done ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_done  = (& \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d );
  assign {lizzieLet11_1_4QNode_Bool_1_argbuf_r,
          \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ,
          \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ,
          \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ,
          \call_map''_map''_Bool_Bool_Bool_goMux1_r } = (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? \call_map''_map''_Bool_Bool_Bool_goMux1_select_d  :
                                                         5'd0);
  assign go_6_goMux_data_d = ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [0] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \call_map''_map''_Bool_Bool_Bool_goMux1_d  :
                              ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [1] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d  :
                               ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [2] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d  :
                                ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [3] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d  :
                                 ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [4] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? lizzieLet11_1_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_6_goMux_choice_d = ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [0] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [1] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [2] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [3] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [4] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_map''_map''_Bool_Bool_Bool_initBuf,Go) > [(call_map''_map''_Bool_Bool_Bool_unlockFork1,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork2,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork3,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork4,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork5,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork6,Go)] */
  logic [5:0] \call_map''_map''_Bool_Bool_Bool_initBuf_emitted ;
  logic [5:0] \call_map''_map''_Bool_Bool_Bool_initBuf_done ;
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork1_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork2_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [1]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork3_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [2]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork4_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [3]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork5_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [4]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork6_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [5]));
  assign \call_map''_map''_Bool_Bool_Bool_initBuf_done  = (\call_map''_map''_Bool_Bool_Bool_initBuf_emitted  | ({\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0]} & {\call_map''_map''_Bool_Bool_Bool_unlockFork6_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork5_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork4_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork3_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork2_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork1_r }));
  assign \call_map''_map''_Bool_Bool_Bool_initBuf_r  = (& \call_map''_map''_Bool_Bool_Bool_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_initBuf_emitted  <= 6'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_initBuf_emitted  <= (\call_map''_map''_Bool_Bool_Bool_initBuf_r  ? 6'd0 :
                                                            \call_map''_map''_Bool_Bool_Bool_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_map''_map''_Bool_Bool_Bool_initBufi,Go) > (call_map''_map''_Bool_Bool_Bool_initBuf,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_initBufi_r  = ((! \call_map''_map''_Bool_Bool_Bool_initBuf_d [0]) || \call_map''_map''_Bool_Bool_Bool_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_map''_map''_Bool_Bool_Bool_initBufi_r )
        \call_map''_map''_Bool_Bool_Bool_initBuf_d  <= \call_map''_map''_Bool_Bool_Bool_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_map''_map''_Bool_Bool_Bool_unlockFork1,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6,Go)] > (call_map''_map''_Bool_Bool_Bool_goMux1,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_r  = (\call_map''_map''_Bool_Bool_Bool_goMux1_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork1_r  = (\call_map''_map''_Bool_Bool_Bool_goMux1_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_6_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork2,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA,MyDTBool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux2,MyDTBool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux2_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_r  = (\call_map''_map''_Bool_Bool_Bool_goMux2_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork2_r  = (\call_map''_map''_Bool_Bool_Bool_goMux2_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacA_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork3,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB,MyDTBool_Bool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux3_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_r  = (\call_map''_map''_Bool_Bool_Bool_goMux3_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork3_r  = (\call_map''_map''_Bool_Bool_Bool_goMux3_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacB_d [0]));
  
  /* mux (Ty Go,
     Ty MyBool) : (call_map''_map''_Bool_Bool_Bool_unlockFork4,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC,MyBool)] > (call_map''_map''_Bool_Bool_Bool_goMux4,MyBool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux4_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d [1:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_r  = (\call_map''_map''_Bool_Bool_Bool_goMux4_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork4_r  = (\call_map''_map''_Bool_Bool_Bool_goMux4_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'acC_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork5,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD,Pointer_QTree_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux5_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d [16:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_r  = (\call_map''_map''_Bool_Bool_Bool_goMux5_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork5_r  = (\call_map''_map''_Bool_Bool_Bool_goMux5_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolmacD_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork6,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux6,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux6_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [16:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r  = (\call_map''_map''_Bool_Bool_Bool_goMux6_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork6_r  = (\call_map''_map''_Bool_Bool_Bool_goMux6_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0]));
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_1_1,MyBool) (lizzieLet11_1_4QVal_Bool_3,Go) > [(es_0_1_1MyFalse,Go),
                                                                     (es_0_1_1MyTrue,Go)] */
  logic [1:0] lizzieLet11_1_4QVal_Bool_3_onehotd;
  always_comb
    if ((es_0_1_1_d[0] && lizzieLet11_1_4QVal_Bool_3_d[0]))
      unique case (es_0_1_1_d[1:1])
        1'd0: lizzieLet11_1_4QVal_Bool_3_onehotd = 2'd1;
        1'd1: lizzieLet11_1_4QVal_Bool_3_onehotd = 2'd2;
        default: lizzieLet11_1_4QVal_Bool_3_onehotd = 2'd0;
      endcase
    else lizzieLet11_1_4QVal_Bool_3_onehotd = 2'd0;
  assign es_0_1_1MyFalse_d = lizzieLet11_1_4QVal_Bool_3_onehotd[0];
  assign es_0_1_1MyTrue_d = lizzieLet11_1_4QVal_Bool_3_onehotd[1];
  assign lizzieLet11_1_4QVal_Bool_3_r = (| (lizzieLet11_1_4QVal_Bool_3_onehotd & {es_0_1_1MyTrue_r,
                                                                                  es_0_1_1MyFalse_r}));
  assign es_0_1_1_r = lizzieLet11_1_4QVal_Bool_3_r;
  
  /* buf (Ty Go) : (es_0_1_1MyFalse,Go) > (es_0_1_1MyFalse_1_argbuf,Go) */
  Go_t es_0_1_1MyFalse_bufchan_d;
  logic es_0_1_1MyFalse_bufchan_r;
  assign es_0_1_1MyFalse_r = ((! es_0_1_1MyFalse_bufchan_d[0]) || es_0_1_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_1_1MyFalse_r)
        es_0_1_1MyFalse_bufchan_d <= es_0_1_1MyFalse_d;
  Go_t es_0_1_1MyFalse_bufchan_buf;
  assign es_0_1_1MyFalse_bufchan_r = (! es_0_1_1MyFalse_bufchan_buf[0]);
  assign es_0_1_1MyFalse_1_argbuf_d = (es_0_1_1MyFalse_bufchan_buf[0] ? es_0_1_1MyFalse_bufchan_buf :
                                       es_0_1_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_1_1MyFalse_1_argbuf_r && es_0_1_1MyFalse_bufchan_buf[0]))
        es_0_1_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_1_1MyFalse_1_argbuf_r) && (! es_0_1_1MyFalse_bufchan_buf[0])))
        es_0_1_1MyFalse_bufchan_buf <= es_0_1_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_1_1MyTrue,Go) > [(es_0_1_1MyTrue_1,Go),
                                      (es_0_1_1MyTrue_2,Go)] */
  logic [1:0] es_0_1_1MyTrue_emitted;
  logic [1:0] es_0_1_1MyTrue_done;
  assign es_0_1_1MyTrue_1_d = (es_0_1_1MyTrue_d[0] && (! es_0_1_1MyTrue_emitted[0]));
  assign es_0_1_1MyTrue_2_d = (es_0_1_1MyTrue_d[0] && (! es_0_1_1MyTrue_emitted[1]));
  assign es_0_1_1MyTrue_done = (es_0_1_1MyTrue_emitted | ({es_0_1_1MyTrue_2_d[0],
                                                           es_0_1_1MyTrue_1_d[0]} & {es_0_1_1MyTrue_2_r,
                                                                                     es_0_1_1MyTrue_1_r}));
  assign es_0_1_1MyTrue_r = (& es_0_1_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_emitted <= 2'd0;
    else
      es_0_1_1MyTrue_emitted <= (es_0_1_1MyTrue_r ? 2'd0 :
                                 es_0_1_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(es_0_1_1MyTrue_1,Go)] > (es_0_1_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign es_0_1_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {es_0_1_1MyTrue_1_d[0]}), es_0_1_1MyTrue_1_d);
  assign {es_0_1_1MyTrue_1_r} = {1 {(es_0_1_1MyTrue_1QNone_Bool_r && es_0_1_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_1_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet14_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1_1MyTrue_1QNone_Bool_bufchan_d;
  logic es_0_1_1MyTrue_1QNone_Bool_bufchan_r;
  assign es_0_1_1MyTrue_1QNone_Bool_r = ((! es_0_1_1MyTrue_1QNone_Bool_bufchan_d[0]) || es_0_1_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_1MyTrue_1QNone_Bool_r)
        es_0_1_1MyTrue_1QNone_Bool_bufchan_d <= es_0_1_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t es_0_1_1MyTrue_1QNone_Bool_bufchan_buf;
  assign es_0_1_1MyTrue_1QNone_Bool_bufchan_r = (! es_0_1_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (es_0_1_1MyTrue_1QNone_Bool_bufchan_buf[0] ? es_0_1_1MyTrue_1QNone_Bool_bufchan_buf :
                                   es_0_1_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && es_0_1_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        es_0_1_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! es_0_1_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        es_0_1_1MyTrue_1QNone_Bool_bufchan_buf <= es_0_1_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (es_0_1_1MyTrue_2,Go) > (es_0_1_1MyTrue_2_argbuf,Go) */
  Go_t es_0_1_1MyTrue_2_bufchan_d;
  logic es_0_1_1MyTrue_2_bufchan_r;
  assign es_0_1_1MyTrue_2_r = ((! es_0_1_1MyTrue_2_bufchan_d[0]) || es_0_1_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_1_1MyTrue_2_r)
        es_0_1_1MyTrue_2_bufchan_d <= es_0_1_1MyTrue_2_d;
  Go_t es_0_1_1MyTrue_2_bufchan_buf;
  assign es_0_1_1MyTrue_2_bufchan_r = (! es_0_1_1MyTrue_2_bufchan_buf[0]);
  assign es_0_1_1MyTrue_2_argbuf_d = (es_0_1_1MyTrue_2_bufchan_buf[0] ? es_0_1_1MyTrue_2_bufchan_buf :
                                      es_0_1_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_1_1MyTrue_2_argbuf_r && es_0_1_1MyTrue_2_bufchan_buf[0]))
        es_0_1_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_1_1MyTrue_2_argbuf_r) && (! es_0_1_1MyTrue_2_bufchan_buf[0])))
        es_0_1_1MyTrue_2_bufchan_buf <= es_0_1_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_1_2,MyBool) (lizzieLet11_1_6QVal_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(es_0_1_2MyFalse,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (es_0_1_2MyTrue,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] lizzieLet11_1_6QVal_Bool_onehotd;
  always_comb
    if ((es_0_1_2_d[0] && lizzieLet11_1_6QVal_Bool_d[0]))
      unique case (es_0_1_2_d[1:1])
        1'd0: lizzieLet11_1_6QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet11_1_6QVal_Bool_onehotd = 2'd2;
        default: lizzieLet11_1_6QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet11_1_6QVal_Bool_onehotd = 2'd0;
  assign es_0_1_2MyFalse_d = {lizzieLet11_1_6QVal_Bool_d[16:1],
                              lizzieLet11_1_6QVal_Bool_onehotd[0]};
  assign es_0_1_2MyTrue_d = {lizzieLet11_1_6QVal_Bool_d[16:1],
                             lizzieLet11_1_6QVal_Bool_onehotd[1]};
  assign lizzieLet11_1_6QVal_Bool_r = (| (lizzieLet11_1_6QVal_Bool_onehotd & {es_0_1_2MyTrue_r,
                                                                              es_0_1_2MyFalse_r}));
  assign es_0_1_2_r = lizzieLet11_1_6QVal_Bool_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_1_2MyFalse,Pointer_CTmap''_map''_Bool_Bool_Bool) > (es_0_1_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyFalse_bufchan_d;
  logic es_0_1_2MyFalse_bufchan_r;
  assign es_0_1_2MyFalse_r = ((! es_0_1_2MyFalse_bufchan_d[0]) || es_0_1_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_1_2MyFalse_r)
        es_0_1_2MyFalse_bufchan_d <= es_0_1_2MyFalse_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyFalse_bufchan_buf;
  assign es_0_1_2MyFalse_bufchan_r = (! es_0_1_2MyFalse_bufchan_buf[0]);
  assign es_0_1_2MyFalse_1_argbuf_d = (es_0_1_2MyFalse_bufchan_buf[0] ? es_0_1_2MyFalse_bufchan_buf :
                                       es_0_1_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_2MyFalse_1_argbuf_r && es_0_1_2MyFalse_bufchan_buf[0]))
        es_0_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_2MyFalse_1_argbuf_r) && (! es_0_1_2MyFalse_bufchan_buf[0])))
        es_0_1_2MyFalse_bufchan_buf <= es_0_1_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_1_2MyTrue,Pointer_CTmap''_map''_Bool_Bool_Bool) > (es_0_1_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyTrue_bufchan_d;
  logic es_0_1_2MyTrue_bufchan_r;
  assign es_0_1_2MyTrue_r = ((! es_0_1_2MyTrue_bufchan_d[0]) || es_0_1_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_1_2MyTrue_r) es_0_1_2MyTrue_bufchan_d <= es_0_1_2MyTrue_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_1_2MyTrue_bufchan_buf;
  assign es_0_1_2MyTrue_bufchan_r = (! es_0_1_2MyTrue_bufchan_buf[0]);
  assign es_0_1_2MyTrue_1_argbuf_d = (es_0_1_2MyTrue_bufchan_buf[0] ? es_0_1_2MyTrue_bufchan_buf :
                                      es_0_1_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_2MyTrue_1_argbuf_r && es_0_1_2MyTrue_bufchan_buf[0]))
        es_0_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_2MyTrue_1_argbuf_r) && (! es_0_1_2MyTrue_bufchan_buf[0])))
        es_0_1_2MyTrue_bufchan_buf <= es_0_1_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (es_0_1_3,MyBool) (xabY_2,MyBool) > [(es_0_1_3MyFalse,MyBool),
                                                         (_43,MyBool)] */
  logic [1:0] xabY_2_onehotd;
  always_comb
    if ((es_0_1_3_d[0] && xabY_2_d[0]))
      unique case (es_0_1_3_d[1:1])
        1'd0: xabY_2_onehotd = 2'd1;
        1'd1: xabY_2_onehotd = 2'd2;
        default: xabY_2_onehotd = 2'd0;
      endcase
    else xabY_2_onehotd = 2'd0;
  assign es_0_1_3MyFalse_d = {xabY_2_d[1:1], xabY_2_onehotd[0]};
  assign _43_d = {xabY_2_d[1:1], xabY_2_onehotd[1]};
  assign xabY_2_r = (| (xabY_2_onehotd & {_43_r,
                                          es_0_1_3MyFalse_r}));
  assign es_0_1_3_r = xabY_2_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(es_0_1_3MyFalse,MyBool)] > (es_0_1_3MyFalse_1QVal_Bool,QTree_Bool) */
  assign es_0_1_3MyFalse_1QVal_Bool_d = QVal_Bool_dc((& {es_0_1_3MyFalse_d[0]}), es_0_1_3MyFalse_d);
  assign {es_0_1_3MyFalse_r} = {1 {(es_0_1_3MyFalse_1QVal_Bool_r && es_0_1_3MyFalse_1QVal_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_1_3MyFalse_1QVal_Bool,QTree_Bool) > (lizzieLet13_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1_3MyFalse_1QVal_Bool_bufchan_d;
  logic es_0_1_3MyFalse_1QVal_Bool_bufchan_r;
  assign es_0_1_3MyFalse_1QVal_Bool_r = ((! es_0_1_3MyFalse_1QVal_Bool_bufchan_d[0]) || es_0_1_3MyFalse_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_3MyFalse_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_3MyFalse_1QVal_Bool_r)
        es_0_1_3MyFalse_1QVal_Bool_bufchan_d <= es_0_1_3MyFalse_1QVal_Bool_d;
  QTree_Bool_t es_0_1_3MyFalse_1QVal_Bool_bufchan_buf;
  assign es_0_1_3MyFalse_1QVal_Bool_bufchan_r = (! es_0_1_3MyFalse_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (es_0_1_3MyFalse_1QVal_Bool_bufchan_buf[0] ? es_0_1_3MyFalse_1QVal_Bool_bufchan_buf :
                                   es_0_1_3MyFalse_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && es_0_1_3MyFalse_1QVal_Bool_bufchan_buf[0]))
        es_0_1_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! es_0_1_3MyFalse_1QVal_Bool_bufchan_buf[0])))
        es_0_1_3MyFalse_1QVal_Bool_bufchan_buf <= es_0_1_3MyFalse_1QVal_Bool_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacB_2_2,MyDTBool_Bool_Bool) > (gacB_2_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacB_2_2_bufchan_d;
  logic gacB_2_2_bufchan_r;
  assign gacB_2_2_r = ((! gacB_2_2_bufchan_d[0]) || gacB_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_2_2_bufchan_d <= 1'd0;
    else if (gacB_2_2_r) gacB_2_2_bufchan_d <= gacB_2_2_d;
  MyDTBool_Bool_Bool_t gacB_2_2_bufchan_buf;
  assign gacB_2_2_bufchan_r = (! gacB_2_2_bufchan_buf[0]);
  assign gacB_2_2_argbuf_d = (gacB_2_2_bufchan_buf[0] ? gacB_2_2_bufchan_buf :
                              gacB_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacB_2_2_argbuf_r && gacB_2_2_bufchan_buf[0]))
        gacB_2_2_bufchan_buf <= 1'd0;
      else if (((! gacB_2_2_argbuf_r) && (! gacB_2_2_bufchan_buf[0])))
        gacB_2_2_bufchan_buf <= gacB_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacB_2_destruct,MyDTBool_Bool_Bool) > [(gacB_2_1,MyDTBool_Bool_Bool),
                                                                       (gacB_2_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacB_2_destruct_emitted;
  logic [1:0] gacB_2_destruct_done;
  assign gacB_2_1_d = (gacB_2_destruct_d[0] && (! gacB_2_destruct_emitted[0]));
  assign gacB_2_2_d = (gacB_2_destruct_d[0] && (! gacB_2_destruct_emitted[1]));
  assign gacB_2_destruct_done = (gacB_2_destruct_emitted | ({gacB_2_2_d[0],
                                                             gacB_2_1_d[0]} & {gacB_2_2_r,
                                                                               gacB_2_1_r}));
  assign gacB_2_destruct_r = (& gacB_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_2_destruct_emitted <= 2'd0;
    else
      gacB_2_destruct_emitted <= (gacB_2_destruct_r ? 2'd0 :
                                  gacB_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacB_3_2,MyDTBool_Bool_Bool) > (gacB_3_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacB_3_2_bufchan_d;
  logic gacB_3_2_bufchan_r;
  assign gacB_3_2_r = ((! gacB_3_2_bufchan_d[0]) || gacB_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_3_2_bufchan_d <= 1'd0;
    else if (gacB_3_2_r) gacB_3_2_bufchan_d <= gacB_3_2_d;
  MyDTBool_Bool_Bool_t gacB_3_2_bufchan_buf;
  assign gacB_3_2_bufchan_r = (! gacB_3_2_bufchan_buf[0]);
  assign gacB_3_2_argbuf_d = (gacB_3_2_bufchan_buf[0] ? gacB_3_2_bufchan_buf :
                              gacB_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacB_3_2_argbuf_r && gacB_3_2_bufchan_buf[0]))
        gacB_3_2_bufchan_buf <= 1'd0;
      else if (((! gacB_3_2_argbuf_r) && (! gacB_3_2_bufchan_buf[0])))
        gacB_3_2_bufchan_buf <= gacB_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacB_3_destruct,MyDTBool_Bool_Bool) > [(gacB_3_1,MyDTBool_Bool_Bool),
                                                                       (gacB_3_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacB_3_destruct_emitted;
  logic [1:0] gacB_3_destruct_done;
  assign gacB_3_1_d = (gacB_3_destruct_d[0] && (! gacB_3_destruct_emitted[0]));
  assign gacB_3_2_d = (gacB_3_destruct_d[0] && (! gacB_3_destruct_emitted[1]));
  assign gacB_3_destruct_done = (gacB_3_destruct_emitted | ({gacB_3_2_d[0],
                                                             gacB_3_1_d[0]} & {gacB_3_2_r,
                                                                               gacB_3_1_r}));
  assign gacB_3_destruct_r = (& gacB_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_3_destruct_emitted <= 2'd0;
    else
      gacB_3_destruct_emitted <= (gacB_3_destruct_r ? 2'd0 :
                                  gacB_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacB_4_destruct,MyDTBool_Bool_Bool) > (gacB_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacB_4_destruct_bufchan_d;
  logic gacB_4_destruct_bufchan_r;
  assign gacB_4_destruct_r = ((! gacB_4_destruct_bufchan_d[0]) || gacB_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacB_4_destruct_r)
        gacB_4_destruct_bufchan_d <= gacB_4_destruct_d;
  MyDTBool_Bool_Bool_t gacB_4_destruct_bufchan_buf;
  assign gacB_4_destruct_bufchan_r = (! gacB_4_destruct_bufchan_buf[0]);
  assign gacB_4_1_argbuf_d = (gacB_4_destruct_bufchan_buf[0] ? gacB_4_destruct_bufchan_buf :
                              gacB_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacB_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacB_4_1_argbuf_r && gacB_4_destruct_bufchan_buf[0]))
        gacB_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacB_4_1_argbuf_r) && (! gacB_4_destruct_bufchan_buf[0])))
        gacB_4_destruct_bufchan_buf <= gacB_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacK_2_2,MyDTBool_Bool_Bool) > (gacK_2_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacK_2_2_bufchan_d;
  logic gacK_2_2_bufchan_r;
  assign gacK_2_2_r = ((! gacK_2_2_bufchan_d[0]) || gacK_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_2_2_bufchan_d <= 1'd0;
    else if (gacK_2_2_r) gacK_2_2_bufchan_d <= gacK_2_2_d;
  MyDTBool_Bool_Bool_t gacK_2_2_bufchan_buf;
  assign gacK_2_2_bufchan_r = (! gacK_2_2_bufchan_buf[0]);
  assign gacK_2_2_argbuf_d = (gacK_2_2_bufchan_buf[0] ? gacK_2_2_bufchan_buf :
                              gacK_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacK_2_2_argbuf_r && gacK_2_2_bufchan_buf[0]))
        gacK_2_2_bufchan_buf <= 1'd0;
      else if (((! gacK_2_2_argbuf_r) && (! gacK_2_2_bufchan_buf[0])))
        gacK_2_2_bufchan_buf <= gacK_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacK_2_destruct,MyDTBool_Bool_Bool) > [(gacK_2_1,MyDTBool_Bool_Bool),
                                                                       (gacK_2_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacK_2_destruct_emitted;
  logic [1:0] gacK_2_destruct_done;
  assign gacK_2_1_d = (gacK_2_destruct_d[0] && (! gacK_2_destruct_emitted[0]));
  assign gacK_2_2_d = (gacK_2_destruct_d[0] && (! gacK_2_destruct_emitted[1]));
  assign gacK_2_destruct_done = (gacK_2_destruct_emitted | ({gacK_2_2_d[0],
                                                             gacK_2_1_d[0]} & {gacK_2_2_r,
                                                                               gacK_2_1_r}));
  assign gacK_2_destruct_r = (& gacK_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_2_destruct_emitted <= 2'd0;
    else
      gacK_2_destruct_emitted <= (gacK_2_destruct_r ? 2'd0 :
                                  gacK_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacK_3_2,MyDTBool_Bool_Bool) > (gacK_3_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacK_3_2_bufchan_d;
  logic gacK_3_2_bufchan_r;
  assign gacK_3_2_r = ((! gacK_3_2_bufchan_d[0]) || gacK_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_3_2_bufchan_d <= 1'd0;
    else if (gacK_3_2_r) gacK_3_2_bufchan_d <= gacK_3_2_d;
  MyDTBool_Bool_Bool_t gacK_3_2_bufchan_buf;
  assign gacK_3_2_bufchan_r = (! gacK_3_2_bufchan_buf[0]);
  assign gacK_3_2_argbuf_d = (gacK_3_2_bufchan_buf[0] ? gacK_3_2_bufchan_buf :
                              gacK_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacK_3_2_argbuf_r && gacK_3_2_bufchan_buf[0]))
        gacK_3_2_bufchan_buf <= 1'd0;
      else if (((! gacK_3_2_argbuf_r) && (! gacK_3_2_bufchan_buf[0])))
        gacK_3_2_bufchan_buf <= gacK_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacK_3_destruct,MyDTBool_Bool_Bool) > [(gacK_3_1,MyDTBool_Bool_Bool),
                                                                       (gacK_3_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacK_3_destruct_emitted;
  logic [1:0] gacK_3_destruct_done;
  assign gacK_3_1_d = (gacK_3_destruct_d[0] && (! gacK_3_destruct_emitted[0]));
  assign gacK_3_2_d = (gacK_3_destruct_d[0] && (! gacK_3_destruct_emitted[1]));
  assign gacK_3_destruct_done = (gacK_3_destruct_emitted | ({gacK_3_2_d[0],
                                                             gacK_3_1_d[0]} & {gacK_3_2_r,
                                                                               gacK_3_1_r}));
  assign gacK_3_destruct_r = (& gacK_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_3_destruct_emitted <= 2'd0;
    else
      gacK_3_destruct_emitted <= (gacK_3_destruct_r ? 2'd0 :
                                  gacK_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacK_4_destruct,MyDTBool_Bool_Bool) > (gacK_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacK_4_destruct_bufchan_d;
  logic gacK_4_destruct_bufchan_r;
  assign gacK_4_destruct_r = ((! gacK_4_destruct_bufchan_d[0]) || gacK_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacK_4_destruct_r)
        gacK_4_destruct_bufchan_d <= gacK_4_destruct_d;
  MyDTBool_Bool_Bool_t gacK_4_destruct_bufchan_buf;
  assign gacK_4_destruct_bufchan_r = (! gacK_4_destruct_bufchan_buf[0]);
  assign gacK_4_1_argbuf_d = (gacK_4_destruct_bufchan_buf[0] ? gacK_4_destruct_bufchan_buf :
                              gacK_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacK_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacK_4_1_argbuf_r && gacK_4_destruct_bufchan_buf[0]))
        gacK_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacK_4_1_argbuf_r) && (! gacK_4_destruct_bufchan_buf[0])))
        gacK_4_destruct_bufchan_buf <= gacK_4_destruct_bufchan_d;
  
  /* dcon (Ty MyDTBool_Bool_Bool,
      Dcon Dcon_&&) : [(go_1,Go)] > (go_1Dcon_&&,MyDTBool_Bool_Bool) */
  assign \go_1Dcon_&&_d  = \Dcon_&&_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_&&_r  && \go_1Dcon_&&_d [0])}};
  
  /* fork (Ty C4) : (go_10_goMux_choice,C4) > [(go_10_goMux_choice_1,C4),
                                          (go_10_goMux_choice_2,C4)] */
  logic [1:0] go_10_goMux_choice_emitted;
  logic [1:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[2:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[2:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 2'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 2'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Pointer_QTree_Bool) : (go_10_goMux_choice_1,C4) [(lizzieLet10_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet11_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet12_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet10_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet11_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet12_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet12_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (go_10_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (go_10_goMux_choice_2,C4) [(lizzieLet0_7QNone_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (sc_0_6_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (lizzieLet0_7QVal_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (lizzieLet0_7QError_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (scfarg_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet0_7QNone_Bool_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet0_7QVal_Bool_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet0_7QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet0_7QError_Bool_1_argbuf_r,
          lizzieLet0_7QVal_Bool_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet0_7QNone_Bool_1_argbuf_r} = (go_10_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                                4'd0);
  
  /* fork (Ty C6) : (go_11_goMux_choice,C6) > [(go_11_goMux_choice_1,C6),
                                          (go_11_goMux_choice_2,C6)] */
  logic [1:0] go_11_goMux_choice_emitted;
  logic [1:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 2'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 2'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Bool) : (go_11_goMux_choice_1,C6) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet4_5MQVal_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [5:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet4_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet4_5MQVal_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_11_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTmain_mask_Bool) : (go_11_goMux_choice_2,C6) [(lizzieLet4_6MQNone_1_argbuf,Pointer_CTmain_mask_Bool),
                                                               (sc_0_10_1_argbuf,Pointer_CTmain_mask_Bool),
                                                               (lizzieLet4_6MQVal_1_argbuf,Pointer_CTmain_mask_Bool),
                                                               (lizzieLet4_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTmain_mask_Bool),
                                                               (lizzieLet4_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTmain_mask_Bool),
                                                               (lizzieLet4_4MQNode_4QError_Bool_1_argbuf,Pointer_CTmain_mask_Bool)] > (scfarg_0_1_goMux_mux,Pointer_CTmain_mask_Bool) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [5:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet4_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   sc_0_10_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet4_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_d};
      3'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet4_4MQNode_4QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet4_4MQNode_4QError_Bool_1_argbuf_r,
          lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_r,
          lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_r,
          lizzieLet4_6MQVal_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet4_6MQNone_1_argbuf_r} = (go_11_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                            6'd0);
  
  /* fork (Ty C5) : (go_12_goMux_choice,C5) > [(go_12_goMux_choice_1,C5),
                                          (go_12_goMux_choice_2,C5)] */
  logic [1:0] go_12_goMux_choice_emitted;
  logic [1:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 2'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 2'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_12_goMux_choice_1,C5) [(lizzieLet5_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [4:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet5_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet6_1_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet7_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet8_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0])};
  assign go_12_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = (go_12_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (go_12_goMux_choice_2,C5) [(lizzieLet11_1_6QNone_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (sc_0_14_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (es_0_1_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (es_0_1_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (lizzieLet11_1_6QError_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (scfarg_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [4:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet11_1_6QNone_Bool_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   sc_0_14_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   es_0_1_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   es_0_1_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet11_1_6QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0])};
  assign go_12_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet11_1_6QError_Bool_1_argbuf_r,
          es_0_1_2MyTrue_1_argbuf_r,
          es_0_1_2MyFalse_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet11_1_6QNone_Bool_1_argbuf_r} = (go_12_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                   5'd0);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (go_1Dcon_&&,MyDTBool_Bool_Bool) > (es_3_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \go_1Dcon_&&_bufchan_d ;
  logic \go_1Dcon_&&_bufchan_r ;
  assign \go_1Dcon_&&_r  = ((! \go_1Dcon_&&_bufchan_d [0]) || \go_1Dcon_&&_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_&&_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_&&_r ) \go_1Dcon_&&_bufchan_d  <= \go_1Dcon_&&_d ;
  MyDTBool_Bool_Bool_t \go_1Dcon_&&_bufchan_buf ;
  assign \go_1Dcon_&&_bufchan_r  = (! \go_1Dcon_&&_bufchan_buf [0]);
  assign es_3_1_argbuf_d = (\go_1Dcon_&&_bufchan_buf [0] ? \go_1Dcon_&&_bufchan_buf  :
                            \go_1Dcon_&&_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_&&_bufchan_buf  <= 1'd0;
    else
      if ((es_3_1_argbuf_r && \go_1Dcon_&&_bufchan_buf [0]))
        \go_1Dcon_&&_bufchan_buf  <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! \go_1Dcon_&&_bufchan_buf [0])))
        \go_1Dcon_&&_bufchan_buf  <= \go_1Dcon_&&_bufchan_d ;
  
  /* dcon (Ty MyDTBool_Bool,
      Dcon Dcon_main1) : [(go_2,Go)] > (go_2Dcon_main1,MyDTBool_Bool) */
  assign go_2Dcon_main1_d = Dcon_main1_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_main1_r && go_2Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTBool_Bool) : (go_2Dcon_main1,MyDTBool_Bool) > (es_2_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t go_2Dcon_main1_bufchan_d;
  logic go_2Dcon_main1_bufchan_r;
  assign go_2Dcon_main1_r = ((! go_2Dcon_main1_bufchan_d[0]) || go_2Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_main1_r) go_2Dcon_main1_bufchan_d <= go_2Dcon_main1_d;
  MyDTBool_Bool_t go_2Dcon_main1_bufchan_buf;
  assign go_2Dcon_main1_bufchan_r = (! go_2Dcon_main1_bufchan_buf[0]);
  assign es_2_1_argbuf_d = (go_2Dcon_main1_bufchan_buf[0] ? go_2Dcon_main1_bufchan_buf :
                            go_2Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_argbuf_r && go_2Dcon_main1_bufchan_buf[0]))
        go_2Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_2_1_argbuf_r) && (! go_2Dcon_main1_bufchan_buf[0])))
        go_2Dcon_main1_bufchan_buf <= go_2Dcon_main1_bufchan_d;
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(go_3_argbuf,Go),
                                                                                                    (es_2_1_argbuf,MyDTBool_Bool),
                                                                                                    (es_3_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                    (m2acT_1,Pointer_QTree_Bool),
                                                                                                    (m3acU_2,Pointer_QTree_Bool)] > (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {go_3_argbuf_d[0],
                                                                                                                                                                                                                        es_2_1_argbuf_d[0],
                                                                                                                                                                                                                        es_3_1_argbuf_d[0],
                                                                                                                                                                                                                        m2acT_1_d[0],
                                                                                                                                                                                                                        m3acU_2_d[0]}), go_3_argbuf_d, es_2_1_argbuf_d, es_3_1_argbuf_d, m2acT_1_d, m3acU_2_d);
  assign {go_3_argbuf_r,
          es_2_1_argbuf_r,
          es_3_1_argbuf_r,
          m2acT_1_r,
          m3acU_2_r} = {5 {(kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0])}};
  
  /* buf (Ty Go) : (go_4,Go) > (go_4_argbuf,Go) */
  Go_t go_4_bufchan_d;
  logic go_4_bufchan_r;
  assign go_4_r = ((! go_4_bufchan_d[0]) || go_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_d <= 1'd0;
    else if (go_4_r) go_4_bufchan_d <= go_4_d;
  Go_t go_4_bufchan_buf;
  assign go_4_bufchan_r = (! go_4_bufchan_buf[0]);
  assign go_4_argbuf_d = (go_4_bufchan_buf[0] ? go_4_bufchan_buf :
                          go_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_buf <= 1'd0;
    else
      if ((go_4_argbuf_r && go_4_bufchan_buf[0]))
        go_4_bufchan_buf <= 1'd0;
      else if (((! go_4_argbuf_r) && (! go_4_bufchan_buf[0])))
        go_4_bufchan_buf <= go_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) : [(go_4_argbuf,Go),
                                                              (es_0_1_argbuf,Pointer_QTree_Bool),
                                                              (m1acS_0,Pointer_MaskQTree)] > (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) */
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d = TupGo___Pointer_QTree_Bool___Pointer_MaskQTree_dc((& {go_4_argbuf_d[0],
                                                                                                                                  es_0_1_argbuf_d[0],
                                                                                                                                  m1acS_0_d[0]}), go_4_argbuf_d, es_0_1_argbuf_d, m1acS_0_d);
  assign {go_4_argbuf_r,
          es_0_1_argbuf_r,
          m1acS_0_r} = {3 {(main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0])}};
  
  /* fork (Ty C5) : (go_4_goMux_choice,C5) > [(go_4_goMux_choice_1,C5),
                                         (go_4_goMux_choice_2,C5),
                                         (go_4_goMux_choice_3,C5),
                                         (go_4_goMux_choice_4,C5),
                                         (go_4_goMux_choice_5,C5)] */
  logic [4:0] go_4_goMux_choice_emitted;
  logic [4:0] go_4_goMux_choice_done;
  assign go_4_goMux_choice_1_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[0]))};
  assign go_4_goMux_choice_2_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[1]))};
  assign go_4_goMux_choice_3_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[2]))};
  assign go_4_goMux_choice_4_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[3]))};
  assign go_4_goMux_choice_5_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[4]))};
  assign go_4_goMux_choice_done = (go_4_goMux_choice_emitted | ({go_4_goMux_choice_5_d[0],
                                                                 go_4_goMux_choice_4_d[0],
                                                                 go_4_goMux_choice_3_d[0],
                                                                 go_4_goMux_choice_2_d[0],
                                                                 go_4_goMux_choice_1_d[0]} & {go_4_goMux_choice_5_r,
                                                                                              go_4_goMux_choice_4_r,
                                                                                              go_4_goMux_choice_3_r,
                                                                                              go_4_goMux_choice_2_r,
                                                                                              go_4_goMux_choice_1_r}));
  assign go_4_goMux_choice_r = (& go_4_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_goMux_choice_emitted <= 5'd0;
    else
      go_4_goMux_choice_emitted <= (go_4_goMux_choice_r ? 5'd0 :
                                    go_4_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool) : (go_4_goMux_choice_1,C5) [(call_kron_kron_Bool_Bool_Bool_goMux2,MyDTBool_Bool),
                                                   (isZacJ_2_2_argbuf,MyDTBool_Bool),
                                                   (isZacJ_3_2_argbuf,MyDTBool_Bool),
                                                   (isZacJ_4_1_argbuf,MyDTBool_Bool),
                                                   (lizzieLet0_5QNode_Bool_2_argbuf,MyDTBool_Bool)] > (isZacJ_goMux_mux,MyDTBool_Bool) */
  logic [0:0] isZacJ_goMux_mux_mux;
  logic [4:0] isZacJ_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_1_d[3:1])
      3'd0:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Bool_Bool_Bool_goMux2_d};
      3'd1:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd2,
                                                           isZacJ_2_2_argbuf_d};
      3'd2:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd4,
                                                           isZacJ_3_2_argbuf_d};
      3'd3:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd8,
                                                           isZacJ_4_1_argbuf_d};
      3'd4:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd16,
                                                           lizzieLet0_5QNode_Bool_2_argbuf_d};
      default:
        {isZacJ_goMux_mux_onehot, isZacJ_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacJ_goMux_mux_d = (isZacJ_goMux_mux_mux[0] && go_4_goMux_choice_1_d[0]);
  assign go_4_goMux_choice_1_r = (isZacJ_goMux_mux_d[0] && isZacJ_goMux_mux_r);
  assign {lizzieLet0_5QNode_Bool_2_argbuf_r,
          isZacJ_4_1_argbuf_r,
          isZacJ_3_2_argbuf_r,
          isZacJ_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux2_r} = (go_4_goMux_choice_1_r ? isZacJ_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool_Bool) : (go_4_goMux_choice_2,C5) [(call_kron_kron_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool),
                                                        (gacK_2_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacK_3_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacK_4_1_argbuf,MyDTBool_Bool_Bool),
                                                        (lizzieLet0_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool)] > (gacK_goMux_mux,MyDTBool_Bool_Bool) */
  logic [0:0] gacK_goMux_mux_mux;
  logic [4:0] gacK_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_2_d[3:1])
      3'd0:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Bool_Bool_Bool_goMux3_d};
      3'd1:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd2,
                                                       gacK_2_2_argbuf_d};
      3'd2:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd4,
                                                       gacK_3_2_argbuf_d};
      3'd3:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd8,
                                                       gacK_4_1_argbuf_d};
      3'd4:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd16,
                                                       lizzieLet0_3QNode_Bool_2_argbuf_d};
      default:
        {gacK_goMux_mux_onehot, gacK_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacK_goMux_mux_d = (gacK_goMux_mux_mux[0] && go_4_goMux_choice_2_d[0]);
  assign go_4_goMux_choice_2_r = (gacK_goMux_mux_d[0] && gacK_goMux_mux_r);
  assign {lizzieLet0_3QNode_Bool_2_argbuf_r,
          gacK_4_1_argbuf_r,
          gacK_3_2_argbuf_r,
          gacK_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux3_r} = (go_4_goMux_choice_2_r ? gacK_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_4_goMux_choice_3,C5) [(call_kron_kron_Bool_Bool_Bool_goMux4,Pointer_QTree_Bool),
                                                        (q3acQ_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2acP_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1acO_3_1_argbuf,Pointer_QTree_Bool),
                                                        (q4acR_1_argbuf,Pointer_QTree_Bool)] > (m1acL_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m1acL_goMux_mux_mux;
  logic [4:0] m1acL_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_3_d[3:1])
      3'd0:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Bool_Bool_Bool_goMux4_d};
      3'd1:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd2,
                                                         q3acQ_1_1_argbuf_d};
      3'd2:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd4,
                                                         q2acP_2_1_argbuf_d};
      3'd3:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd8,
                                                         q1acO_3_1_argbuf_d};
      3'd4:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd16,
                                                         q4acR_1_argbuf_d};
      default:
        {m1acL_goMux_mux_onehot, m1acL_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1acL_goMux_mux_d = {m1acL_goMux_mux_mux[16:1],
                              (m1acL_goMux_mux_mux[0] && go_4_goMux_choice_3_d[0])};
  assign go_4_goMux_choice_3_r = (m1acL_goMux_mux_d[0] && m1acL_goMux_mux_r);
  assign {q4acR_1_argbuf_r,
          q1acO_3_1_argbuf_r,
          q2acP_2_1_argbuf_r,
          q3acQ_1_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux4_r} = (go_4_goMux_choice_3_r ? m1acL_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_4_goMux_choice_4,C5) [(call_kron_kron_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool),
                                                        (m2acM_2_2_argbuf,Pointer_QTree_Bool),
                                                        (m2acM_3_2_argbuf,Pointer_QTree_Bool),
                                                        (m2acM_4_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet0_6QNode_Bool_2_argbuf,Pointer_QTree_Bool)] > (m2acM_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m2acM_goMux_mux_mux;
  logic [4:0] m2acM_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_4_d[3:1])
      3'd0:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Bool_Bool_Bool_goMux5_d};
      3'd1:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd2,
                                                         m2acM_2_2_argbuf_d};
      3'd2:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd4,
                                                         m2acM_3_2_argbuf_d};
      3'd3:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd8,
                                                         m2acM_4_1_argbuf_d};
      3'd4:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd16,
                                                         lizzieLet0_6QNode_Bool_2_argbuf_d};
      default:
        {m2acM_goMux_mux_onehot, m2acM_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2acM_goMux_mux_d = {m2acM_goMux_mux_mux[16:1],
                              (m2acM_goMux_mux_mux[0] && go_4_goMux_choice_4_d[0])};
  assign go_4_goMux_choice_4_r = (m2acM_goMux_mux_d[0] && m2acM_goMux_mux_r);
  assign {lizzieLet0_6QNode_Bool_2_argbuf_r,
          m2acM_4_1_argbuf_r,
          m2acM_3_2_argbuf_r,
          m2acM_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux5_r} = (go_4_goMux_choice_4_r ? m2acM_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (go_4_goMux_choice_5,C5) [(call_kron_kron_Bool_Bool_Bool_goMux6,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca3_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (sc_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Bool_Bool_Bool_goMux6_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_4_goMux_choice_5_d[0])};
  assign go_4_goMux_choice_5_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux6_r} = (go_4_goMux_choice_5_r ? sc_0_goMux_mux_onehot :
                                                     5'd0);
  
  /* fork (Ty C5) : (go_5_goMux_choice,C5) > [(go_5_goMux_choice_1,C5),
                                         (go_5_goMux_choice_2,C5),
                                         (go_5_goMux_choice_3,C5)] */
  logic [2:0] go_5_goMux_choice_emitted;
  logic [2:0] go_5_goMux_choice_done;
  assign go_5_goMux_choice_1_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[0]))};
  assign go_5_goMux_choice_2_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[1]))};
  assign go_5_goMux_choice_3_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[2]))};
  assign go_5_goMux_choice_done = (go_5_goMux_choice_emitted | ({go_5_goMux_choice_3_d[0],
                                                                 go_5_goMux_choice_2_d[0],
                                                                 go_5_goMux_choice_1_d[0]} & {go_5_goMux_choice_3_r,
                                                                                              go_5_goMux_choice_2_r,
                                                                                              go_5_goMux_choice_1_r}));
  assign go_5_goMux_choice_r = (& go_5_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_goMux_choice_emitted <= 3'd0;
    else
      go_5_goMux_choice_emitted <= (go_5_goMux_choice_r ? 3'd0 :
                                    go_5_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_5_goMux_choice_1,C5) [(call_main_mask_Bool_goMux2,Pointer_QTree_Bool),
                                                        (t3acr_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2acq_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1acp_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4acs_1_argbuf,Pointer_QTree_Bool)] > (maci_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] maci_goMux_mux_mux;
  logic [4:0] maci_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_1_d[3:1])
      3'd0:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd1,
                                                       call_main_mask_Bool_goMux2_d};
      3'd1:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd2,
                                                       t3acr_1_1_argbuf_d};
      3'd2:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd4,
                                                       t2acq_2_1_argbuf_d};
      3'd3:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd8,
                                                       t1acp_3_1_argbuf_d};
      3'd4:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd16,
                                                       t4acs_1_argbuf_d};
      default:
        {maci_goMux_mux_onehot, maci_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign maci_goMux_mux_d = {maci_goMux_mux_mux[16:1],
                             (maci_goMux_mux_mux[0] && go_5_goMux_choice_1_d[0])};
  assign go_5_goMux_choice_1_r = (maci_goMux_mux_d[0] && maci_goMux_mux_r);
  assign {t4acs_1_argbuf_r,
          t1acp_3_1_argbuf_r,
          t2acq_2_1_argbuf_r,
          t3acr_1_1_argbuf_r,
          call_main_mask_Bool_goMux2_r} = (go_5_goMux_choice_1_r ? maci_goMux_mux_onehot :
                                           5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_5_goMux_choice_2,C5) [(call_main_mask_Bool_goMux3,Pointer_MaskQTree),
                                                       (q3acm_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2acl_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1ack_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet4_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree)] > (mskacj_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] mskacj_goMux_mux_mux;
  logic [4:0] mskacj_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_2_d[3:1])
      3'd0:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Bool_goMux3_d};
      3'd1:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd2,
                                                           q3acm_1_1_argbuf_d};
      3'd2:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd4,
                                                           q2acl_2_1_argbuf_d};
      3'd3:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd8,
                                                           q1ack_3_1_argbuf_d};
      3'd4:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd16,
                                                           lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_d};
      default:
        {mskacj_goMux_mux_onehot, mskacj_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign mskacj_goMux_mux_d = {mskacj_goMux_mux_mux[16:1],
                               (mskacj_goMux_mux_mux[0] && go_5_goMux_choice_2_d[0])};
  assign go_5_goMux_choice_2_r = (mskacj_goMux_mux_d[0] && mskacj_goMux_mux_r);
  assign {lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_r,
          q1ack_3_1_argbuf_r,
          q2acl_2_1_argbuf_r,
          q3acm_1_1_argbuf_r,
          call_main_mask_Bool_goMux3_r} = (go_5_goMux_choice_2_r ? mskacj_goMux_mux_onehot :
                                           5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_mask_Bool) : (go_5_goMux_choice_3,C5) [(call_main_mask_Bool_goMux4,Pointer_CTmain_mask_Bool),
                                                              (sca2_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca1_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca0_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca3_1_1_argbuf,Pointer_CTmain_mask_Bool)] > (sc_0_1_goMux_mux,Pointer_CTmain_mask_Bool) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Bool_goMux4_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_5_goMux_choice_3_d[0])};
  assign go_5_goMux_choice_3_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_main_mask_Bool_goMux4_r} = (go_5_goMux_choice_3_r ? sc_0_1_goMux_mux_onehot :
                                           5'd0);
  
  /* fork (Ty C5) : (go_6_goMux_choice,C5) > [(go_6_goMux_choice_1,C5),
                                         (go_6_goMux_choice_2,C5),
                                         (go_6_goMux_choice_3,C5),
                                         (go_6_goMux_choice_4,C5),
                                         (go_6_goMux_choice_5,C5)] */
  logic [4:0] go_6_goMux_choice_emitted;
  logic [4:0] go_6_goMux_choice_done;
  assign go_6_goMux_choice_1_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[0]))};
  assign go_6_goMux_choice_2_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[1]))};
  assign go_6_goMux_choice_3_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[2]))};
  assign go_6_goMux_choice_4_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[3]))};
  assign go_6_goMux_choice_5_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[4]))};
  assign go_6_goMux_choice_done = (go_6_goMux_choice_emitted | ({go_6_goMux_choice_5_d[0],
                                                                 go_6_goMux_choice_4_d[0],
                                                                 go_6_goMux_choice_3_d[0],
                                                                 go_6_goMux_choice_2_d[0],
                                                                 go_6_goMux_choice_1_d[0]} & {go_6_goMux_choice_5_r,
                                                                                              go_6_goMux_choice_4_r,
                                                                                              go_6_goMux_choice_3_r,
                                                                                              go_6_goMux_choice_2_r,
                                                                                              go_6_goMux_choice_1_r}));
  assign go_6_goMux_choice_r = (& go_6_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_goMux_choice_emitted <= 5'd0;
    else
      go_6_goMux_choice_emitted <= (go_6_goMux_choice_r ? 5'd0 :
                                    go_6_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool) : (go_6_goMux_choice_1,C5) [(call_map''_map''_Bool_Bool_Bool_goMux2,MyDTBool_Bool),
                                                   (isZacA_2_2_argbuf,MyDTBool_Bool),
                                                   (isZacA_3_2_argbuf,MyDTBool_Bool),
                                                   (isZacA_4_1_argbuf,MyDTBool_Bool),
                                                   (lizzieLet11_1_5QNode_Bool_2_argbuf,MyDTBool_Bool)] > (isZacA_goMux_mux,MyDTBool_Bool) */
  logic [0:0] isZacA_goMux_mux_mux;
  logic [4:0] isZacA_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_1_d[3:1])
      3'd0:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Bool_Bool_Bool_goMux2_d };
      3'd1:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd2,
                                                           isZacA_2_2_argbuf_d};
      3'd2:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd4,
                                                           isZacA_3_2_argbuf_d};
      3'd3:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd8,
                                                           isZacA_4_1_argbuf_d};
      3'd4:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd16,
                                                           lizzieLet11_1_5QNode_Bool_2_argbuf_d};
      default:
        {isZacA_goMux_mux_onehot, isZacA_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacA_goMux_mux_d = (isZacA_goMux_mux_mux[0] && go_6_goMux_choice_1_d[0]);
  assign go_6_goMux_choice_1_r = (isZacA_goMux_mux_d[0] && isZacA_goMux_mux_r);
  assign {lizzieLet11_1_5QNode_Bool_2_argbuf_r,
          isZacA_4_1_argbuf_r,
          isZacA_3_2_argbuf_r,
          isZacA_2_2_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux2_r } = (go_6_goMux_choice_1_r ? isZacA_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool_Bool) : (go_6_goMux_choice_2,C5) [(call_map''_map''_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool),
                                                        (gacB_2_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacB_3_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacB_4_1_argbuf,MyDTBool_Bool_Bool),
                                                        (lizzieLet11_1_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool)] > (gacB_goMux_mux,MyDTBool_Bool_Bool) */
  logic [0:0] gacB_goMux_mux_mux;
  logic [4:0] gacB_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_2_d[3:1])
      3'd0:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Bool_Bool_Bool_goMux3_d };
      3'd1:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd2,
                                                       gacB_2_2_argbuf_d};
      3'd2:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd4,
                                                       gacB_3_2_argbuf_d};
      3'd3:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd8,
                                                       gacB_4_1_argbuf_d};
      3'd4:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd16,
                                                       lizzieLet11_1_3QNode_Bool_2_argbuf_d};
      default:
        {gacB_goMux_mux_onehot, gacB_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacB_goMux_mux_d = (gacB_goMux_mux_mux[0] && go_6_goMux_choice_2_d[0]);
  assign go_6_goMux_choice_2_r = (gacB_goMux_mux_d[0] && gacB_goMux_mux_r);
  assign {lizzieLet11_1_3QNode_Bool_2_argbuf_r,
          gacB_4_1_argbuf_r,
          gacB_3_2_argbuf_r,
          gacB_2_2_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux3_r } = (go_6_goMux_choice_2_r ? gacB_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty MyBool) : (go_6_goMux_choice_3,C5) [(call_map''_map''_Bool_Bool_Bool_goMux4,MyBool),
                                            (v'acC_2_2_argbuf,MyBool),
                                            (v'acC_3_2_argbuf,MyBool),
                                            (v'acC_4_1_argbuf,MyBool),
                                            (lizzieLet11_1_7QNode_Bool_2_argbuf,MyBool)] > (v'acC_goMux_mux,MyBool) */
  logic [1:0] \v'acC_goMux_mux_mux ;
  logic [4:0] \v'acC_goMux_mux_onehot ;
  always_comb
    unique case (go_6_goMux_choice_3_d[3:1])
      3'd0:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd1,
                                                             \call_map''_map''_Bool_Bool_Bool_goMux4_d };
      3'd1:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd2,
                                                             \v'acC_2_2_argbuf_d };
      3'd2:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd4,
                                                             \v'acC_3_2_argbuf_d };
      3'd3:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd8,
                                                             \v'acC_4_1_argbuf_d };
      3'd4:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd16,
                                                             lizzieLet11_1_7QNode_Bool_2_argbuf_d};
      default:
        {\v'acC_goMux_mux_onehot , \v'acC_goMux_mux_mux } = {5'd0,
                                                             {1'd0, 1'd0}};
    endcase
  assign \v'acC_goMux_mux_d  = {\v'acC_goMux_mux_mux [1:1],
                                (\v'acC_goMux_mux_mux [0] && go_6_goMux_choice_3_d[0])};
  assign go_6_goMux_choice_3_r = (\v'acC_goMux_mux_d [0] && \v'acC_goMux_mux_r );
  assign {lizzieLet11_1_7QNode_Bool_2_argbuf_r,
          \v'acC_4_1_argbuf_r ,
          \v'acC_3_2_argbuf_r ,
          \v'acC_2_2_argbuf_r ,
          \call_map''_map''_Bool_Bool_Bool_goMux4_r } = (go_6_goMux_choice_3_r ? \v'acC_goMux_mux_onehot  :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_6_goMux_choice_4,C5) [(call_map''_map''_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool),
                                                        (q3acH_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2acG_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1acF_3_1_argbuf,Pointer_QTree_Bool),
                                                        (q4acI_1_argbuf,Pointer_QTree_Bool)] > (macD_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] macD_goMux_mux_mux;
  logic [4:0] macD_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_4_d[3:1])
      3'd0:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Bool_Bool_Bool_goMux5_d };
      3'd1:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd2,
                                                       q3acH_1_1_argbuf_d};
      3'd2:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd4,
                                                       q2acG_2_1_argbuf_d};
      3'd3:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd8,
                                                       q1acF_3_1_argbuf_d};
      3'd4:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd16,
                                                       q4acI_1_argbuf_d};
      default:
        {macD_goMux_mux_onehot, macD_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign macD_goMux_mux_d = {macD_goMux_mux_mux[16:1],
                             (macD_goMux_mux_mux[0] && go_6_goMux_choice_4_d[0])};
  assign go_6_goMux_choice_4_r = (macD_goMux_mux_d[0] && macD_goMux_mux_r);
  assign {q4acI_1_argbuf_r,
          q1acF_3_1_argbuf_r,
          q2acG_2_1_argbuf_r,
          q3acH_1_1_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux5_r } = (go_6_goMux_choice_4_r ? macD_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (go_6_goMux_choice_5,C5) [(call_map''_map''_Bool_Bool_Bool_goMux6,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca2_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca1_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca3_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (sc_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Bool_Bool_Bool_goMux6_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_6_goMux_choice_5_d[0])};
  assign go_6_goMux_choice_5_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux6_r } = (go_6_goMux_choice_5_r ? sc_0_2_goMux_mux_onehot :
                                                         5'd0);
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lkron_kron_Bool_Bool_Boolsbos) : [(go_7_1,Go)] > (go_7_1Lkron_kron_Bool_Bool_Boolsbos,CTkron_kron_Bool_Bool_Bool) */
  assign go_7_1Lkron_kron_Bool_Bool_Boolsbos_d = Lkron_kron_Bool_Bool_Boolsbos_dc((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(go_7_1Lkron_kron_Bool_Bool_Boolsbos_r && go_7_1Lkron_kron_Bool_Bool_Boolsbos_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (go_7_1Lkron_kron_Bool_Bool_Boolsbos,CTkron_kron_Bool_Bool_Bool) > (lizzieLet17_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d;
  logic go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r;
  assign go_7_1Lkron_kron_Bool_Bool_Boolsbos_r = ((! go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d[0]) || go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d <= {83'd0, 1'd0};
    else
      if (go_7_1Lkron_kron_Bool_Bool_Boolsbos_r)
        go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d <= go_7_1Lkron_kron_Bool_Bool_Boolsbos_d;
  CTkron_kron_Bool_Bool_Bool_t go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf;
  assign go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r = (! go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0] ? go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf :
                                   go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= {83'd0, 1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0]))
        go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= {83'd0, 1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0])))
        go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= go_7_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_7_2,Go) > (go_7_2_argbuf,Go) */
  Go_t go_7_2_bufchan_d;
  logic go_7_2_bufchan_r;
  assign go_7_2_r = ((! go_7_2_bufchan_d[0]) || go_7_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_d <= 1'd0;
    else if (go_7_2_r) go_7_2_bufchan_d <= go_7_2_d;
  Go_t go_7_2_bufchan_buf;
  assign go_7_2_bufchan_r = (! go_7_2_bufchan_buf[0]);
  assign go_7_2_argbuf_d = (go_7_2_bufchan_buf[0] ? go_7_2_bufchan_buf :
                            go_7_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_buf <= 1'd0;
    else
      if ((go_7_2_argbuf_r && go_7_2_bufchan_buf[0]))
        go_7_2_bufchan_buf <= 1'd0;
      else if (((! go_7_2_argbuf_r) && (! go_7_2_bufchan_buf[0])))
        go_7_2_bufchan_buf <= go_7_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) : [(go_7_2_argbuf,Go),
                                                                                                                                         (isZacJ_1_1_argbuf,MyDTBool_Bool),
                                                                                                                                         (gacK_1_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                                                         (m1acL_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                                         (m2acM_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                                         (lizzieLet13_1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_dc((& {go_7_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       isZacJ_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       gacK_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       m1acL_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       m2acM_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       lizzieLet13_1_1_argbuf_d[0]}), go_7_2_argbuf_d, isZacJ_1_1_argbuf_d, gacK_1_1_argbuf_d, m1acL_1_1_argbuf_d, m2acM_1_1_argbuf_d, lizzieLet13_1_1_argbuf_d);
  assign {go_7_2_argbuf_r,
          isZacJ_1_1_argbuf_r,
          gacK_1_1_argbuf_r,
          m1acL_1_1_argbuf_r,
          m2acM_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r} = {6 {(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0])}};
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lmain_mask_Boolsbos) : [(go_8_1,Go)] > (go_8_1Lmain_mask_Boolsbos,CTmain_mask_Bool) */
  assign go_8_1Lmain_mask_Boolsbos_d = Lmain_mask_Boolsbos_dc((& {go_8_1_d[0]}), go_8_1_d);
  assign {go_8_1_r} = {1 {(go_8_1Lmain_mask_Boolsbos_r && go_8_1Lmain_mask_Boolsbos_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (go_8_1Lmain_mask_Boolsbos,CTmain_mask_Bool) > (lizzieLet18_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t go_8_1Lmain_mask_Boolsbos_bufchan_d;
  logic go_8_1Lmain_mask_Boolsbos_bufchan_r;
  assign go_8_1Lmain_mask_Boolsbos_r = ((! go_8_1Lmain_mask_Boolsbos_bufchan_d[0]) || go_8_1Lmain_mask_Boolsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_8_1Lmain_mask_Boolsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_8_1Lmain_mask_Boolsbos_r)
        go_8_1Lmain_mask_Boolsbos_bufchan_d <= go_8_1Lmain_mask_Boolsbos_d;
  CTmain_mask_Bool_t go_8_1Lmain_mask_Boolsbos_bufchan_buf;
  assign go_8_1Lmain_mask_Boolsbos_bufchan_r = (! go_8_1Lmain_mask_Boolsbos_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (go_8_1Lmain_mask_Boolsbos_bufchan_buf[0] ? go_8_1Lmain_mask_Boolsbos_bufchan_buf :
                                   go_8_1Lmain_mask_Boolsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_8_1Lmain_mask_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && go_8_1Lmain_mask_Boolsbos_bufchan_buf[0]))
        go_8_1Lmain_mask_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! go_8_1Lmain_mask_Boolsbos_bufchan_buf[0])))
        go_8_1Lmain_mask_Boolsbos_bufchan_buf <= go_8_1Lmain_mask_Boolsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_8_2,Go) > (go_8_2_argbuf,Go) */
  Go_t go_8_2_bufchan_d;
  logic go_8_2_bufchan_r;
  assign go_8_2_r = ((! go_8_2_bufchan_d[0]) || go_8_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_d <= 1'd0;
    else if (go_8_2_r) go_8_2_bufchan_d <= go_8_2_d;
  Go_t go_8_2_bufchan_buf;
  assign go_8_2_bufchan_r = (! go_8_2_bufchan_buf[0]);
  assign go_8_2_argbuf_d = (go_8_2_bufchan_buf[0] ? go_8_2_bufchan_buf :
                            go_8_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_buf <= 1'd0;
    else
      if ((go_8_2_argbuf_r && go_8_2_bufchan_buf[0]))
        go_8_2_bufchan_buf <= 1'd0;
      else if (((! go_8_2_argbuf_r) && (! go_8_2_bufchan_buf[0])))
        go_8_2_bufchan_buf <= go_8_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) : [(go_8_2_argbuf,Go),
                                                                                         (maci_1_1_argbuf,Pointer_QTree_Bool),
                                                                                         (mskacj_1_1_argbuf,Pointer_MaskQTree),
                                                                                         (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Bool)] > (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) */
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d = TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_dc((& {go_8_2_argbuf_d[0],
                                                                                                                                                                                             maci_1_1_argbuf_d[0],
                                                                                                                                                                                             mskacj_1_1_argbuf_d[0],
                                                                                                                                                                                             lizzieLet4_1_1_argbuf_d[0]}), go_8_2_argbuf_d, maci_1_1_argbuf_d, mskacj_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_8_2_argbuf_r,
          maci_1_1_argbuf_r,
          mskacj_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {4 {(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0])}};
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lmap''_map''_Bool_Bool_Boolsbos) : [(go_9_1,Go)] > (go_9_1Lmap''_map''_Bool_Bool_Boolsbos,CTmap''_map''_Bool_Bool_Bool) */
  assign \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_d  = \Lmap''_map''_Bool_Bool_Boolsbos_dc ((& {go_9_1_d[0]}), go_9_1_d);
  assign {go_9_1_r} = {1 {(\go_9_1Lmap''_map''_Bool_Bool_Boolsbos_r  && \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (go_9_1Lmap''_map''_Bool_Bool_Boolsbos,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet19_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d ;
  logic \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r ;
  assign \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_r  = ((! \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d [0]) || \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d  <= {68'd0, 1'd0};
    else
      if (\go_9_1Lmap''_map''_Bool_Bool_Boolsbos_r )
        \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d  <= \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf ;
  assign \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r  = (! \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0]);
  assign lizzieLet19_1_argbuf_d = (\go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0] ? \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  :
                                   \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= {68'd0,
                                                              1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0]))
        \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= {68'd0,
                                                                1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0])))
        \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= \go_9_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_9_2,Go) > (go_9_2_argbuf,Go) */
  Go_t go_9_2_bufchan_d;
  logic go_9_2_bufchan_r;
  assign go_9_2_r = ((! go_9_2_bufchan_d[0]) || go_9_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_2_bufchan_d <= 1'd0;
    else if (go_9_2_r) go_9_2_bufchan_d <= go_9_2_d;
  Go_t go_9_2_bufchan_buf;
  assign go_9_2_bufchan_r = (! go_9_2_bufchan_buf[0]);
  assign go_9_2_argbuf_d = (go_9_2_bufchan_buf[0] ? go_9_2_bufchan_buf :
                            go_9_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_2_bufchan_buf <= 1'd0;
    else
      if ((go_9_2_argbuf_r && go_9_2_bufchan_buf[0]))
        go_9_2_bufchan_buf <= 1'd0;
      else if (((! go_9_2_argbuf_r) && (! go_9_2_bufchan_buf[0])))
        go_9_2_bufchan_buf <= go_9_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) : [(go_9_2_argbuf,Go),
                                                                                                                               (isZacA_1_1_argbuf,MyDTBool_Bool),
                                                                                                                               (gacB_1_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                                               (v'acC_1_1_argbuf,MyBool),
                                                                                                                               (macD_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                               (lizzieLet9_1_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d  = \TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_dc ((& {go_9_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                         isZacA_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         gacB_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         \v'acC_1_1_argbuf_d [0],
                                                                                                                                                                                                                                                                                         macD_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         lizzieLet9_1_1_argbuf_d[0]}), go_9_2_argbuf_d, isZacA_1_1_argbuf_d, gacB_1_1_argbuf_d, \v'acC_1_1_argbuf_d , macD_1_1_argbuf_d, lizzieLet9_1_1_argbuf_d);
  assign {go_9_2_argbuf_r,
          isZacA_1_1_argbuf_r,
          gacB_1_1_argbuf_r,
          \v'acC_1_1_argbuf_r ,
          macD_1_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r} = {6 {(\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0])}};
  
  /* buf (Ty MyDTBool_Bool) : (isZacA_2_2,MyDTBool_Bool) > (isZacA_2_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacA_2_2_bufchan_d;
  logic isZacA_2_2_bufchan_r;
  assign isZacA_2_2_r = ((! isZacA_2_2_bufchan_d[0]) || isZacA_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_2_2_bufchan_d <= 1'd0;
    else if (isZacA_2_2_r) isZacA_2_2_bufchan_d <= isZacA_2_2_d;
  MyDTBool_Bool_t isZacA_2_2_bufchan_buf;
  assign isZacA_2_2_bufchan_r = (! isZacA_2_2_bufchan_buf[0]);
  assign isZacA_2_2_argbuf_d = (isZacA_2_2_bufchan_buf[0] ? isZacA_2_2_bufchan_buf :
                                isZacA_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacA_2_2_argbuf_r && isZacA_2_2_bufchan_buf[0]))
        isZacA_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacA_2_2_argbuf_r) && (! isZacA_2_2_bufchan_buf[0])))
        isZacA_2_2_bufchan_buf <= isZacA_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacA_2_destruct,MyDTBool_Bool) > [(isZacA_2_1,MyDTBool_Bool),
                                                               (isZacA_2_2,MyDTBool_Bool)] */
  logic [1:0] isZacA_2_destruct_emitted;
  logic [1:0] isZacA_2_destruct_done;
  assign isZacA_2_1_d = (isZacA_2_destruct_d[0] && (! isZacA_2_destruct_emitted[0]));
  assign isZacA_2_2_d = (isZacA_2_destruct_d[0] && (! isZacA_2_destruct_emitted[1]));
  assign isZacA_2_destruct_done = (isZacA_2_destruct_emitted | ({isZacA_2_2_d[0],
                                                                 isZacA_2_1_d[0]} & {isZacA_2_2_r,
                                                                                     isZacA_2_1_r}));
  assign isZacA_2_destruct_r = (& isZacA_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_2_destruct_emitted <= 2'd0;
    else
      isZacA_2_destruct_emitted <= (isZacA_2_destruct_r ? 2'd0 :
                                    isZacA_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacA_3_2,MyDTBool_Bool) > (isZacA_3_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacA_3_2_bufchan_d;
  logic isZacA_3_2_bufchan_r;
  assign isZacA_3_2_r = ((! isZacA_3_2_bufchan_d[0]) || isZacA_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_3_2_bufchan_d <= 1'd0;
    else if (isZacA_3_2_r) isZacA_3_2_bufchan_d <= isZacA_3_2_d;
  MyDTBool_Bool_t isZacA_3_2_bufchan_buf;
  assign isZacA_3_2_bufchan_r = (! isZacA_3_2_bufchan_buf[0]);
  assign isZacA_3_2_argbuf_d = (isZacA_3_2_bufchan_buf[0] ? isZacA_3_2_bufchan_buf :
                                isZacA_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacA_3_2_argbuf_r && isZacA_3_2_bufchan_buf[0]))
        isZacA_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacA_3_2_argbuf_r) && (! isZacA_3_2_bufchan_buf[0])))
        isZacA_3_2_bufchan_buf <= isZacA_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacA_3_destruct,MyDTBool_Bool) > [(isZacA_3_1,MyDTBool_Bool),
                                                               (isZacA_3_2,MyDTBool_Bool)] */
  logic [1:0] isZacA_3_destruct_emitted;
  logic [1:0] isZacA_3_destruct_done;
  assign isZacA_3_1_d = (isZacA_3_destruct_d[0] && (! isZacA_3_destruct_emitted[0]));
  assign isZacA_3_2_d = (isZacA_3_destruct_d[0] && (! isZacA_3_destruct_emitted[1]));
  assign isZacA_3_destruct_done = (isZacA_3_destruct_emitted | ({isZacA_3_2_d[0],
                                                                 isZacA_3_1_d[0]} & {isZacA_3_2_r,
                                                                                     isZacA_3_1_r}));
  assign isZacA_3_destruct_r = (& isZacA_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_3_destruct_emitted <= 2'd0;
    else
      isZacA_3_destruct_emitted <= (isZacA_3_destruct_r ? 2'd0 :
                                    isZacA_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacA_4_destruct,MyDTBool_Bool) > (isZacA_4_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacA_4_destruct_bufchan_d;
  logic isZacA_4_destruct_bufchan_r;
  assign isZacA_4_destruct_r = ((! isZacA_4_destruct_bufchan_d[0]) || isZacA_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacA_4_destruct_r)
        isZacA_4_destruct_bufchan_d <= isZacA_4_destruct_d;
  MyDTBool_Bool_t isZacA_4_destruct_bufchan_buf;
  assign isZacA_4_destruct_bufchan_r = (! isZacA_4_destruct_bufchan_buf[0]);
  assign isZacA_4_1_argbuf_d = (isZacA_4_destruct_bufchan_buf[0] ? isZacA_4_destruct_bufchan_buf :
                                isZacA_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacA_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacA_4_1_argbuf_r && isZacA_4_destruct_bufchan_buf[0]))
        isZacA_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacA_4_1_argbuf_r) && (! isZacA_4_destruct_bufchan_buf[0])))
        isZacA_4_destruct_bufchan_buf <= isZacA_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (isZacJ_2_2,MyDTBool_Bool) > (isZacJ_2_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacJ_2_2_bufchan_d;
  logic isZacJ_2_2_bufchan_r;
  assign isZacJ_2_2_r = ((! isZacJ_2_2_bufchan_d[0]) || isZacJ_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_2_2_bufchan_d <= 1'd0;
    else if (isZacJ_2_2_r) isZacJ_2_2_bufchan_d <= isZacJ_2_2_d;
  MyDTBool_Bool_t isZacJ_2_2_bufchan_buf;
  assign isZacJ_2_2_bufchan_r = (! isZacJ_2_2_bufchan_buf[0]);
  assign isZacJ_2_2_argbuf_d = (isZacJ_2_2_bufchan_buf[0] ? isZacJ_2_2_bufchan_buf :
                                isZacJ_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacJ_2_2_argbuf_r && isZacJ_2_2_bufchan_buf[0]))
        isZacJ_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacJ_2_2_argbuf_r) && (! isZacJ_2_2_bufchan_buf[0])))
        isZacJ_2_2_bufchan_buf <= isZacJ_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacJ_2_destruct,MyDTBool_Bool) > [(isZacJ_2_1,MyDTBool_Bool),
                                                               (isZacJ_2_2,MyDTBool_Bool)] */
  logic [1:0] isZacJ_2_destruct_emitted;
  logic [1:0] isZacJ_2_destruct_done;
  assign isZacJ_2_1_d = (isZacJ_2_destruct_d[0] && (! isZacJ_2_destruct_emitted[0]));
  assign isZacJ_2_2_d = (isZacJ_2_destruct_d[0] && (! isZacJ_2_destruct_emitted[1]));
  assign isZacJ_2_destruct_done = (isZacJ_2_destruct_emitted | ({isZacJ_2_2_d[0],
                                                                 isZacJ_2_1_d[0]} & {isZacJ_2_2_r,
                                                                                     isZacJ_2_1_r}));
  assign isZacJ_2_destruct_r = (& isZacJ_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_2_destruct_emitted <= 2'd0;
    else
      isZacJ_2_destruct_emitted <= (isZacJ_2_destruct_r ? 2'd0 :
                                    isZacJ_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacJ_3_2,MyDTBool_Bool) > (isZacJ_3_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacJ_3_2_bufchan_d;
  logic isZacJ_3_2_bufchan_r;
  assign isZacJ_3_2_r = ((! isZacJ_3_2_bufchan_d[0]) || isZacJ_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_3_2_bufchan_d <= 1'd0;
    else if (isZacJ_3_2_r) isZacJ_3_2_bufchan_d <= isZacJ_3_2_d;
  MyDTBool_Bool_t isZacJ_3_2_bufchan_buf;
  assign isZacJ_3_2_bufchan_r = (! isZacJ_3_2_bufchan_buf[0]);
  assign isZacJ_3_2_argbuf_d = (isZacJ_3_2_bufchan_buf[0] ? isZacJ_3_2_bufchan_buf :
                                isZacJ_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacJ_3_2_argbuf_r && isZacJ_3_2_bufchan_buf[0]))
        isZacJ_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacJ_3_2_argbuf_r) && (! isZacJ_3_2_bufchan_buf[0])))
        isZacJ_3_2_bufchan_buf <= isZacJ_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacJ_3_destruct,MyDTBool_Bool) > [(isZacJ_3_1,MyDTBool_Bool),
                                                               (isZacJ_3_2,MyDTBool_Bool)] */
  logic [1:0] isZacJ_3_destruct_emitted;
  logic [1:0] isZacJ_3_destruct_done;
  assign isZacJ_3_1_d = (isZacJ_3_destruct_d[0] && (! isZacJ_3_destruct_emitted[0]));
  assign isZacJ_3_2_d = (isZacJ_3_destruct_d[0] && (! isZacJ_3_destruct_emitted[1]));
  assign isZacJ_3_destruct_done = (isZacJ_3_destruct_emitted | ({isZacJ_3_2_d[0],
                                                                 isZacJ_3_1_d[0]} & {isZacJ_3_2_r,
                                                                                     isZacJ_3_1_r}));
  assign isZacJ_3_destruct_r = (& isZacJ_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_3_destruct_emitted <= 2'd0;
    else
      isZacJ_3_destruct_emitted <= (isZacJ_3_destruct_r ? 2'd0 :
                                    isZacJ_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacJ_4_destruct,MyDTBool_Bool) > (isZacJ_4_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacJ_4_destruct_bufchan_d;
  logic isZacJ_4_destruct_bufchan_r;
  assign isZacJ_4_destruct_r = ((! isZacJ_4_destruct_bufchan_d[0]) || isZacJ_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacJ_4_destruct_r)
        isZacJ_4_destruct_bufchan_d <= isZacJ_4_destruct_d;
  MyDTBool_Bool_t isZacJ_4_destruct_bufchan_buf;
  assign isZacJ_4_destruct_bufchan_r = (! isZacJ_4_destruct_bufchan_buf[0]);
  assign isZacJ_4_1_argbuf_d = (isZacJ_4_destruct_bufchan_buf[0] ? isZacJ_4_destruct_bufchan_buf :
                                isZacJ_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacJ_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacJ_4_1_argbuf_r && isZacJ_4_destruct_bufchan_buf[0]))
        isZacJ_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacJ_4_1_argbuf_r) && (! isZacJ_4_destruct_bufchan_buf[0])))
        isZacJ_4_destruct_bufchan_buf <= isZacJ_4_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7,Go),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1,Pointer_QTree_Bool)] */
  logic [4:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted;
  logic [4:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[0]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[1]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[2]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_d = {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[16:1],
                                                                                                                                  (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[3]))};
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_d = {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[32:17],
                                                                                                                                  (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[4]))};
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted | ({kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_d[0]} & {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_r}));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r = (& kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= 5'd0;
    else
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ? 5'd0 :
                                                                                                                                 kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1,MyDTBool_Bool_Bool) > (gacK_1_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_d;
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf[0]);
  assign gacK_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf :
                              kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf <= 1'd0;
    else
      if ((gacK_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf <= 1'd0;
      else if (((! gacK_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolgacK_1_bufchan_d;
  
  /* fork (Ty Go) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7,Go) > [(go_7_1,Go),
                                                                                                                                        (go_7_2,Go)] */
  logic [1:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted;
  logic [1:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_done;
  assign go_7_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted[0]));
  assign go_7_2_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted[1]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_done = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted | ({go_7_2_d[0],
                                                                                                                                                                                                                                                               go_7_1_d[0]} & {go_7_2_r,
                                                                                                                                                                                                                                                                               go_7_1_r}));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_r = (& kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted <= 2'd0;
    else
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_emitted <= (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_r ? 2'd0 :
                                                                                                                                   kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_7_done);
  
  /* buf (Ty MyDTBool_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1,MyDTBool_Bool) > (isZacJ_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_d;
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf[0]);
  assign isZacJ_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf :
                                kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf <= 1'd0;
    else
      if ((isZacJ_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf <= 1'd0;
      else if (((! isZacJ_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZacJ_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1,Pointer_QTree_Bool) > (m1acL_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d <= {16'd0,
                                                                                                                                        1'd0};
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf[0]);
  assign m1acL_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf :
                               kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf <= {16'd0,
                                                                                                                                          1'd0};
    else
      if ((m1acL_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf <= {16'd0,
                                                                                                                                            1'd0};
      else if (((! m1acL_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1acL_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1,Pointer_QTree_Bool) > (m2acM_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d <= {16'd0,
                                                                                                                                        1'd0};
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf[0]);
  assign m2acM_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf :
                               kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf <= {16'd0,
                                                                                                                                          1'd0};
    else
      if ((m2acM_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf <= {16'd0,
                                                                                                                                            1'd0};
      else if (((! m2acM_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2acM_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) > (es_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_bufchan_d;
  logic kron_kron_Bool_Bool_Bool_resbuf_bufchan_r;
  assign kron_kron_Bool_Bool_Bool_resbuf_r = ((! kron_kron_Bool_Bool_Bool_resbuf_bufchan_d[0]) || kron_kron_Bool_Bool_Bool_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_Bool_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (kron_kron_Bool_Bool_Bool_resbuf_r)
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_d <= kron_kron_Bool_Bool_Bool_resbuf_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf;
  assign kron_kron_Bool_Bool_Bool_resbuf_bufchan_r = (! kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0] ? kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf :
                            kron_kron_Bool_Bool_Bool_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0]))
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0])))
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= kron_kron_Bool_Bool_Bool_resbuf_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet0_1QNode_Bool,QTree_Bool) > [(q1acO_destruct,Pointer_QTree_Bool),
                                                                    (q2acP_destruct,Pointer_QTree_Bool),
                                                                    (q3acQ_destruct,Pointer_QTree_Bool),
                                                                    (q4acR_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet0_1QNode_Bool_emitted;
  logic [3:0] lizzieLet0_1QNode_Bool_done;
  assign q1acO_destruct_d = {lizzieLet0_1QNode_Bool_d[18:3],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[0]))};
  assign q2acP_destruct_d = {lizzieLet0_1QNode_Bool_d[34:19],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[1]))};
  assign q3acQ_destruct_d = {lizzieLet0_1QNode_Bool_d[50:35],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[2]))};
  assign q4acR_destruct_d = {lizzieLet0_1QNode_Bool_d[66:51],
                             (lizzieLet0_1QNode_Bool_d[0] && (! lizzieLet0_1QNode_Bool_emitted[3]))};
  assign lizzieLet0_1QNode_Bool_done = (lizzieLet0_1QNode_Bool_emitted | ({q4acR_destruct_d[0],
                                                                           q3acQ_destruct_d[0],
                                                                           q2acP_destruct_d[0],
                                                                           q1acO_destruct_d[0]} & {q4acR_destruct_r,
                                                                                                   q3acQ_destruct_r,
                                                                                                   q2acP_destruct_r,
                                                                                                   q1acO_destruct_r}));
  assign lizzieLet0_1QNode_Bool_r = (& lizzieLet0_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet0_1QNode_Bool_emitted <= (lizzieLet0_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet0_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet0_1QVal_Bool,QTree_Bool) > [(vacN_destruct,MyBool)] */
  assign vacN_destruct_d = {lizzieLet0_1QVal_Bool_d[3:3],
                            lizzieLet0_1QVal_Bool_d[0]};
  assign lizzieLet0_1QVal_Bool_r = vacN_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet0_2,QTree_Bool) (lizzieLet0_1,QTree_Bool) > [(_42,QTree_Bool),
                                                                               (lizzieLet0_1QVal_Bool,QTree_Bool),
                                                                               (lizzieLet0_1QNode_Bool,QTree_Bool),
                                                                               (_41,QTree_Bool)] */
  logic [3:0] lizzieLet0_1_onehotd;
  always_comb
    if ((lizzieLet0_2_d[0] && lizzieLet0_1_d[0]))
      unique case (lizzieLet0_2_d[2:1])
        2'd0: lizzieLet0_1_onehotd = 4'd1;
        2'd1: lizzieLet0_1_onehotd = 4'd2;
        2'd2: lizzieLet0_1_onehotd = 4'd4;
        2'd3: lizzieLet0_1_onehotd = 4'd8;
        default: lizzieLet0_1_onehotd = 4'd0;
      endcase
    else lizzieLet0_1_onehotd = 4'd0;
  assign _42_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[0]};
  assign lizzieLet0_1QVal_Bool_d = {lizzieLet0_1_d[66:1],
                                    lizzieLet0_1_onehotd[1]};
  assign lizzieLet0_1QNode_Bool_d = {lizzieLet0_1_d[66:1],
                                     lizzieLet0_1_onehotd[2]};
  assign _41_d = {lizzieLet0_1_d[66:1], lizzieLet0_1_onehotd[3]};
  assign lizzieLet0_1_r = (| (lizzieLet0_1_onehotd & {_41_r,
                                                      lizzieLet0_1QNode_Bool_r,
                                                      lizzieLet0_1QVal_Bool_r,
                                                      _42_r}));
  assign lizzieLet0_2_r = lizzieLet0_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet0_3,QTree_Bool) (gacK_goMux_mux,MyDTBool_Bool_Bool) > [(_40,MyDTBool_Bool_Bool),
                                                                                                 (lizzieLet0_3QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                 (lizzieLet0_3QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                 (_39,MyDTBool_Bool_Bool)] */
  logic [3:0] gacK_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_3_d[0] && gacK_goMux_mux_d[0]))
      unique case (lizzieLet0_3_d[2:1])
        2'd0: gacK_goMux_mux_onehotd = 4'd1;
        2'd1: gacK_goMux_mux_onehotd = 4'd2;
        2'd2: gacK_goMux_mux_onehotd = 4'd4;
        2'd3: gacK_goMux_mux_onehotd = 4'd8;
        default: gacK_goMux_mux_onehotd = 4'd0;
      endcase
    else gacK_goMux_mux_onehotd = 4'd0;
  assign _40_d = gacK_goMux_mux_onehotd[0];
  assign lizzieLet0_3QVal_Bool_d = gacK_goMux_mux_onehotd[1];
  assign lizzieLet0_3QNode_Bool_d = gacK_goMux_mux_onehotd[2];
  assign _39_d = gacK_goMux_mux_onehotd[3];
  assign gacK_goMux_mux_r = (| (gacK_goMux_mux_onehotd & {_39_r,
                                                          lizzieLet0_3QNode_Bool_r,
                                                          lizzieLet0_3QVal_Bool_r,
                                                          _40_r}));
  assign lizzieLet0_3_r = gacK_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (lizzieLet0_3QNode_Bool,MyDTBool_Bool_Bool) > [(lizzieLet0_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                                              (lizzieLet0_3QNode_Bool_2,MyDTBool_Bool_Bool)] */
  logic [1:0] lizzieLet0_3QNode_Bool_emitted;
  logic [1:0] lizzieLet0_3QNode_Bool_done;
  assign lizzieLet0_3QNode_Bool_1_d = (lizzieLet0_3QNode_Bool_d[0] && (! lizzieLet0_3QNode_Bool_emitted[0]));
  assign lizzieLet0_3QNode_Bool_2_d = (lizzieLet0_3QNode_Bool_d[0] && (! lizzieLet0_3QNode_Bool_emitted[1]));
  assign lizzieLet0_3QNode_Bool_done = (lizzieLet0_3QNode_Bool_emitted | ({lizzieLet0_3QNode_Bool_2_d[0],
                                                                           lizzieLet0_3QNode_Bool_1_d[0]} & {lizzieLet0_3QNode_Bool_2_r,
                                                                                                             lizzieLet0_3QNode_Bool_1_r}));
  assign lizzieLet0_3QNode_Bool_r = (& lizzieLet0_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_3QNode_Bool_emitted <= (lizzieLet0_3QNode_Bool_r ? 2'd0 :
                                         lizzieLet0_3QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet0_3QNode_Bool_2,MyDTBool_Bool_Bool) > (lizzieLet0_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_2_bufchan_d;
  logic lizzieLet0_3QNode_Bool_2_bufchan_r;
  assign lizzieLet0_3QNode_Bool_2_r = ((! lizzieLet0_3QNode_Bool_2_bufchan_d[0]) || lizzieLet0_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3QNode_Bool_2_r)
        lizzieLet0_3QNode_Bool_2_bufchan_d <= lizzieLet0_3QNode_Bool_2_d;
  MyDTBool_Bool_Bool_t lizzieLet0_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_3QNode_Bool_2_bufchan_r = (! lizzieLet0_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_3QNode_Bool_2_argbuf_d = (lizzieLet0_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_3QNode_Bool_2_bufchan_buf :
                                              lizzieLet0_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3QNode_Bool_2_argbuf_r && lizzieLet0_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3QNode_Bool_2_argbuf_r) && (! lizzieLet0_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_3QNode_Bool_2_bufchan_buf <= lizzieLet0_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet0_3QVal_Bool,MyDTBool_Bool_Bool) > (lizzieLet0_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet0_3QVal_Bool_bufchan_d;
  logic lizzieLet0_3QVal_Bool_bufchan_r;
  assign lizzieLet0_3QVal_Bool_r = ((! lizzieLet0_3QVal_Bool_bufchan_d[0]) || lizzieLet0_3QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_3QVal_Bool_r)
        lizzieLet0_3QVal_Bool_bufchan_d <= lizzieLet0_3QVal_Bool_d;
  MyDTBool_Bool_Bool_t lizzieLet0_3QVal_Bool_bufchan_buf;
  assign lizzieLet0_3QVal_Bool_bufchan_r = (! lizzieLet0_3QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_3QVal_Bool_1_argbuf_d = (lizzieLet0_3QVal_Bool_bufchan_buf[0] ? lizzieLet0_3QVal_Bool_bufchan_buf :
                                             lizzieLet0_3QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_3QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_3QVal_Bool_1_argbuf_r && lizzieLet0_3QVal_Bool_bufchan_buf[0]))
        lizzieLet0_3QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_3QVal_Bool_1_argbuf_r) && (! lizzieLet0_3QVal_Bool_bufchan_buf[0])))
        lizzieLet0_3QVal_Bool_bufchan_buf <= lizzieLet0_3QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet0_4,QTree_Bool) (go_4_goMux_data,Go) > [(lizzieLet0_4QNone_Bool,Go),
                                                                  (lizzieLet0_4QVal_Bool,Go),
                                                                  (lizzieLet0_4QNode_Bool,Go),
                                                                  (lizzieLet0_4QError_Bool,Go)] */
  logic [3:0] go_4_goMux_data_onehotd;
  always_comb
    if ((lizzieLet0_4_d[0] && go_4_goMux_data_d[0]))
      unique case (lizzieLet0_4_d[2:1])
        2'd0: go_4_goMux_data_onehotd = 4'd1;
        2'd1: go_4_goMux_data_onehotd = 4'd2;
        2'd2: go_4_goMux_data_onehotd = 4'd4;
        2'd3: go_4_goMux_data_onehotd = 4'd8;
        default: go_4_goMux_data_onehotd = 4'd0;
      endcase
    else go_4_goMux_data_onehotd = 4'd0;
  assign lizzieLet0_4QNone_Bool_d = go_4_goMux_data_onehotd[0];
  assign lizzieLet0_4QVal_Bool_d = go_4_goMux_data_onehotd[1];
  assign lizzieLet0_4QNode_Bool_d = go_4_goMux_data_onehotd[2];
  assign lizzieLet0_4QError_Bool_d = go_4_goMux_data_onehotd[3];
  assign go_4_goMux_data_r = (| (go_4_goMux_data_onehotd & {lizzieLet0_4QError_Bool_r,
                                                            lizzieLet0_4QNode_Bool_r,
                                                            lizzieLet0_4QVal_Bool_r,
                                                            lizzieLet0_4QNone_Bool_r}));
  assign lizzieLet0_4_r = go_4_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet0_4QError_Bool,Go) > [(lizzieLet0_4QError_Bool_1,Go),
                                               (lizzieLet0_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QError_Bool_emitted;
  logic [1:0] lizzieLet0_4QError_Bool_done;
  assign lizzieLet0_4QError_Bool_1_d = (lizzieLet0_4QError_Bool_d[0] && (! lizzieLet0_4QError_Bool_emitted[0]));
  assign lizzieLet0_4QError_Bool_2_d = (lizzieLet0_4QError_Bool_d[0] && (! lizzieLet0_4QError_Bool_emitted[1]));
  assign lizzieLet0_4QError_Bool_done = (lizzieLet0_4QError_Bool_emitted | ({lizzieLet0_4QError_Bool_2_d[0],
                                                                             lizzieLet0_4QError_Bool_1_d[0]} & {lizzieLet0_4QError_Bool_2_r,
                                                                                                                lizzieLet0_4QError_Bool_1_r}));
  assign lizzieLet0_4QError_Bool_r = (& lizzieLet0_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QError_Bool_emitted <= (lizzieLet0_4QError_Bool_r ? 2'd0 :
                                          lizzieLet0_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet0_4QError_Bool_1,Go)] > (lizzieLet0_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet0_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet0_4QError_Bool_1_d[0]}), lizzieLet0_4QError_Bool_1_d);
  assign {lizzieLet0_4QError_Bool_1_r} = {1 {(lizzieLet0_4QError_Bool_1QError_Bool_r && lizzieLet0_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet3_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet0_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet0_4QError_Bool_1QError_Bool_r = ((! lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet0_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_4QError_Bool_1QError_Bool_r)
        lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet0_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet0_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet3_1_argbuf_d = (lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet3_1_argbuf_r && lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet3_1_argbuf_r) && (! lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet0_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet0_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QError_Bool_2,Go) > (lizzieLet0_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QError_Bool_2_bufchan_d;
  logic lizzieLet0_4QError_Bool_2_bufchan_r;
  assign lizzieLet0_4QError_Bool_2_r = ((! lizzieLet0_4QError_Bool_2_bufchan_d[0]) || lizzieLet0_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QError_Bool_2_r)
        lizzieLet0_4QError_Bool_2_bufchan_d <= lizzieLet0_4QError_Bool_2_d;
  Go_t lizzieLet0_4QError_Bool_2_bufchan_buf;
  assign lizzieLet0_4QError_Bool_2_bufchan_r = (! lizzieLet0_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QError_Bool_2_argbuf_d = (lizzieLet0_4QError_Bool_2_bufchan_buf[0] ? lizzieLet0_4QError_Bool_2_bufchan_buf :
                                               lizzieLet0_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QError_Bool_2_argbuf_r && lizzieLet0_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QError_Bool_2_argbuf_r) && (! lizzieLet0_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QError_Bool_2_bufchan_buf <= lizzieLet0_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNode_Bool,Go) > (lizzieLet0_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QNode_Bool_bufchan_d;
  logic lizzieLet0_4QNode_Bool_bufchan_r;
  assign lizzieLet0_4QNode_Bool_r = ((! lizzieLet0_4QNode_Bool_bufchan_d[0]) || lizzieLet0_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNode_Bool_r)
        lizzieLet0_4QNode_Bool_bufchan_d <= lizzieLet0_4QNode_Bool_d;
  Go_t lizzieLet0_4QNode_Bool_bufchan_buf;
  assign lizzieLet0_4QNode_Bool_bufchan_r = (! lizzieLet0_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet0_4QNode_Bool_1_argbuf_d = (lizzieLet0_4QNode_Bool_bufchan_buf[0] ? lizzieLet0_4QNode_Bool_bufchan_buf :
                                              lizzieLet0_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNode_Bool_1_argbuf_r && lizzieLet0_4QNode_Bool_bufchan_buf[0]))
        lizzieLet0_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNode_Bool_1_argbuf_r) && (! lizzieLet0_4QNode_Bool_bufchan_buf[0])))
        lizzieLet0_4QNode_Bool_bufchan_buf <= lizzieLet0_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet0_4QNone_Bool,Go) > [(lizzieLet0_4QNone_Bool_1,Go),
                                              (lizzieLet0_4QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QNone_Bool_emitted;
  logic [1:0] lizzieLet0_4QNone_Bool_done;
  assign lizzieLet0_4QNone_Bool_1_d = (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[0]));
  assign lizzieLet0_4QNone_Bool_2_d = (lizzieLet0_4QNone_Bool_d[0] && (! lizzieLet0_4QNone_Bool_emitted[1]));
  assign lizzieLet0_4QNone_Bool_done = (lizzieLet0_4QNone_Bool_emitted | ({lizzieLet0_4QNone_Bool_2_d[0],
                                                                           lizzieLet0_4QNone_Bool_1_d[0]} & {lizzieLet0_4QNone_Bool_2_r,
                                                                                                             lizzieLet0_4QNone_Bool_1_r}));
  assign lizzieLet0_4QNone_Bool_r = (& lizzieLet0_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_emitted <= (lizzieLet0_4QNone_Bool_r ? 2'd0 :
                                         lizzieLet0_4QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet0_4QNone_Bool_1,Go)] > (lizzieLet0_4QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet0_4QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet0_4QNone_Bool_1_d[0]}), lizzieLet0_4QNone_Bool_1_d);
  assign {lizzieLet0_4QNone_Bool_1_r} = {1 {(lizzieLet0_4QNone_Bool_1QNone_Bool_r && lizzieLet0_4QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_4QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet0_4QNone_Bool_1QNone_Bool_r = ((! lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_4QNone_Bool_1QNone_Bool_r)
        lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet0_4QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_1_argbuf_d = (lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf :
                                  lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet1_1_argbuf_r && lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet1_1_argbuf_r) && (! lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet0_4QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet0_4QNone_Bool_2,Go) > (lizzieLet0_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QNone_Bool_2_bufchan_d;
  logic lizzieLet0_4QNone_Bool_2_bufchan_r;
  assign lizzieLet0_4QNone_Bool_2_r = ((! lizzieLet0_4QNone_Bool_2_bufchan_d[0]) || lizzieLet0_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QNone_Bool_2_r)
        lizzieLet0_4QNone_Bool_2_bufchan_d <= lizzieLet0_4QNone_Bool_2_d;
  Go_t lizzieLet0_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet0_4QNone_Bool_2_bufchan_r = (! lizzieLet0_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QNone_Bool_2_argbuf_d = (lizzieLet0_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet0_4QNone_Bool_2_bufchan_buf :
                                              lizzieLet0_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QNone_Bool_2_argbuf_r && lizzieLet0_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QNone_Bool_2_argbuf_r) && (! lizzieLet0_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QNone_Bool_2_bufchan_buf <= lizzieLet0_4QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet0_4QNone_Bool_2_argbuf,Go),
                           (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf,Go),
                           (lizzieLet0_4QVal_Bool_2_argbuf,Go),
                           (lizzieLet0_4QError_Bool_2_argbuf,Go)] > (go_10_goMux_choice,C4) (go_10_goMux_data,Go) */
  logic [3:0] lizzieLet0_4QNone_Bool_2_argbuf_select_d;
  assign lizzieLet0_4QNone_Bool_2_argbuf_select_d = ((| lizzieLet0_4QNone_Bool_2_argbuf_select_q) ? lizzieLet0_4QNone_Bool_2_argbuf_select_q :
                                                     (lizzieLet0_4QNone_Bool_2_argbuf_d[0] ? 4'd1 :
                                                      (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d[0] ? 4'd2 :
                                                       (lizzieLet0_4QVal_Bool_2_argbuf_d[0] ? 4'd4 :
                                                        (lizzieLet0_4QError_Bool_2_argbuf_d[0] ? 4'd8 :
                                                         4'd0)))));
  logic [3:0] lizzieLet0_4QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet0_4QNone_Bool_2_argbuf_select_q <= (lizzieLet0_4QNone_Bool_2_argbuf_done ? 4'd0 :
                                                   lizzieLet0_4QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet0_4QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_4QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_4QNone_Bool_2_argbuf_emit_q <= (lizzieLet0_4QNone_Bool_2_argbuf_done ? 2'd0 :
                                                 lizzieLet0_4QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet0_4QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet0_4QNone_Bool_2_argbuf_emit_d = (lizzieLet0_4QNone_Bool_2_argbuf_emit_q | ({go_10_goMux_choice_d[0],
                                                                                              go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                                        go_10_goMux_data_r}));
  logic lizzieLet0_4QNone_Bool_2_argbuf_done;
  assign lizzieLet0_4QNone_Bool_2_argbuf_done = (& lizzieLet0_4QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet0_4QError_Bool_2_argbuf_r,
          lizzieLet0_4QVal_Bool_2_argbuf_r,
          lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r,
          lizzieLet0_4QNone_Bool_2_argbuf_r} = (lizzieLet0_4QNone_Bool_2_argbuf_done ? lizzieLet0_4QNone_Bool_2_argbuf_select_d :
                                                4'd0);
  assign go_10_goMux_data_d = ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet0_4QNone_Bool_2_argbuf_d :
                               ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d :
                                ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet0_4QVal_Bool_2_argbuf_d :
                                 ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet0_4QError_Bool_2_argbuf_d :
                                  1'd0))));
  assign go_10_goMux_choice_d = ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet0_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet0_4QNone_Bool_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet0_4QVal_Bool,Go) > [(lizzieLet0_4QVal_Bool_1,Go),
                                             (lizzieLet0_4QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet0_4QVal_Bool_emitted;
  logic [1:0] lizzieLet0_4QVal_Bool_done;
  assign lizzieLet0_4QVal_Bool_1_d = (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[0]));
  assign lizzieLet0_4QVal_Bool_2_d = (lizzieLet0_4QVal_Bool_d[0] && (! lizzieLet0_4QVal_Bool_emitted[1]));
  assign lizzieLet0_4QVal_Bool_done = (lizzieLet0_4QVal_Bool_emitted | ({lizzieLet0_4QVal_Bool_2_d[0],
                                                                         lizzieLet0_4QVal_Bool_1_d[0]} & {lizzieLet0_4QVal_Bool_2_r,
                                                                                                          lizzieLet0_4QVal_Bool_1_r}));
  assign lizzieLet0_4QVal_Bool_r = (& lizzieLet0_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet0_4QVal_Bool_emitted <= (lizzieLet0_4QVal_Bool_r ? 2'd0 :
                                        lizzieLet0_4QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_1,Go) > (lizzieLet0_4QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_1_bufchan_d;
  logic lizzieLet0_4QVal_Bool_1_bufchan_r;
  assign lizzieLet0_4QVal_Bool_1_r = ((! lizzieLet0_4QVal_Bool_1_bufchan_d[0]) || lizzieLet0_4QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_1_r)
        lizzieLet0_4QVal_Bool_1_bufchan_d <= lizzieLet0_4QVal_Bool_1_d;
  Go_t lizzieLet0_4QVal_Bool_1_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_1_bufchan_r = (! lizzieLet0_4QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_1_argbuf_d = (lizzieLet0_4QVal_Bool_1_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_1_bufchan_buf :
                                             lizzieLet0_4QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_1_argbuf_r && lizzieLet0_4QVal_Bool_1_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_1_argbuf_r) && (! lizzieLet0_4QVal_Bool_1_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_1_bufchan_buf <= lizzieLet0_4QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) : [(lizzieLet0_4QVal_Bool_1_argbuf,Go),
                                                                                        (lizzieLet0_5QVal_Bool_1_argbuf,MyDTBool_Bool),
                                                                                        (lizzieLet0_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool),
                                                                                        (vacN_1_argbuf,MyBool),
                                                                                        (lizzieLet0_6QVal_Bool_1_argbuf,Pointer_QTree_Bool)] > (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) */
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d  = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_dc((& {lizzieLet0_4QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet0_5QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet0_3QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    vacN_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet0_6QVal_Bool_1_argbuf_d[0]}), lizzieLet0_4QVal_Bool_1_argbuf_d, lizzieLet0_5QVal_Bool_1_argbuf_d, lizzieLet0_3QVal_Bool_1_argbuf_d, vacN_1_argbuf_d, lizzieLet0_6QVal_Bool_1_argbuf_d);
  assign {lizzieLet0_4QVal_Bool_1_argbuf_r,
          lizzieLet0_5QVal_Bool_1_argbuf_r,
          lizzieLet0_3QVal_Bool_1_argbuf_r,
          vacN_1_argbuf_r,
          lizzieLet0_6QVal_Bool_1_argbuf_r} = {5 {(\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet0_4QVal_Bool_2,Go) > (lizzieLet0_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet0_4QVal_Bool_2_bufchan_d;
  logic lizzieLet0_4QVal_Bool_2_bufchan_r;
  assign lizzieLet0_4QVal_Bool_2_r = ((! lizzieLet0_4QVal_Bool_2_bufchan_d[0]) || lizzieLet0_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_4QVal_Bool_2_r)
        lizzieLet0_4QVal_Bool_2_bufchan_d <= lizzieLet0_4QVal_Bool_2_d;
  Go_t lizzieLet0_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet0_4QVal_Bool_2_bufchan_r = (! lizzieLet0_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_4QVal_Bool_2_argbuf_d = (lizzieLet0_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet0_4QVal_Bool_2_bufchan_buf :
                                             lizzieLet0_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_4QVal_Bool_2_argbuf_r && lizzieLet0_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet0_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_4QVal_Bool_2_argbuf_r) && (! lizzieLet0_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet0_4QVal_Bool_2_bufchan_buf <= lizzieLet0_4QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool) : (lizzieLet0_5,QTree_Bool) (isZacJ_goMux_mux,MyDTBool_Bool) > [(_38,MyDTBool_Bool),
                                                                                         (lizzieLet0_5QVal_Bool,MyDTBool_Bool),
                                                                                         (lizzieLet0_5QNode_Bool,MyDTBool_Bool),
                                                                                         (_37,MyDTBool_Bool)] */
  logic [3:0] isZacJ_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_5_d[0] && isZacJ_goMux_mux_d[0]))
      unique case (lizzieLet0_5_d[2:1])
        2'd0: isZacJ_goMux_mux_onehotd = 4'd1;
        2'd1: isZacJ_goMux_mux_onehotd = 4'd2;
        2'd2: isZacJ_goMux_mux_onehotd = 4'd4;
        2'd3: isZacJ_goMux_mux_onehotd = 4'd8;
        default: isZacJ_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacJ_goMux_mux_onehotd = 4'd0;
  assign _38_d = isZacJ_goMux_mux_onehotd[0];
  assign lizzieLet0_5QVal_Bool_d = isZacJ_goMux_mux_onehotd[1];
  assign lizzieLet0_5QNode_Bool_d = isZacJ_goMux_mux_onehotd[2];
  assign _37_d = isZacJ_goMux_mux_onehotd[3];
  assign isZacJ_goMux_mux_r = (| (isZacJ_goMux_mux_onehotd & {_37_r,
                                                              lizzieLet0_5QNode_Bool_r,
                                                              lizzieLet0_5QVal_Bool_r,
                                                              _38_r}));
  assign lizzieLet0_5_r = isZacJ_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool) : (lizzieLet0_5QNode_Bool,MyDTBool_Bool) > [(lizzieLet0_5QNode_Bool_1,MyDTBool_Bool),
                                                                    (lizzieLet0_5QNode_Bool_2,MyDTBool_Bool)] */
  logic [1:0] lizzieLet0_5QNode_Bool_emitted;
  logic [1:0] lizzieLet0_5QNode_Bool_done;
  assign lizzieLet0_5QNode_Bool_1_d = (lizzieLet0_5QNode_Bool_d[0] && (! lizzieLet0_5QNode_Bool_emitted[0]));
  assign lizzieLet0_5QNode_Bool_2_d = (lizzieLet0_5QNode_Bool_d[0] && (! lizzieLet0_5QNode_Bool_emitted[1]));
  assign lizzieLet0_5QNode_Bool_done = (lizzieLet0_5QNode_Bool_emitted | ({lizzieLet0_5QNode_Bool_2_d[0],
                                                                           lizzieLet0_5QNode_Bool_1_d[0]} & {lizzieLet0_5QNode_Bool_2_r,
                                                                                                             lizzieLet0_5QNode_Bool_1_r}));
  assign lizzieLet0_5QNode_Bool_r = (& lizzieLet0_5QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_5QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_5QNode_Bool_emitted <= (lizzieLet0_5QNode_Bool_r ? 2'd0 :
                                         lizzieLet0_5QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet0_5QNode_Bool_2,MyDTBool_Bool) > (lizzieLet0_5QNode_Bool_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_2_bufchan_d;
  logic lizzieLet0_5QNode_Bool_2_bufchan_r;
  assign lizzieLet0_5QNode_Bool_2_r = ((! lizzieLet0_5QNode_Bool_2_bufchan_d[0]) || lizzieLet0_5QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_5QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_5QNode_Bool_2_r)
        lizzieLet0_5QNode_Bool_2_bufchan_d <= lizzieLet0_5QNode_Bool_2_d;
  MyDTBool_Bool_t lizzieLet0_5QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_5QNode_Bool_2_bufchan_r = (! lizzieLet0_5QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_5QNode_Bool_2_argbuf_d = (lizzieLet0_5QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_5QNode_Bool_2_bufchan_buf :
                                              lizzieLet0_5QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_5QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_5QNode_Bool_2_argbuf_r && lizzieLet0_5QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_5QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_5QNode_Bool_2_argbuf_r) && (! lizzieLet0_5QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_5QNode_Bool_2_bufchan_buf <= lizzieLet0_5QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet0_5QVal_Bool,MyDTBool_Bool) > (lizzieLet0_5QVal_Bool_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet0_5QVal_Bool_bufchan_d;
  logic lizzieLet0_5QVal_Bool_bufchan_r;
  assign lizzieLet0_5QVal_Bool_r = ((! lizzieLet0_5QVal_Bool_bufchan_d[0]) || lizzieLet0_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_5QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet0_5QVal_Bool_r)
        lizzieLet0_5QVal_Bool_bufchan_d <= lizzieLet0_5QVal_Bool_d;
  MyDTBool_Bool_t lizzieLet0_5QVal_Bool_bufchan_buf;
  assign lizzieLet0_5QVal_Bool_bufchan_r = (! lizzieLet0_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_5QVal_Bool_1_argbuf_d = (lizzieLet0_5QVal_Bool_bufchan_buf[0] ? lizzieLet0_5QVal_Bool_bufchan_buf :
                                             lizzieLet0_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_5QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet0_5QVal_Bool_1_argbuf_r && lizzieLet0_5QVal_Bool_bufchan_buf[0]))
        lizzieLet0_5QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet0_5QVal_Bool_1_argbuf_r) && (! lizzieLet0_5QVal_Bool_bufchan_buf[0])))
        lizzieLet0_5QVal_Bool_bufchan_buf <= lizzieLet0_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet0_6,QTree_Bool) (m2acM_goMux_mux,Pointer_QTree_Bool) > [(_36,Pointer_QTree_Bool),
                                                                                                  (lizzieLet0_6QVal_Bool,Pointer_QTree_Bool),
                                                                                                  (lizzieLet0_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                  (_35,Pointer_QTree_Bool)] */
  logic [3:0] m2acM_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_6_d[0] && m2acM_goMux_mux_d[0]))
      unique case (lizzieLet0_6_d[2:1])
        2'd0: m2acM_goMux_mux_onehotd = 4'd1;
        2'd1: m2acM_goMux_mux_onehotd = 4'd2;
        2'd2: m2acM_goMux_mux_onehotd = 4'd4;
        2'd3: m2acM_goMux_mux_onehotd = 4'd8;
        default: m2acM_goMux_mux_onehotd = 4'd0;
      endcase
    else m2acM_goMux_mux_onehotd = 4'd0;
  assign _36_d = {m2acM_goMux_mux_d[16:1],
                  m2acM_goMux_mux_onehotd[0]};
  assign lizzieLet0_6QVal_Bool_d = {m2acM_goMux_mux_d[16:1],
                                    m2acM_goMux_mux_onehotd[1]};
  assign lizzieLet0_6QNode_Bool_d = {m2acM_goMux_mux_d[16:1],
                                     m2acM_goMux_mux_onehotd[2]};
  assign _35_d = {m2acM_goMux_mux_d[16:1],
                  m2acM_goMux_mux_onehotd[3]};
  assign m2acM_goMux_mux_r = (| (m2acM_goMux_mux_onehotd & {_35_r,
                                                            lizzieLet0_6QNode_Bool_r,
                                                            lizzieLet0_6QVal_Bool_r,
                                                            _36_r}));
  assign lizzieLet0_6_r = m2acM_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet0_6QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet0_6QNode_Bool_1,Pointer_QTree_Bool),
                                                                              (lizzieLet0_6QNode_Bool_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet0_6QNode_Bool_emitted;
  logic [1:0] lizzieLet0_6QNode_Bool_done;
  assign lizzieLet0_6QNode_Bool_1_d = {lizzieLet0_6QNode_Bool_d[16:1],
                                       (lizzieLet0_6QNode_Bool_d[0] && (! lizzieLet0_6QNode_Bool_emitted[0]))};
  assign lizzieLet0_6QNode_Bool_2_d = {lizzieLet0_6QNode_Bool_d[16:1],
                                       (lizzieLet0_6QNode_Bool_d[0] && (! lizzieLet0_6QNode_Bool_emitted[1]))};
  assign lizzieLet0_6QNode_Bool_done = (lizzieLet0_6QNode_Bool_emitted | ({lizzieLet0_6QNode_Bool_2_d[0],
                                                                           lizzieLet0_6QNode_Bool_1_d[0]} & {lizzieLet0_6QNode_Bool_2_r,
                                                                                                             lizzieLet0_6QNode_Bool_1_r}));
  assign lizzieLet0_6QNode_Bool_r = (& lizzieLet0_6QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_6QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet0_6QNode_Bool_emitted <= (lizzieLet0_6QNode_Bool_r ? 2'd0 :
                                         lizzieLet0_6QNode_Bool_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_6QNode_Bool_2,Pointer_QTree_Bool) > (lizzieLet0_6QNode_Bool_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_2_bufchan_d;
  logic lizzieLet0_6QNode_Bool_2_bufchan_r;
  assign lizzieLet0_6QNode_Bool_2_r = ((! lizzieLet0_6QNode_Bool_2_bufchan_d[0]) || lizzieLet0_6QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_6QNode_Bool_2_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_6QNode_Bool_2_r)
        lizzieLet0_6QNode_Bool_2_bufchan_d <= lizzieLet0_6QNode_Bool_2_d;
  Pointer_QTree_Bool_t lizzieLet0_6QNode_Bool_2_bufchan_buf;
  assign lizzieLet0_6QNode_Bool_2_bufchan_r = (! lizzieLet0_6QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet0_6QNode_Bool_2_argbuf_d = (lizzieLet0_6QNode_Bool_2_bufchan_buf[0] ? lizzieLet0_6QNode_Bool_2_bufchan_buf :
                                              lizzieLet0_6QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_6QNode_Bool_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_6QNode_Bool_2_argbuf_r && lizzieLet0_6QNode_Bool_2_bufchan_buf[0]))
        lizzieLet0_6QNode_Bool_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_6QNode_Bool_2_argbuf_r) && (! lizzieLet0_6QNode_Bool_2_bufchan_buf[0])))
        lizzieLet0_6QNode_Bool_2_bufchan_buf <= lizzieLet0_6QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet0_6QVal_Bool,Pointer_QTree_Bool) > (lizzieLet0_6QVal_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet0_6QVal_Bool_bufchan_d;
  logic lizzieLet0_6QVal_Bool_bufchan_r;
  assign lizzieLet0_6QVal_Bool_r = ((! lizzieLet0_6QVal_Bool_bufchan_d[0]) || lizzieLet0_6QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_6QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_6QVal_Bool_r)
        lizzieLet0_6QVal_Bool_bufchan_d <= lizzieLet0_6QVal_Bool_d;
  Pointer_QTree_Bool_t lizzieLet0_6QVal_Bool_bufchan_buf;
  assign lizzieLet0_6QVal_Bool_bufchan_r = (! lizzieLet0_6QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_6QVal_Bool_1_argbuf_d = (lizzieLet0_6QVal_Bool_bufchan_buf[0] ? lizzieLet0_6QVal_Bool_bufchan_buf :
                                             lizzieLet0_6QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_6QVal_Bool_1_argbuf_r && lizzieLet0_6QVal_Bool_bufchan_buf[0]))
        lizzieLet0_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_6QVal_Bool_1_argbuf_r) && (! lizzieLet0_6QVal_Bool_bufchan_buf[0])))
        lizzieLet0_6QVal_Bool_bufchan_buf <= lizzieLet0_6QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet0_7,QTree_Bool) (sc_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) > [(lizzieLet0_7QNone_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet0_7QVal_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet0_7QNode_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet0_7QError_Bool,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet0_7_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet0_7_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet0_7QNone_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet0_7QVal_Bool_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet0_7QNode_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet0_7QError_Bool_d = {sc_0_goMux_mux_d[16:1],
                                      sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet0_7QError_Bool_r,
                                                          lizzieLet0_7QNode_Bool_r,
                                                          lizzieLet0_7QVal_Bool_r,
                                                          lizzieLet0_7QNone_Bool_r}));
  assign lizzieLet0_7_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet0_7QError_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet0_7QError_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QError_Bool_bufchan_d;
  logic lizzieLet0_7QError_Bool_bufchan_r;
  assign lizzieLet0_7QError_Bool_r = ((! lizzieLet0_7QError_Bool_bufchan_d[0]) || lizzieLet0_7QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_7QError_Bool_r)
        lizzieLet0_7QError_Bool_bufchan_d <= lizzieLet0_7QError_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QError_Bool_bufchan_buf;
  assign lizzieLet0_7QError_Bool_bufchan_r = (! lizzieLet0_7QError_Bool_bufchan_buf[0]);
  assign lizzieLet0_7QError_Bool_1_argbuf_d = (lizzieLet0_7QError_Bool_bufchan_buf[0] ? lizzieLet0_7QError_Bool_bufchan_buf :
                                               lizzieLet0_7QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_7QError_Bool_1_argbuf_r && lizzieLet0_7QError_Bool_bufchan_buf[0]))
        lizzieLet0_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_7QError_Bool_1_argbuf_r) && (! lizzieLet0_7QError_Bool_bufchan_buf[0])))
        lizzieLet0_7QError_Bool_bufchan_buf <= lizzieLet0_7QError_Bool_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool3) : [(lizzieLet0_7QNode_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (lizzieLet0_5QNode_Bool_1,MyDTBool_Bool),
                                               (lizzieLet0_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                               (q1acO_destruct,Pointer_QTree_Bool),
                                               (lizzieLet0_6QNode_Bool_1,Pointer_QTree_Bool),
                                               (q2acP_destruct,Pointer_QTree_Bool),
                                               (q3acQ_destruct,Pointer_QTree_Bool)] > (lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_d = Lcall_kron_kron_Bool_Bool_Bool3_dc((& {lizzieLet0_7QNode_Bool_d[0],
                                                                                                                                                                                                         lizzieLet0_5QNode_Bool_1_d[0],
                                                                                                                                                                                                         lizzieLet0_3QNode_Bool_1_d[0],
                                                                                                                                                                                                         q1acO_destruct_d[0],
                                                                                                                                                                                                         lizzieLet0_6QNode_Bool_1_d[0],
                                                                                                                                                                                                         q2acP_destruct_d[0],
                                                                                                                                                                                                         q3acQ_destruct_d[0]}), lizzieLet0_7QNode_Bool_d, lizzieLet0_5QNode_Bool_1_d, lizzieLet0_3QNode_Bool_1_d, q1acO_destruct_d, lizzieLet0_6QNode_Bool_1_d, q2acP_destruct_d, q3acQ_destruct_d);
  assign {lizzieLet0_7QNode_Bool_r,
          lizzieLet0_5QNode_Bool_1_r,
          lizzieLet0_3QNode_Bool_1_r,
          q1acO_destruct_r,
          lizzieLet0_6QNode_Bool_1_r,
          q2acP_destruct_r,
          q3acQ_destruct_r} = {7 {(lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_r && lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) > (lizzieLet2_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  logic lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r;
  assign lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_r = ((! lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d[0]) || lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= {83'd0,
                                                                                                                                                                         1'd0};
    else
      if (lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_r)
        lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf;
  assign lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r = (! lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0] ? lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf :
                                  lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= {83'd0,
                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]))
        lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= {83'd0,
                                                                                                                                                                             1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0])))
        lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= lizzieLet0_7QNode_Bool_1lizzieLet0_5QNode_Bool_1lizzieLet0_3QNode_Bool_1q1acO_1lizzieLet0_6QNode_Bool_1q2acP_1q3acQ_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet0_7QNone_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet0_7QNone_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNone_Bool_bufchan_d;
  logic lizzieLet0_7QNone_Bool_bufchan_r;
  assign lizzieLet0_7QNone_Bool_r = ((! lizzieLet0_7QNone_Bool_bufchan_d[0]) || lizzieLet0_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_7QNone_Bool_r)
        lizzieLet0_7QNone_Bool_bufchan_d <= lizzieLet0_7QNone_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QNone_Bool_bufchan_buf;
  assign lizzieLet0_7QNone_Bool_bufchan_r = (! lizzieLet0_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet0_7QNone_Bool_1_argbuf_d = (lizzieLet0_7QNone_Bool_bufchan_buf[0] ? lizzieLet0_7QNone_Bool_bufchan_buf :
                                              lizzieLet0_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_7QNone_Bool_1_argbuf_r && lizzieLet0_7QNone_Bool_bufchan_buf[0]))
        lizzieLet0_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_7QNone_Bool_1_argbuf_r) && (! lizzieLet0_7QNone_Bool_bufchan_buf[0])))
        lizzieLet0_7QNone_Bool_bufchan_buf <= lizzieLet0_7QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet0_7QVal_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet0_7QVal_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QVal_Bool_bufchan_d;
  logic lizzieLet0_7QVal_Bool_bufchan_r;
  assign lizzieLet0_7QVal_Bool_r = ((! lizzieLet0_7QVal_Bool_bufchan_d[0]) || lizzieLet0_7QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet0_7QVal_Bool_r)
        lizzieLet0_7QVal_Bool_bufchan_d <= lizzieLet0_7QVal_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet0_7QVal_Bool_bufchan_buf;
  assign lizzieLet0_7QVal_Bool_bufchan_r = (! lizzieLet0_7QVal_Bool_bufchan_buf[0]);
  assign lizzieLet0_7QVal_Bool_1_argbuf_d = (lizzieLet0_7QVal_Bool_bufchan_buf[0] ? lizzieLet0_7QVal_Bool_bufchan_buf :
                                             lizzieLet0_7QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_7QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_7QVal_Bool_1_argbuf_r && lizzieLet0_7QVal_Bool_bufchan_buf[0]))
        lizzieLet0_7QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_7QVal_Bool_1_argbuf_r) && (! lizzieLet0_7QVal_Bool_bufchan_buf[0])))
        lizzieLet0_7QVal_Bool_bufchan_buf <= lizzieLet0_7QVal_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet11_1_1QNode_Bool,QTree_Bool) > [(q1acF_destruct,Pointer_QTree_Bool),
                                                                       (q2acG_destruct,Pointer_QTree_Bool),
                                                                       (q3acH_destruct,Pointer_QTree_Bool),
                                                                       (q4acI_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet11_1_1QNode_Bool_emitted;
  logic [3:0] lizzieLet11_1_1QNode_Bool_done;
  assign q1acF_destruct_d = {lizzieLet11_1_1QNode_Bool_d[18:3],
                             (lizzieLet11_1_1QNode_Bool_d[0] && (! lizzieLet11_1_1QNode_Bool_emitted[0]))};
  assign q2acG_destruct_d = {lizzieLet11_1_1QNode_Bool_d[34:19],
                             (lizzieLet11_1_1QNode_Bool_d[0] && (! lizzieLet11_1_1QNode_Bool_emitted[1]))};
  assign q3acH_destruct_d = {lizzieLet11_1_1QNode_Bool_d[50:35],
                             (lizzieLet11_1_1QNode_Bool_d[0] && (! lizzieLet11_1_1QNode_Bool_emitted[2]))};
  assign q4acI_destruct_d = {lizzieLet11_1_1QNode_Bool_d[66:51],
                             (lizzieLet11_1_1QNode_Bool_d[0] && (! lizzieLet11_1_1QNode_Bool_emitted[3]))};
  assign lizzieLet11_1_1QNode_Bool_done = (lizzieLet11_1_1QNode_Bool_emitted | ({q4acI_destruct_d[0],
                                                                                 q3acH_destruct_d[0],
                                                                                 q2acG_destruct_d[0],
                                                                                 q1acF_destruct_d[0]} & {q4acI_destruct_r,
                                                                                                         q3acH_destruct_r,
                                                                                                         q2acG_destruct_r,
                                                                                                         q1acF_destruct_r}));
  assign lizzieLet11_1_1QNode_Bool_r = (& lizzieLet11_1_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet11_1_1QNode_Bool_emitted <= (lizzieLet11_1_1QNode_Bool_r ? 4'd0 :
                                            lizzieLet11_1_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet11_1_1QVal_Bool,QTree_Bool) > [(vacE_destruct,MyBool)] */
  assign vacE_destruct_d = {lizzieLet11_1_1QVal_Bool_d[3:3],
                            lizzieLet11_1_1QVal_Bool_d[0]};
  assign lizzieLet11_1_1QVal_Bool_r = vacE_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet11_1_2,QTree_Bool) (lizzieLet11_1_1,QTree_Bool) > [(_34,QTree_Bool),
                                                                                     (lizzieLet11_1_1QVal_Bool,QTree_Bool),
                                                                                     (lizzieLet11_1_1QNode_Bool,QTree_Bool),
                                                                                     (_33,QTree_Bool)] */
  logic [3:0] lizzieLet11_1_1_onehotd;
  always_comb
    if ((lizzieLet11_1_2_d[0] && lizzieLet11_1_1_d[0]))
      unique case (lizzieLet11_1_2_d[2:1])
        2'd0: lizzieLet11_1_1_onehotd = 4'd1;
        2'd1: lizzieLet11_1_1_onehotd = 4'd2;
        2'd2: lizzieLet11_1_1_onehotd = 4'd4;
        2'd3: lizzieLet11_1_1_onehotd = 4'd8;
        default: lizzieLet11_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet11_1_1_onehotd = 4'd0;
  assign _34_d = {lizzieLet11_1_1_d[66:1],
                  lizzieLet11_1_1_onehotd[0]};
  assign lizzieLet11_1_1QVal_Bool_d = {lizzieLet11_1_1_d[66:1],
                                       lizzieLet11_1_1_onehotd[1]};
  assign lizzieLet11_1_1QNode_Bool_d = {lizzieLet11_1_1_d[66:1],
                                        lizzieLet11_1_1_onehotd[2]};
  assign _33_d = {lizzieLet11_1_1_d[66:1],
                  lizzieLet11_1_1_onehotd[3]};
  assign lizzieLet11_1_1_r = (| (lizzieLet11_1_1_onehotd & {_33_r,
                                                            lizzieLet11_1_1QNode_Bool_r,
                                                            lizzieLet11_1_1QVal_Bool_r,
                                                            _34_r}));
  assign lizzieLet11_1_2_r = lizzieLet11_1_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet11_1_3,QTree_Bool) (gacB_goMux_mux,MyDTBool_Bool_Bool) > [(_32,MyDTBool_Bool_Bool),
                                                                                                    (lizzieLet11_1_3QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                    (lizzieLet11_1_3QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                    (_31,MyDTBool_Bool_Bool)] */
  logic [3:0] gacB_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet11_1_3_d[0] && gacB_goMux_mux_d[0]))
      unique case (lizzieLet11_1_3_d[2:1])
        2'd0: gacB_goMux_mux_onehotd = 4'd1;
        2'd1: gacB_goMux_mux_onehotd = 4'd2;
        2'd2: gacB_goMux_mux_onehotd = 4'd4;
        2'd3: gacB_goMux_mux_onehotd = 4'd8;
        default: gacB_goMux_mux_onehotd = 4'd0;
      endcase
    else gacB_goMux_mux_onehotd = 4'd0;
  assign _32_d = gacB_goMux_mux_onehotd[0];
  assign lizzieLet11_1_3QVal_Bool_d = gacB_goMux_mux_onehotd[1];
  assign lizzieLet11_1_3QNode_Bool_d = gacB_goMux_mux_onehotd[2];
  assign _31_d = gacB_goMux_mux_onehotd[3];
  assign gacB_goMux_mux_r = (| (gacB_goMux_mux_onehotd & {_31_r,
                                                          lizzieLet11_1_3QNode_Bool_r,
                                                          lizzieLet11_1_3QVal_Bool_r,
                                                          _32_r}));
  assign lizzieLet11_1_3_r = gacB_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (lizzieLet11_1_3QNode_Bool,MyDTBool_Bool_Bool) > [(lizzieLet11_1_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                                                 (lizzieLet11_1_3QNode_Bool_2,MyDTBool_Bool_Bool)] */
  logic [1:0] lizzieLet11_1_3QNode_Bool_emitted;
  logic [1:0] lizzieLet11_1_3QNode_Bool_done;
  assign lizzieLet11_1_3QNode_Bool_1_d = (lizzieLet11_1_3QNode_Bool_d[0] && (! lizzieLet11_1_3QNode_Bool_emitted[0]));
  assign lizzieLet11_1_3QNode_Bool_2_d = (lizzieLet11_1_3QNode_Bool_d[0] && (! lizzieLet11_1_3QNode_Bool_emitted[1]));
  assign lizzieLet11_1_3QNode_Bool_done = (lizzieLet11_1_3QNode_Bool_emitted | ({lizzieLet11_1_3QNode_Bool_2_d[0],
                                                                                 lizzieLet11_1_3QNode_Bool_1_d[0]} & {lizzieLet11_1_3QNode_Bool_2_r,
                                                                                                                      lizzieLet11_1_3QNode_Bool_1_r}));
  assign lizzieLet11_1_3QNode_Bool_r = (& lizzieLet11_1_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_3QNode_Bool_emitted <= (lizzieLet11_1_3QNode_Bool_r ? 2'd0 :
                                            lizzieLet11_1_3QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet11_1_3QNode_Bool_2,MyDTBool_Bool_Bool) > (lizzieLet11_1_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_2_bufchan_d;
  logic lizzieLet11_1_3QNode_Bool_2_bufchan_r;
  assign lizzieLet11_1_3QNode_Bool_2_r = ((! lizzieLet11_1_3QNode_Bool_2_bufchan_d[0]) || lizzieLet11_1_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_3QNode_Bool_2_r)
        lizzieLet11_1_3QNode_Bool_2_bufchan_d <= lizzieLet11_1_3QNode_Bool_2_d;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet11_1_3QNode_Bool_2_bufchan_r = (! lizzieLet11_1_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_3QNode_Bool_2_argbuf_d = (lizzieLet11_1_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet11_1_3QNode_Bool_2_bufchan_buf :
                                                 lizzieLet11_1_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_3QNode_Bool_2_argbuf_r && lizzieLet11_1_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_3QNode_Bool_2_argbuf_r) && (! lizzieLet11_1_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_3QNode_Bool_2_bufchan_buf <= lizzieLet11_1_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet11_1_3QVal_Bool,MyDTBool_Bool_Bool) > (lizzieLet11_1_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QVal_Bool_bufchan_d;
  logic lizzieLet11_1_3QVal_Bool_bufchan_r;
  assign lizzieLet11_1_3QVal_Bool_r = ((! lizzieLet11_1_3QVal_Bool_bufchan_d[0]) || lizzieLet11_1_3QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_3QVal_Bool_r)
        lizzieLet11_1_3QVal_Bool_bufchan_d <= lizzieLet11_1_3QVal_Bool_d;
  MyDTBool_Bool_Bool_t lizzieLet11_1_3QVal_Bool_bufchan_buf;
  assign lizzieLet11_1_3QVal_Bool_bufchan_r = (! lizzieLet11_1_3QVal_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_3QVal_Bool_1_argbuf_d = (lizzieLet11_1_3QVal_Bool_bufchan_buf[0] ? lizzieLet11_1_3QVal_Bool_bufchan_buf :
                                                lizzieLet11_1_3QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_3QVal_Bool_1_argbuf_r && lizzieLet11_1_3QVal_Bool_bufchan_buf[0]))
        lizzieLet11_1_3QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_3QVal_Bool_1_argbuf_r) && (! lizzieLet11_1_3QVal_Bool_bufchan_buf[0])))
        lizzieLet11_1_3QVal_Bool_bufchan_buf <= lizzieLet11_1_3QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet11_1_4,QTree_Bool) (go_6_goMux_data,Go) > [(lizzieLet11_1_4QNone_Bool,Go),
                                                                     (lizzieLet11_1_4QVal_Bool,Go),
                                                                     (lizzieLet11_1_4QNode_Bool,Go),
                                                                     (lizzieLet11_1_4QError_Bool,Go)] */
  logic [3:0] go_6_goMux_data_onehotd;
  always_comb
    if ((lizzieLet11_1_4_d[0] && go_6_goMux_data_d[0]))
      unique case (lizzieLet11_1_4_d[2:1])
        2'd0: go_6_goMux_data_onehotd = 4'd1;
        2'd1: go_6_goMux_data_onehotd = 4'd2;
        2'd2: go_6_goMux_data_onehotd = 4'd4;
        2'd3: go_6_goMux_data_onehotd = 4'd8;
        default: go_6_goMux_data_onehotd = 4'd0;
      endcase
    else go_6_goMux_data_onehotd = 4'd0;
  assign lizzieLet11_1_4QNone_Bool_d = go_6_goMux_data_onehotd[0];
  assign lizzieLet11_1_4QVal_Bool_d = go_6_goMux_data_onehotd[1];
  assign lizzieLet11_1_4QNode_Bool_d = go_6_goMux_data_onehotd[2];
  assign lizzieLet11_1_4QError_Bool_d = go_6_goMux_data_onehotd[3];
  assign go_6_goMux_data_r = (| (go_6_goMux_data_onehotd & {lizzieLet11_1_4QError_Bool_r,
                                                            lizzieLet11_1_4QNode_Bool_r,
                                                            lizzieLet11_1_4QVal_Bool_r,
                                                            lizzieLet11_1_4QNone_Bool_r}));
  assign lizzieLet11_1_4_r = go_6_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet11_1_4QError_Bool,Go) > [(lizzieLet11_1_4QError_Bool_1,Go),
                                                  (lizzieLet11_1_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet11_1_4QError_Bool_emitted;
  logic [1:0] lizzieLet11_1_4QError_Bool_done;
  assign lizzieLet11_1_4QError_Bool_1_d = (lizzieLet11_1_4QError_Bool_d[0] && (! lizzieLet11_1_4QError_Bool_emitted[0]));
  assign lizzieLet11_1_4QError_Bool_2_d = (lizzieLet11_1_4QError_Bool_d[0] && (! lizzieLet11_1_4QError_Bool_emitted[1]));
  assign lizzieLet11_1_4QError_Bool_done = (lizzieLet11_1_4QError_Bool_emitted | ({lizzieLet11_1_4QError_Bool_2_d[0],
                                                                                   lizzieLet11_1_4QError_Bool_1_d[0]} & {lizzieLet11_1_4QError_Bool_2_r,
                                                                                                                         lizzieLet11_1_4QError_Bool_1_r}));
  assign lizzieLet11_1_4QError_Bool_r = (& lizzieLet11_1_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_4QError_Bool_emitted <= (lizzieLet11_1_4QError_Bool_r ? 2'd0 :
                                             lizzieLet11_1_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet11_1_4QError_Bool_1,Go)] > (lizzieLet11_1_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet11_1_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet11_1_4QError_Bool_1_d[0]}), lizzieLet11_1_4QError_Bool_1_d);
  assign {lizzieLet11_1_4QError_Bool_1_r} = {1 {(lizzieLet11_1_4QError_Bool_1QError_Bool_r && lizzieLet11_1_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet16_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet11_1_4QError_Bool_1QError_Bool_r = ((! lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet11_1_4QError_Bool_1QError_Bool_r)
        lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet11_1_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                              1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet11_1_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4QError_Bool_2,Go) > (lizzieLet11_1_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4QError_Bool_2_bufchan_d;
  logic lizzieLet11_1_4QError_Bool_2_bufchan_r;
  assign lizzieLet11_1_4QError_Bool_2_r = ((! lizzieLet11_1_4QError_Bool_2_bufchan_d[0]) || lizzieLet11_1_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4QError_Bool_2_r)
        lizzieLet11_1_4QError_Bool_2_bufchan_d <= lizzieLet11_1_4QError_Bool_2_d;
  Go_t lizzieLet11_1_4QError_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4QError_Bool_2_bufchan_r = (! lizzieLet11_1_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4QError_Bool_2_argbuf_d = (lizzieLet11_1_4QError_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4QError_Bool_2_bufchan_buf :
                                                  lizzieLet11_1_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4QError_Bool_2_argbuf_r && lizzieLet11_1_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4QError_Bool_2_argbuf_r) && (! lizzieLet11_1_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4QError_Bool_2_bufchan_buf <= lizzieLet11_1_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4QNode_Bool,Go) > (lizzieLet11_1_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet11_1_4QNode_Bool_bufchan_d;
  logic lizzieLet11_1_4QNode_Bool_bufchan_r;
  assign lizzieLet11_1_4QNode_Bool_r = ((! lizzieLet11_1_4QNode_Bool_bufchan_d[0]) || lizzieLet11_1_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4QNode_Bool_r)
        lizzieLet11_1_4QNode_Bool_bufchan_d <= lizzieLet11_1_4QNode_Bool_d;
  Go_t lizzieLet11_1_4QNode_Bool_bufchan_buf;
  assign lizzieLet11_1_4QNode_Bool_bufchan_r = (! lizzieLet11_1_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4QNode_Bool_1_argbuf_d = (lizzieLet11_1_4QNode_Bool_bufchan_buf[0] ? lizzieLet11_1_4QNode_Bool_bufchan_buf :
                                                 lizzieLet11_1_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4QNode_Bool_1_argbuf_r && lizzieLet11_1_4QNode_Bool_bufchan_buf[0]))
        lizzieLet11_1_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4QNode_Bool_1_argbuf_r) && (! lizzieLet11_1_4QNode_Bool_bufchan_buf[0])))
        lizzieLet11_1_4QNode_Bool_bufchan_buf <= lizzieLet11_1_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet11_1_4QNone_Bool,Go) > [(lizzieLet11_1_4QNone_Bool_1,Go),
                                                 (lizzieLet11_1_4QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet11_1_4QNone_Bool_emitted;
  logic [1:0] lizzieLet11_1_4QNone_Bool_done;
  assign lizzieLet11_1_4QNone_Bool_1_d = (lizzieLet11_1_4QNone_Bool_d[0] && (! lizzieLet11_1_4QNone_Bool_emitted[0]));
  assign lizzieLet11_1_4QNone_Bool_2_d = (lizzieLet11_1_4QNone_Bool_d[0] && (! lizzieLet11_1_4QNone_Bool_emitted[1]));
  assign lizzieLet11_1_4QNone_Bool_done = (lizzieLet11_1_4QNone_Bool_emitted | ({lizzieLet11_1_4QNone_Bool_2_d[0],
                                                                                 lizzieLet11_1_4QNone_Bool_1_d[0]} & {lizzieLet11_1_4QNone_Bool_2_r,
                                                                                                                      lizzieLet11_1_4QNone_Bool_1_r}));
  assign lizzieLet11_1_4QNone_Bool_r = (& lizzieLet11_1_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_4QNone_Bool_emitted <= (lizzieLet11_1_4QNone_Bool_r ? 2'd0 :
                                            lizzieLet11_1_4QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet11_1_4QNone_Bool_1,Go)] > (lizzieLet11_1_4QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet11_1_4QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet11_1_4QNone_Bool_1_d[0]}), lizzieLet11_1_4QNone_Bool_1_d);
  assign {lizzieLet11_1_4QNone_Bool_1_r} = {1 {(lizzieLet11_1_4QNone_Bool_1QNone_Bool_r && lizzieLet11_1_4QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_4QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet12_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet11_1_4QNone_Bool_1QNone_Bool_r = ((! lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet11_1_4QNone_Bool_1QNone_Bool_r)
        lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet11_1_4QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf :
                                     lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet11_1_4QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4QNone_Bool_2,Go) > (lizzieLet11_1_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4QNone_Bool_2_bufchan_d;
  logic lizzieLet11_1_4QNone_Bool_2_bufchan_r;
  assign lizzieLet11_1_4QNone_Bool_2_r = ((! lizzieLet11_1_4QNone_Bool_2_bufchan_d[0]) || lizzieLet11_1_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4QNone_Bool_2_r)
        lizzieLet11_1_4QNone_Bool_2_bufchan_d <= lizzieLet11_1_4QNone_Bool_2_d;
  Go_t lizzieLet11_1_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4QNone_Bool_2_bufchan_r = (! lizzieLet11_1_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4QNone_Bool_2_argbuf_d = (lizzieLet11_1_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4QNone_Bool_2_bufchan_buf :
                                                 lizzieLet11_1_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4QNone_Bool_2_argbuf_r && lizzieLet11_1_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4QNone_Bool_2_argbuf_r) && (! lizzieLet11_1_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4QNone_Bool_2_bufchan_buf <= lizzieLet11_1_4QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet11_1_4QNone_Bool_2_argbuf,Go),
                           (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf,Go),
                           (es_0_1_1MyFalse_1_argbuf,Go),
                           (es_0_1_1MyTrue_2_argbuf,Go),
                           (lizzieLet11_1_4QError_Bool_2_argbuf,Go)] > (go_12_goMux_choice,C5) (go_12_goMux_data,Go) */
  logic [4:0] lizzieLet11_1_4QNone_Bool_2_argbuf_select_d;
  assign lizzieLet11_1_4QNone_Bool_2_argbuf_select_d = ((| lizzieLet11_1_4QNone_Bool_2_argbuf_select_q) ? lizzieLet11_1_4QNone_Bool_2_argbuf_select_q :
                                                        (lizzieLet11_1_4QNone_Bool_2_argbuf_d[0] ? 5'd1 :
                                                         (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d [0] ? 5'd2 :
                                                          (es_0_1_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                           (es_0_1_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                            (lizzieLet11_1_4QError_Bool_2_argbuf_d[0] ? 5'd16 :
                                                             5'd0))))));
  logic [4:0] lizzieLet11_1_4QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QNone_Bool_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet11_1_4QNone_Bool_2_argbuf_select_q <= (lizzieLet11_1_4QNone_Bool_2_argbuf_done ? 5'd0 :
                                                      lizzieLet11_1_4QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q <= (lizzieLet11_1_4QNone_Bool_2_argbuf_done ? 2'd0 :
                                                    lizzieLet11_1_4QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_4QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet11_1_4QNone_Bool_2_argbuf_emit_d = (lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q | ({go_12_goMux_choice_d[0],
                                                                                                    go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                                                              go_12_goMux_data_r}));
  logic lizzieLet11_1_4QNone_Bool_2_argbuf_done;
  assign lizzieLet11_1_4QNone_Bool_2_argbuf_done = (& lizzieLet11_1_4QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet11_1_4QError_Bool_2_argbuf_r,
          es_0_1_1MyTrue_2_argbuf_r,
          es_0_1_1MyFalse_1_argbuf_r,
          \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ,
          lizzieLet11_1_4QNone_Bool_2_argbuf_r} = (lizzieLet11_1_4QNone_Bool_2_argbuf_done ? lizzieLet11_1_4QNone_Bool_2_argbuf_select_d :
                                                   5'd0);
  assign go_12_goMux_data_d = ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet11_1_4QNone_Bool_2_argbuf_d :
                               ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[0])) ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d  :
                                ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_1_1MyFalse_1_argbuf_d :
                                 ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_1_1MyTrue_2_argbuf_d :
                                  ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet11_1_4QError_Bool_2_argbuf_d :
                                   1'd0)))));
  assign go_12_goMux_choice_d = ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet11_1_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet11_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet11_1_4QVal_Bool,Go) > [(lizzieLet11_1_4QVal_Bool_1,Go),
                                                (lizzieLet11_1_4QVal_Bool_2,Go),
                                                (lizzieLet11_1_4QVal_Bool_3,Go)] */
  logic [2:0] lizzieLet11_1_4QVal_Bool_emitted;
  logic [2:0] lizzieLet11_1_4QVal_Bool_done;
  assign lizzieLet11_1_4QVal_Bool_1_d = (lizzieLet11_1_4QVal_Bool_d[0] && (! lizzieLet11_1_4QVal_Bool_emitted[0]));
  assign lizzieLet11_1_4QVal_Bool_2_d = (lizzieLet11_1_4QVal_Bool_d[0] && (! lizzieLet11_1_4QVal_Bool_emitted[1]));
  assign lizzieLet11_1_4QVal_Bool_3_d = (lizzieLet11_1_4QVal_Bool_d[0] && (! lizzieLet11_1_4QVal_Bool_emitted[2]));
  assign lizzieLet11_1_4QVal_Bool_done = (lizzieLet11_1_4QVal_Bool_emitted | ({lizzieLet11_1_4QVal_Bool_3_d[0],
                                                                               lizzieLet11_1_4QVal_Bool_2_d[0],
                                                                               lizzieLet11_1_4QVal_Bool_1_d[0]} & {lizzieLet11_1_4QVal_Bool_3_r,
                                                                                                                   lizzieLet11_1_4QVal_Bool_2_r,
                                                                                                                   lizzieLet11_1_4QVal_Bool_1_r}));
  assign lizzieLet11_1_4QVal_Bool_r = (& lizzieLet11_1_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet11_1_4QVal_Bool_emitted <= (lizzieLet11_1_4QVal_Bool_r ? 3'd0 :
                                           lizzieLet11_1_4QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet11_1_4QVal_Bool_1,Go) > (lizzieLet11_1_4QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet11_1_4QVal_Bool_1_bufchan_d;
  logic lizzieLet11_1_4QVal_Bool_1_bufchan_r;
  assign lizzieLet11_1_4QVal_Bool_1_r = ((! lizzieLet11_1_4QVal_Bool_1_bufchan_d[0]) || lizzieLet11_1_4QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4QVal_Bool_1_r)
        lizzieLet11_1_4QVal_Bool_1_bufchan_d <= lizzieLet11_1_4QVal_Bool_1_d;
  Go_t lizzieLet11_1_4QVal_Bool_1_bufchan_buf;
  assign lizzieLet11_1_4QVal_Bool_1_bufchan_r = (! lizzieLet11_1_4QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet11_1_4QVal_Bool_1_argbuf_d = (lizzieLet11_1_4QVal_Bool_1_bufchan_buf[0] ? lizzieLet11_1_4QVal_Bool_1_bufchan_buf :
                                                lizzieLet11_1_4QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4QVal_Bool_1_argbuf_r && lizzieLet11_1_4QVal_Bool_1_bufchan_buf[0]))
        lizzieLet11_1_4QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4QVal_Bool_1_argbuf_r) && (! lizzieLet11_1_4QVal_Bool_1_bufchan_buf[0])))
        lizzieLet11_1_4QVal_Bool_1_bufchan_buf <= lizzieLet11_1_4QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
      Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : [(lizzieLet11_1_4QVal_Bool_1_argbuf,Go),
                                                            (lizzieLet11_1_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool),
                                                            (lizzieLet11_1_7QVal_Bool_1_argbuf,MyBool),
                                                            (vacE_1_argbuf,MyBool)] > (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) */
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d = TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_dc((& {lizzieLet11_1_4QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet11_1_3QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet11_1_7QVal_Bool_1_argbuf_d[0],
                                                                                                                                       vacE_1_argbuf_d[0]}), lizzieLet11_1_4QVal_Bool_1_argbuf_d, lizzieLet11_1_3QVal_Bool_1_argbuf_d, lizzieLet11_1_7QVal_Bool_1_argbuf_d, vacE_1_argbuf_d);
  assign {lizzieLet11_1_4QVal_Bool_1_argbuf_r,
          lizzieLet11_1_3QVal_Bool_1_argbuf_r,
          lizzieLet11_1_7QVal_Bool_1_argbuf_r,
          vacE_1_argbuf_r} = {4 {(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet11_1_4QVal_Bool_2,Go) > (lizzieLet11_1_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4QVal_Bool_2_bufchan_d;
  logic lizzieLet11_1_4QVal_Bool_2_bufchan_r;
  assign lizzieLet11_1_4QVal_Bool_2_r = ((! lizzieLet11_1_4QVal_Bool_2_bufchan_d[0]) || lizzieLet11_1_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4QVal_Bool_2_r)
        lizzieLet11_1_4QVal_Bool_2_bufchan_d <= lizzieLet11_1_4QVal_Bool_2_d;
  Go_t lizzieLet11_1_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4QVal_Bool_2_bufchan_r = (! lizzieLet11_1_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4QVal_Bool_2_argbuf_d = (lizzieLet11_1_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4QVal_Bool_2_bufchan_buf :
                                                lizzieLet11_1_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4QVal_Bool_2_argbuf_r && lizzieLet11_1_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4QVal_Bool_2_argbuf_r) && (! lizzieLet11_1_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4QVal_Bool_2_bufchan_buf <= lizzieLet11_1_4QVal_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyBool,
      Dcon TupGo___MyDTBool_Bool___MyBool) : [(lizzieLet11_1_4QVal_Bool_2_argbuf,Go),
                                              (lizzieLet11_1_5QVal_Bool_1_argbuf,MyDTBool_Bool),
                                              (xabY_1_argbuf,MyBool)] > (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) */
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d = TupGo___MyDTBool_Bool___MyBool_dc((& {lizzieLet11_1_4QVal_Bool_2_argbuf_d[0],
                                                                                                      lizzieLet11_1_5QVal_Bool_1_argbuf_d[0],
                                                                                                      xabY_1_argbuf_d[0]}), lizzieLet11_1_4QVal_Bool_2_argbuf_d, lizzieLet11_1_5QVal_Bool_1_argbuf_d, xabY_1_argbuf_d);
  assign {lizzieLet11_1_4QVal_Bool_2_argbuf_r,
          lizzieLet11_1_5QVal_Bool_1_argbuf_r,
          xabY_1_argbuf_r} = {3 {(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0])}};
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool) : (lizzieLet11_1_5,QTree_Bool) (isZacA_goMux_mux,MyDTBool_Bool) > [(_30,MyDTBool_Bool),
                                                                                            (lizzieLet11_1_5QVal_Bool,MyDTBool_Bool),
                                                                                            (lizzieLet11_1_5QNode_Bool,MyDTBool_Bool),
                                                                                            (_29,MyDTBool_Bool)] */
  logic [3:0] isZacA_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet11_1_5_d[0] && isZacA_goMux_mux_d[0]))
      unique case (lizzieLet11_1_5_d[2:1])
        2'd0: isZacA_goMux_mux_onehotd = 4'd1;
        2'd1: isZacA_goMux_mux_onehotd = 4'd2;
        2'd2: isZacA_goMux_mux_onehotd = 4'd4;
        2'd3: isZacA_goMux_mux_onehotd = 4'd8;
        default: isZacA_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacA_goMux_mux_onehotd = 4'd0;
  assign _30_d = isZacA_goMux_mux_onehotd[0];
  assign lizzieLet11_1_5QVal_Bool_d = isZacA_goMux_mux_onehotd[1];
  assign lizzieLet11_1_5QNode_Bool_d = isZacA_goMux_mux_onehotd[2];
  assign _29_d = isZacA_goMux_mux_onehotd[3];
  assign isZacA_goMux_mux_r = (| (isZacA_goMux_mux_onehotd & {_29_r,
                                                              lizzieLet11_1_5QNode_Bool_r,
                                                              lizzieLet11_1_5QVal_Bool_r,
                                                              _30_r}));
  assign lizzieLet11_1_5_r = isZacA_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool) : (lizzieLet11_1_5QNode_Bool,MyDTBool_Bool) > [(lizzieLet11_1_5QNode_Bool_1,MyDTBool_Bool),
                                                                       (lizzieLet11_1_5QNode_Bool_2,MyDTBool_Bool)] */
  logic [1:0] lizzieLet11_1_5QNode_Bool_emitted;
  logic [1:0] lizzieLet11_1_5QNode_Bool_done;
  assign lizzieLet11_1_5QNode_Bool_1_d = (lizzieLet11_1_5QNode_Bool_d[0] && (! lizzieLet11_1_5QNode_Bool_emitted[0]));
  assign lizzieLet11_1_5QNode_Bool_2_d = (lizzieLet11_1_5QNode_Bool_d[0] && (! lizzieLet11_1_5QNode_Bool_emitted[1]));
  assign lizzieLet11_1_5QNode_Bool_done = (lizzieLet11_1_5QNode_Bool_emitted | ({lizzieLet11_1_5QNode_Bool_2_d[0],
                                                                                 lizzieLet11_1_5QNode_Bool_1_d[0]} & {lizzieLet11_1_5QNode_Bool_2_r,
                                                                                                                      lizzieLet11_1_5QNode_Bool_1_r}));
  assign lizzieLet11_1_5QNode_Bool_r = (& lizzieLet11_1_5QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_5QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_5QNode_Bool_emitted <= (lizzieLet11_1_5QNode_Bool_r ? 2'd0 :
                                            lizzieLet11_1_5QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet11_1_5QNode_Bool_2,MyDTBool_Bool) > (lizzieLet11_1_5QNode_Bool_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_2_bufchan_d;
  logic lizzieLet11_1_5QNode_Bool_2_bufchan_r;
  assign lizzieLet11_1_5QNode_Bool_2_r = ((! lizzieLet11_1_5QNode_Bool_2_bufchan_d[0]) || lizzieLet11_1_5QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_5QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_5QNode_Bool_2_r)
        lizzieLet11_1_5QNode_Bool_2_bufchan_d <= lizzieLet11_1_5QNode_Bool_2_d;
  MyDTBool_Bool_t lizzieLet11_1_5QNode_Bool_2_bufchan_buf;
  assign lizzieLet11_1_5QNode_Bool_2_bufchan_r = (! lizzieLet11_1_5QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_5QNode_Bool_2_argbuf_d = (lizzieLet11_1_5QNode_Bool_2_bufchan_buf[0] ? lizzieLet11_1_5QNode_Bool_2_bufchan_buf :
                                                 lizzieLet11_1_5QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_5QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_5QNode_Bool_2_argbuf_r && lizzieLet11_1_5QNode_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_5QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_5QNode_Bool_2_argbuf_r) && (! lizzieLet11_1_5QNode_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_5QNode_Bool_2_bufchan_buf <= lizzieLet11_1_5QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet11_1_5QVal_Bool,MyDTBool_Bool) > (lizzieLet11_1_5QVal_Bool_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet11_1_5QVal_Bool_bufchan_d;
  logic lizzieLet11_1_5QVal_Bool_bufchan_r;
  assign lizzieLet11_1_5QVal_Bool_r = ((! lizzieLet11_1_5QVal_Bool_bufchan_d[0]) || lizzieLet11_1_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_5QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_5QVal_Bool_r)
        lizzieLet11_1_5QVal_Bool_bufchan_d <= lizzieLet11_1_5QVal_Bool_d;
  MyDTBool_Bool_t lizzieLet11_1_5QVal_Bool_bufchan_buf;
  assign lizzieLet11_1_5QVal_Bool_bufchan_r = (! lizzieLet11_1_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_5QVal_Bool_1_argbuf_d = (lizzieLet11_1_5QVal_Bool_bufchan_buf[0] ? lizzieLet11_1_5QVal_Bool_bufchan_buf :
                                                lizzieLet11_1_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_5QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_5QVal_Bool_1_argbuf_r && lizzieLet11_1_5QVal_Bool_bufchan_buf[0]))
        lizzieLet11_1_5QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_5QVal_Bool_1_argbuf_r) && (! lizzieLet11_1_5QVal_Bool_bufchan_buf[0])))
        lizzieLet11_1_5QVal_Bool_bufchan_buf <= lizzieLet11_1_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet11_1_6,QTree_Bool) (sc_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(lizzieLet11_1_6QNone_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet11_1_6QVal_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet11_1_6QNode_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet11_1_6QError_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet11_1_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet11_1_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet11_1_6QNone_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                        sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet11_1_6QVal_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                       sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet11_1_6QNode_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                        sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet11_1_6QError_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                         sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet11_1_6QError_Bool_r,
                                                              lizzieLet11_1_6QNode_Bool_r,
                                                              lizzieLet11_1_6QVal_Bool_r,
                                                              lizzieLet11_1_6QNone_Bool_r}));
  assign lizzieLet11_1_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet11_1_6QError_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet11_1_6QError_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QError_Bool_bufchan_d;
  logic lizzieLet11_1_6QError_Bool_bufchan_r;
  assign lizzieLet11_1_6QError_Bool_r = ((! lizzieLet11_1_6QError_Bool_bufchan_d[0]) || lizzieLet11_1_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_6QError_Bool_r)
        lizzieLet11_1_6QError_Bool_bufchan_d <= lizzieLet11_1_6QError_Bool_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QError_Bool_bufchan_buf;
  assign lizzieLet11_1_6QError_Bool_bufchan_r = (! lizzieLet11_1_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_6QError_Bool_1_argbuf_d = (lizzieLet11_1_6QError_Bool_bufchan_buf[0] ? lizzieLet11_1_6QError_Bool_bufchan_buf :
                                                  lizzieLet11_1_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_6QError_Bool_1_argbuf_r && lizzieLet11_1_6QError_Bool_bufchan_buf[0]))
        lizzieLet11_1_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_6QError_Bool_1_argbuf_r) && (! lizzieLet11_1_6QError_Bool_bufchan_buf[0])))
        lizzieLet11_1_6QError_Bool_bufchan_buf <= lizzieLet11_1_6QError_Bool_bufchan_d;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool3) : [(lizzieLet11_1_6QNode_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (lizzieLet11_1_5QNode_Bool_1,MyDTBool_Bool),
                                                 (lizzieLet11_1_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                 (lizzieLet11_1_7QNode_Bool_1,MyBool),
                                                 (q1acF_destruct,Pointer_QTree_Bool),
                                                 (q2acG_destruct,Pointer_QTree_Bool),
                                                 (q3acH_destruct,Pointer_QTree_Bool)] > (lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_d  = \Lcall_map''_map''_Bool_Bool_Bool3_dc ((& {lizzieLet11_1_6QNode_Bool_d[0],
                                                                                                                                                                                                                             lizzieLet11_1_5QNode_Bool_1_d[0],
                                                                                                                                                                                                                             lizzieLet11_1_3QNode_Bool_1_d[0],
                                                                                                                                                                                                                             lizzieLet11_1_7QNode_Bool_1_d[0],
                                                                                                                                                                                                                             q1acF_destruct_d[0],
                                                                                                                                                                                                                             q2acG_destruct_d[0],
                                                                                                                                                                                                                             q3acH_destruct_d[0]}), lizzieLet11_1_6QNode_Bool_d, lizzieLet11_1_5QNode_Bool_1_d, lizzieLet11_1_3QNode_Bool_1_d, lizzieLet11_1_7QNode_Bool_1_d, q1acF_destruct_d, q2acG_destruct_d, q3acH_destruct_d);
  assign {lizzieLet11_1_6QNode_Bool_r,
          lizzieLet11_1_5QNode_Bool_1_r,
          lizzieLet11_1_3QNode_Bool_1_r,
          lizzieLet11_1_7QNode_Bool_1_r,
          q1acF_destruct_r,
          q2acG_destruct_r,
          q3acH_destruct_r} = {7 {(\lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_r  && \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet15_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  logic \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r ;
  assign \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_r  = ((! \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d [0]) || \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= {68'd0,
                                                                                                                                                                                         1'd0};
    else
      if (\lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_r )
        \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf ;
  assign \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r  = (! \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]);
  assign lizzieLet15_1_argbuf_d = (\lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0] ? \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  :
                                   \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= {68'd0,
                                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]))
        \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= {68'd0,
                                                                                                                                                                                             1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0])))
        \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= \lizzieLet11_1_6QNode_Bool_1lizzieLet11_1_5QNode_Bool_1lizzieLet11_1_3QNode_Bool_1lizzieLet11_1_7QNode_Bool_1q1acF_1q2acG_1q3acH_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet11_1_6QNone_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet11_1_6QNone_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QNone_Bool_bufchan_d;
  logic lizzieLet11_1_6QNone_Bool_bufchan_r;
  assign lizzieLet11_1_6QNone_Bool_r = ((! lizzieLet11_1_6QNone_Bool_bufchan_d[0]) || lizzieLet11_1_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_6QNone_Bool_r)
        lizzieLet11_1_6QNone_Bool_bufchan_d <= lizzieLet11_1_6QNone_Bool_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet11_1_6QNone_Bool_bufchan_buf;
  assign lizzieLet11_1_6QNone_Bool_bufchan_r = (! lizzieLet11_1_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_6QNone_Bool_1_argbuf_d = (lizzieLet11_1_6QNone_Bool_bufchan_buf[0] ? lizzieLet11_1_6QNone_Bool_bufchan_buf :
                                                 lizzieLet11_1_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_6QNone_Bool_1_argbuf_r && lizzieLet11_1_6QNone_Bool_bufchan_buf[0]))
        lizzieLet11_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_6QNone_Bool_1_argbuf_r) && (! lizzieLet11_1_6QNone_Bool_bufchan_buf[0])))
        lizzieLet11_1_6QNone_Bool_bufchan_buf <= lizzieLet11_1_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet11_1_7,QTree_Bool) (v'acC_goMux_mux,MyBool) > [(_28,MyBool),
                                                                             (lizzieLet11_1_7QVal_Bool,MyBool),
                                                                             (lizzieLet11_1_7QNode_Bool,MyBool),
                                                                             (_27,MyBool)] */
  logic [3:0] \v'acC_goMux_mux_onehotd ;
  always_comb
    if ((lizzieLet11_1_7_d[0] && \v'acC_goMux_mux_d [0]))
      unique case (lizzieLet11_1_7_d[2:1])
        2'd0: \v'acC_goMux_mux_onehotd  = 4'd1;
        2'd1: \v'acC_goMux_mux_onehotd  = 4'd2;
        2'd2: \v'acC_goMux_mux_onehotd  = 4'd4;
        2'd3: \v'acC_goMux_mux_onehotd  = 4'd8;
        default: \v'acC_goMux_mux_onehotd  = 4'd0;
      endcase
    else \v'acC_goMux_mux_onehotd  = 4'd0;
  assign _28_d = {\v'acC_goMux_mux_d [1:1],
                  \v'acC_goMux_mux_onehotd [0]};
  assign lizzieLet11_1_7QVal_Bool_d = {\v'acC_goMux_mux_d [1:1],
                                       \v'acC_goMux_mux_onehotd [1]};
  assign lizzieLet11_1_7QNode_Bool_d = {\v'acC_goMux_mux_d [1:1],
                                        \v'acC_goMux_mux_onehotd [2]};
  assign _27_d = {\v'acC_goMux_mux_d [1:1],
                  \v'acC_goMux_mux_onehotd [3]};
  assign \v'acC_goMux_mux_r  = (| (\v'acC_goMux_mux_onehotd  & {_27_r,
                                                                lizzieLet11_1_7QNode_Bool_r,
                                                                lizzieLet11_1_7QVal_Bool_r,
                                                                _28_r}));
  assign lizzieLet11_1_7_r = \v'acC_goMux_mux_r ;
  
  /* fork (Ty MyBool) : (lizzieLet11_1_7QNode_Bool,MyBool) > [(lizzieLet11_1_7QNode_Bool_1,MyBool),
                                                         (lizzieLet11_1_7QNode_Bool_2,MyBool)] */
  logic [1:0] lizzieLet11_1_7QNode_Bool_emitted;
  logic [1:0] lizzieLet11_1_7QNode_Bool_done;
  assign lizzieLet11_1_7QNode_Bool_1_d = {lizzieLet11_1_7QNode_Bool_d[1:1],
                                          (lizzieLet11_1_7QNode_Bool_d[0] && (! lizzieLet11_1_7QNode_Bool_emitted[0]))};
  assign lizzieLet11_1_7QNode_Bool_2_d = {lizzieLet11_1_7QNode_Bool_d[1:1],
                                          (lizzieLet11_1_7QNode_Bool_d[0] && (! lizzieLet11_1_7QNode_Bool_emitted[1]))};
  assign lizzieLet11_1_7QNode_Bool_done = (lizzieLet11_1_7QNode_Bool_emitted | ({lizzieLet11_1_7QNode_Bool_2_d[0],
                                                                                 lizzieLet11_1_7QNode_Bool_1_d[0]} & {lizzieLet11_1_7QNode_Bool_2_r,
                                                                                                                      lizzieLet11_1_7QNode_Bool_1_r}));
  assign lizzieLet11_1_7QNode_Bool_r = (& lizzieLet11_1_7QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_7QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_7QNode_Bool_emitted <= (lizzieLet11_1_7QNode_Bool_r ? 2'd0 :
                                            lizzieLet11_1_7QNode_Bool_done);
  
  /* buf (Ty MyBool) : (lizzieLet11_1_7QNode_Bool_2,MyBool) > (lizzieLet11_1_7QNode_Bool_2_argbuf,MyBool) */
  MyBool_t lizzieLet11_1_7QNode_Bool_2_bufchan_d;
  logic lizzieLet11_1_7QNode_Bool_2_bufchan_r;
  assign lizzieLet11_1_7QNode_Bool_2_r = ((! lizzieLet11_1_7QNode_Bool_2_bufchan_d[0]) || lizzieLet11_1_7QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_7QNode_Bool_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet11_1_7QNode_Bool_2_r)
        lizzieLet11_1_7QNode_Bool_2_bufchan_d <= lizzieLet11_1_7QNode_Bool_2_d;
  MyBool_t lizzieLet11_1_7QNode_Bool_2_bufchan_buf;
  assign lizzieLet11_1_7QNode_Bool_2_bufchan_r = (! lizzieLet11_1_7QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_7QNode_Bool_2_argbuf_d = (lizzieLet11_1_7QNode_Bool_2_bufchan_buf[0] ? lizzieLet11_1_7QNode_Bool_2_bufchan_buf :
                                                 lizzieLet11_1_7QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_7QNode_Bool_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet11_1_7QNode_Bool_2_argbuf_r && lizzieLet11_1_7QNode_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_7QNode_Bool_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet11_1_7QNode_Bool_2_argbuf_r) && (! lizzieLet11_1_7QNode_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_7QNode_Bool_2_bufchan_buf <= lizzieLet11_1_7QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyBool) : (lizzieLet11_1_7QVal_Bool,MyBool) > (lizzieLet11_1_7QVal_Bool_1_argbuf,MyBool) */
  MyBool_t lizzieLet11_1_7QVal_Bool_bufchan_d;
  logic lizzieLet11_1_7QVal_Bool_bufchan_r;
  assign lizzieLet11_1_7QVal_Bool_r = ((! lizzieLet11_1_7QVal_Bool_bufchan_d[0]) || lizzieLet11_1_7QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_7QVal_Bool_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet11_1_7QVal_Bool_r)
        lizzieLet11_1_7QVal_Bool_bufchan_d <= lizzieLet11_1_7QVal_Bool_d;
  MyBool_t lizzieLet11_1_7QVal_Bool_bufchan_buf;
  assign lizzieLet11_1_7QVal_Bool_bufchan_r = (! lizzieLet11_1_7QVal_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_7QVal_Bool_1_argbuf_d = (lizzieLet11_1_7QVal_Bool_bufchan_buf[0] ? lizzieLet11_1_7QVal_Bool_bufchan_buf :
                                                lizzieLet11_1_7QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet11_1_7QVal_Bool_1_argbuf_r && lizzieLet11_1_7QVal_Bool_bufchan_buf[0]))
        lizzieLet11_1_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet11_1_7QVal_Bool_1_argbuf_r) && (! lizzieLet11_1_7QVal_Bool_bufchan_buf[0])))
        lizzieLet11_1_7QVal_Bool_bufchan_buf <= lizzieLet11_1_7QVal_Bool_bufchan_d;
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool0) : (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) > [(es_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_2_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_3_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_6_destruct,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted;
  logic [3:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_done;
  assign es_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[19:4],
                            (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[0]))};
  assign es_2_2_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[35:20],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[1]))};
  assign es_3_3_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[51:36],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[67:52],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[3]))};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_done = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted | ({sc_0_6_destruct_d[0],
                                                                                                                       es_3_3_destruct_d[0],
                                                                                                                       es_2_2_destruct_d[0],
                                                                                                                       es_1_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                                                              es_3_3_destruct_r,
                                                                                                                                              es_2_2_destruct_r,
                                                                                                                                              es_1_destruct_r}));
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_r = (& lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted <= 4'd0;
    else
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_emitted <= (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_r ? 4'd0 :
                                                               lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool1) : (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_3_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_5_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZacJ_4_destruct,MyDTBool_Bool),
                                                                                                                               (gacK_4_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1acO_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2acM_4_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted;
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_done;
  assign es_2_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[19:4],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[35:20],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[51:36],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[2]))};
  assign isZacJ_4_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[3]));
  assign gacK_4_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[4]));
  assign q1acO_3_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[67:52],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[5]))};
  assign m2acM_4_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[83:68],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[6]))};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_done = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted | ({m2acM_4_destruct_d[0],
                                                                                                                       q1acO_3_destruct_d[0],
                                                                                                                       gacK_4_destruct_d[0],
                                                                                                                       isZacJ_4_destruct_d[0],
                                                                                                                       sc_0_5_destruct_d[0],
                                                                                                                       es_3_2_destruct_d[0],
                                                                                                                       es_2_1_destruct_d[0]} & {m2acM_4_destruct_r,
                                                                                                                                                q1acO_3_destruct_r,
                                                                                                                                                gacK_4_destruct_r,
                                                                                                                                                isZacJ_4_destruct_r,
                                                                                                                                                sc_0_5_destruct_r,
                                                                                                                                                es_3_2_destruct_r,
                                                                                                                                                es_2_1_destruct_r}));
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_r = (& lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted <= 7'd0;
    else
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_emitted <= (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_r ? 7'd0 :
                                                               lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool2) : (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) > [(es_3_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_4_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZacJ_3_destruct,MyDTBool_Bool),
                                                                                                                               (gacK_3_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1acO_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2acM_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (q2acP_2_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted;
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_done;
  assign es_3_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[19:4],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[35:20],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[1]))};
  assign isZacJ_3_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[2]));
  assign gacK_3_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[3]));
  assign q1acO_2_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[51:36],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[4]))};
  assign m2acM_3_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[67:52],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[5]))};
  assign q2acP_2_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[83:68],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[6]))};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_done = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted | ({q2acP_2_destruct_d[0],
                                                                                                                       m2acM_3_destruct_d[0],
                                                                                                                       q1acO_2_destruct_d[0],
                                                                                                                       gacK_3_destruct_d[0],
                                                                                                                       isZacJ_3_destruct_d[0],
                                                                                                                       sc_0_4_destruct_d[0],
                                                                                                                       es_3_1_destruct_d[0]} & {q2acP_2_destruct_r,
                                                                                                                                                m2acM_3_destruct_r,
                                                                                                                                                q1acO_2_destruct_r,
                                                                                                                                                gacK_3_destruct_r,
                                                                                                                                                isZacJ_3_destruct_r,
                                                                                                                                                sc_0_4_destruct_r,
                                                                                                                                                es_3_1_destruct_r}));
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_r = (& lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted <= 7'd0;
    else
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_emitted <= (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_r ? 7'd0 :
                                                               lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool3) : (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) > [(sc_0_3_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZacJ_2_destruct,MyDTBool_Bool),
                                                                                                                               (gacK_2_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1acO_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2acM_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (q2acP_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (q3acQ_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted;
  logic [6:0] lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_done;
  assign sc_0_3_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[19:4],
                              (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[0]))};
  assign isZacJ_2_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[1]));
  assign gacK_2_destruct_d = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[2]));
  assign q1acO_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[35:20],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[3]))};
  assign m2acM_2_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[51:36],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[4]))};
  assign q2acP_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[67:52],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[5]))};
  assign q3acQ_1_destruct_d = {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[83:68],
                               (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[6]))};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_done = (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted | ({q3acQ_1_destruct_d[0],
                                                                                                                       q2acP_1_destruct_d[0],
                                                                                                                       m2acM_2_destruct_d[0],
                                                                                                                       q1acO_1_destruct_d[0],
                                                                                                                       gacK_2_destruct_d[0],
                                                                                                                       isZacJ_2_destruct_d[0],
                                                                                                                       sc_0_3_destruct_d[0]} & {q3acQ_1_destruct_r,
                                                                                                                                                q2acP_1_destruct_r,
                                                                                                                                                m2acM_2_destruct_r,
                                                                                                                                                q1acO_1_destruct_r,
                                                                                                                                                gacK_2_destruct_r,
                                                                                                                                                isZacJ_2_destruct_r,
                                                                                                                                                sc_0_3_destruct_r}));
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_r = (& lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted <= 7'd0;
    else
      lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_emitted <= (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_r ? 7'd0 :
                                                               lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_done);
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet20_2,CTkron_kron_Bool_Bool_Bool) (lizzieLet20_1,CTkron_kron_Bool_Bool_Bool) > [(_26,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool)] */
  logic [4:0] lizzieLet20_1_onehotd;
  always_comb
    if ((lizzieLet20_2_d[0] && lizzieLet20_1_d[0]))
      unique case (lizzieLet20_2_d[3:1])
        3'd0: lizzieLet20_1_onehotd = 5'd1;
        3'd1: lizzieLet20_1_onehotd = 5'd2;
        3'd2: lizzieLet20_1_onehotd = 5'd4;
        3'd3: lizzieLet20_1_onehotd = 5'd8;
        3'd4: lizzieLet20_1_onehotd = 5'd16;
        default: lizzieLet20_1_onehotd = 5'd0;
      endcase
    else lizzieLet20_1_onehotd = 5'd0;
  assign _26_d = {lizzieLet20_1_d[83:1], lizzieLet20_1_onehotd[0]};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_d = {lizzieLet20_1_d[83:1],
                                                           lizzieLet20_1_onehotd[1]};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_d = {lizzieLet20_1_d[83:1],
                                                           lizzieLet20_1_onehotd[2]};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_d = {lizzieLet20_1_d[83:1],
                                                           lizzieLet20_1_onehotd[3]};
  assign lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_d = {lizzieLet20_1_d[83:1],
                                                           lizzieLet20_1_onehotd[4]};
  assign lizzieLet20_1_r = (| (lizzieLet20_1_onehotd & {lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                        lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                        lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                        lizzieLet20_1Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                        _26_r}));
  assign lizzieLet20_2_r = lizzieLet20_1_r;
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty Go) : (lizzieLet20_3,CTkron_kron_Bool_Bool_Bool) (go_10_goMux_data,Go) > [(_25,Go),
                                                                                    (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3,Go),
                                                                                    (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2,Go),
                                                                                    (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1,Go),
                                                                                    (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0,Go)] */
  logic [4:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet20_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet20_3_d[3:1])
        3'd0: go_10_goMux_data_onehotd = 5'd1;
        3'd1: go_10_goMux_data_onehotd = 5'd2;
        3'd2: go_10_goMux_data_onehotd = 5'd4;
        3'd3: go_10_goMux_data_onehotd = 5'd8;
        3'd4: go_10_goMux_data_onehotd = 5'd16;
        default: go_10_goMux_data_onehotd = 5'd0;
      endcase
    else go_10_goMux_data_onehotd = 5'd0;
  assign _25_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_d = go_10_goMux_data_onehotd[3];
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_d = go_10_goMux_data_onehotd[4];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                              lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                              lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                              lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                              _25_r}));
  assign lizzieLet20_3_r = go_10_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0,Go) > (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf,Go) */
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_r = ((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d[0]) || lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_r)
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_d;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r = (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]);
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d = (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0] ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf :
                                                                    lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r && lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r) && (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0])))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1,Go) > (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf,Go) */
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_r = ((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d[0]) || lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_r)
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_d;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r = (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]);
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d = (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0] ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf :
                                                                    lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r && lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r) && (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0])))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2,Go) > (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf,Go) */
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_r = ((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d[0]) || lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_r)
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_d;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r = (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]);
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d = (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0] ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf :
                                                                    lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r && lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r) && (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0])))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3,Go) > (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf,Go) */
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  logic lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_r = ((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d[0]) || lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= 1'd0;
    else
      if (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_r)
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_d;
  Go_t lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf;
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r = (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]);
  assign lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d = (lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0] ? lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf :
                                                                    lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r && lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r) && (! lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0])))
        lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= lizzieLet20_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet20_4,CTkron_kron_Bool_Bool_Bool) (srtarg_0_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet20_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet20_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                                         srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                                  lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                                  lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                                  lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                                  lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_r}));
  assign lizzieLet20_4_r = srtarg_0_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0,Pointer_QTree_Bool),
                          (es_1_destruct,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_3_destruct,Pointer_QTree_Bool)] > (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) */
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_d[0],
                                                                                                              es_1_destruct_d[0],
                                                                                                              es_2_2_destruct_d[0],
                                                                                                              es_3_3_destruct_d[0]}), lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_d, es_1_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_r,
          es_1_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) > (lizzieLet24_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_r = ((! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d[0]) || lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                                   1'd0};
    else
      if (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_r)
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_d;
  QTree_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r = (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0] ? lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf :
                                   lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                                     1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0]))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                                       1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0])))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool0) : [(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                               (es_2_1_destruct,Pointer_QTree_Bool),
                                               (es_3_2_destruct,Pointer_QTree_Bool),
                                               (sc_0_5_destruct,Pointer_CTkron_kron_Bool_Bool_Bool)] > (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d = Lcall_kron_kron_Bool_Bool_Bool0_dc((& {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_d[0],
                                                                                                                                                          es_2_1_destruct_d[0],
                                                                                                                                                          es_3_2_destruct_d[0],
                                                                                                                                                          sc_0_5_destruct_d[0]}), lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_d, es_2_1_destruct_d, es_3_2_destruct_d, sc_0_5_destruct_d);
  assign {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_r,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_5_destruct_r} = {4 {(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) > (lizzieLet23_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r = ((! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d[0]) || lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= {83'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r)
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r = (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0] ? lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf :
                                   lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= {83'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= {83'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0])))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool1) : [(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                               (es_3_1_destruct,Pointer_QTree_Bool),
                                               (sc_0_4_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (isZacJ_3_1,MyDTBool_Bool),
                                               (gacK_3_1,MyDTBool_Bool_Bool),
                                               (q1acO_2_destruct,Pointer_QTree_Bool),
                                               (m2acM_3_1,Pointer_QTree_Bool)] > (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_d = Lcall_kron_kron_Bool_Bool_Bool1_dc((& {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_d[0],
                                                                                                                                                                                      es_3_1_destruct_d[0],
                                                                                                                                                                                      sc_0_4_destruct_d[0],
                                                                                                                                                                                      isZacJ_3_1_d[0],
                                                                                                                                                                                      gacK_3_1_d[0],
                                                                                                                                                                                      q1acO_2_destruct_d[0],
                                                                                                                                                                                      m2acM_3_1_d[0]}), lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_d, es_3_1_destruct_d, sc_0_4_destruct_d, isZacJ_3_1_d, gacK_3_1_d, q1acO_2_destruct_d, m2acM_3_1_d);
  assign {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_r,
          es_3_1_destruct_r,
          sc_0_4_destruct_r,
          isZacJ_3_1_r,
          gacK_3_1_r,
          q1acO_2_destruct_r,
          m2acM_3_1_r} = {7 {(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) > (lizzieLet22_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_r = ((! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d[0]) || lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= {83'd0,
                                                                                                                                                      1'd0};
    else
      if (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_r)
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r = (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0] ? lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf :
                                   lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= {83'd0,
                                                                                                                                                        1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= {83'd0,
                                                                                                                                                          1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0])))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZacJ_3_1gacK_3_1q1acO_2_1m2acM_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool2) : [(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                               (sc_0_3_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (isZacJ_2_1,MyDTBool_Bool),
                                               (gacK_2_1,MyDTBool_Bool_Bool),
                                               (q1acO_1_destruct,Pointer_QTree_Bool),
                                               (m2acM_2_1,Pointer_QTree_Bool),
                                               (q2acP_1_destruct,Pointer_QTree_Bool)] > (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_d = Lcall_kron_kron_Bool_Bool_Bool2_dc((& {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_d[0],
                                                                                                                                                                                       sc_0_3_destruct_d[0],
                                                                                                                                                                                       isZacJ_2_1_d[0],
                                                                                                                                                                                       gacK_2_1_d[0],
                                                                                                                                                                                       q1acO_1_destruct_d[0],
                                                                                                                                                                                       m2acM_2_1_d[0],
                                                                                                                                                                                       q2acP_1_destruct_d[0]}), lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_d, sc_0_3_destruct_d, isZacJ_2_1_d, gacK_2_1_d, q1acO_1_destruct_d, m2acM_2_1_d, q2acP_1_destruct_d);
  assign {lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_r,
          sc_0_3_destruct_r,
          isZacJ_2_1_r,
          gacK_2_1_r,
          q1acO_1_destruct_r,
          m2acM_2_1_r,
          q2acP_1_destruct_r} = {7 {(lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) > (lizzieLet21_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  logic lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_r = ((! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d[0]) || lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= {83'd0,
                                                                                                                                                       1'd0};
    else
      if (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_r)
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf;
  assign lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r = (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0] ? lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf :
                                   lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= {83'd0,
                                                                                                                                                         1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= {83'd0,
                                                                                                                                                           1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0])))
        lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= lizzieLet20_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZacJ_2_1gacK_2_1q1acO_1_1m2acM_2_1q2acP_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                                  (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted;
  logic [1:0] lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_done;
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d = {lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d[16:1],
                                                                              (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d[0] && (! lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted[0]))};
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d = {lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d[16:1],
                                                                              (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_d[0] && (! lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted[1]))};
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_done = (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted | ({lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d[0],
                                                                                                                   lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r,
                                                                                                                                                                                            lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_r = (& lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted <= 2'd0;
    else
      lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_emitted <= (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_r ? 2'd0 :
                                                             lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_kron_kron_Bool_Bool_Bool_goConst,Go) */
  assign call_kron_kron_Bool_Bool_Bool_goConst_d = lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r = call_kron_kron_Bool_Bool_Bool_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (kron_kron_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r = ((! lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                                    1'd0};
    else
      if (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r)
        lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign kron_kron_Bool_Bool_Bool_resbuf_d = (lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf :
                                              lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                      1'd0};
    else
      if ((kron_kron_Bool_Bool_Bool_resbuf_r && lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                        1'd0};
      else if (((! kron_kron_Bool_Bool_Bool_resbuf_r) && (! lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet20_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool0) : (lizzieLet25_1Lcall_main_mask_Bool0,CTmain_mask_Bool) > [(es_1_1_destruct,Pointer_QTree_Bool),
                                                                                                 (es_2_4_destruct,Pointer_QTree_Bool),
                                                                                                 (es_3_6_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_10_destruct,Pointer_CTmain_mask_Bool)] */
  logic [3:0] lizzieLet25_1Lcall_main_mask_Bool0_emitted;
  logic [3:0] lizzieLet25_1Lcall_main_mask_Bool0_done;
  assign es_1_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool0_d[19:4],
                              (lizzieLet25_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool0_emitted[0]))};
  assign es_2_4_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool0_d[35:20],
                              (lizzieLet25_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool0_emitted[1]))};
  assign es_3_6_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool0_d[51:36],
                              (lizzieLet25_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool0_emitted[2]))};
  assign sc_0_10_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool0_d[67:52],
                               (lizzieLet25_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool0_emitted[3]))};
  assign lizzieLet25_1Lcall_main_mask_Bool0_done = (lizzieLet25_1Lcall_main_mask_Bool0_emitted | ({sc_0_10_destruct_d[0],
                                                                                                   es_3_6_destruct_d[0],
                                                                                                   es_2_4_destruct_d[0],
                                                                                                   es_1_1_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                            es_3_6_destruct_r,
                                                                                                                            es_2_4_destruct_r,
                                                                                                                            es_1_1_destruct_r}));
  assign lizzieLet25_1Lcall_main_mask_Bool0_r = (& lizzieLet25_1Lcall_main_mask_Bool0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1Lcall_main_mask_Bool0_emitted <= 4'd0;
    else
      lizzieLet25_1Lcall_main_mask_Bool0_emitted <= (lizzieLet25_1Lcall_main_mask_Bool0_r ? 4'd0 :
                                                     lizzieLet25_1Lcall_main_mask_Bool0_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool1) : (lizzieLet25_1Lcall_main_mask_Bool1,CTmain_mask_Bool) > [(es_2_3_destruct,Pointer_QTree_Bool),
                                                                                                 (es_3_5_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_9_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1acp_3_destruct,Pointer_QTree_Bool),
                                                                                                 (q1ack_3_destruct,Pointer_MaskQTree)] */
  logic [4:0] lizzieLet25_1Lcall_main_mask_Bool1_emitted;
  logic [4:0] lizzieLet25_1Lcall_main_mask_Bool1_done;
  assign es_2_3_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool1_d[19:4],
                              (lizzieLet25_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool1_emitted[0]))};
  assign es_3_5_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool1_d[35:20],
                              (lizzieLet25_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool1_emitted[1]))};
  assign sc_0_9_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool1_d[51:36],
                              (lizzieLet25_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool1_emitted[2]))};
  assign t1acp_3_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool1_d[67:52],
                               (lizzieLet25_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool1_emitted[3]))};
  assign q1ack_3_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool1_d[83:68],
                               (lizzieLet25_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool1_emitted[4]))};
  assign lizzieLet25_1Lcall_main_mask_Bool1_done = (lizzieLet25_1Lcall_main_mask_Bool1_emitted | ({q1ack_3_destruct_d[0],
                                                                                                   t1acp_3_destruct_d[0],
                                                                                                   sc_0_9_destruct_d[0],
                                                                                                   es_3_5_destruct_d[0],
                                                                                                   es_2_3_destruct_d[0]} & {q1ack_3_destruct_r,
                                                                                                                            t1acp_3_destruct_r,
                                                                                                                            sc_0_9_destruct_r,
                                                                                                                            es_3_5_destruct_r,
                                                                                                                            es_2_3_destruct_r}));
  assign lizzieLet25_1Lcall_main_mask_Bool1_r = (& lizzieLet25_1Lcall_main_mask_Bool1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1Lcall_main_mask_Bool1_emitted <= 5'd0;
    else
      lizzieLet25_1Lcall_main_mask_Bool1_emitted <= (lizzieLet25_1Lcall_main_mask_Bool1_r ? 5'd0 :
                                                     lizzieLet25_1Lcall_main_mask_Bool1_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool2) : (lizzieLet25_1Lcall_main_mask_Bool2,CTmain_mask_Bool) > [(es_3_4_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_8_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1acp_2_destruct,Pointer_QTree_Bool),
                                                                                                 (q1ack_2_destruct,Pointer_MaskQTree),
                                                                                                 (t2acq_2_destruct,Pointer_QTree_Bool),
                                                                                                 (q2acl_2_destruct,Pointer_MaskQTree)] */
  logic [5:0] lizzieLet25_1Lcall_main_mask_Bool2_emitted;
  logic [5:0] lizzieLet25_1Lcall_main_mask_Bool2_done;
  assign es_3_4_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[19:4],
                              (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[0]))};
  assign sc_0_8_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[35:20],
                              (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[1]))};
  assign t1acp_2_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[51:36],
                               (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[2]))};
  assign q1ack_2_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[67:52],
                               (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[3]))};
  assign t2acq_2_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[83:68],
                               (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[4]))};
  assign q2acl_2_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool2_d[99:84],
                               (lizzieLet25_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool2_emitted[5]))};
  assign lizzieLet25_1Lcall_main_mask_Bool2_done = (lizzieLet25_1Lcall_main_mask_Bool2_emitted | ({q2acl_2_destruct_d[0],
                                                                                                   t2acq_2_destruct_d[0],
                                                                                                   q1ack_2_destruct_d[0],
                                                                                                   t1acp_2_destruct_d[0],
                                                                                                   sc_0_8_destruct_d[0],
                                                                                                   es_3_4_destruct_d[0]} & {q2acl_2_destruct_r,
                                                                                                                            t2acq_2_destruct_r,
                                                                                                                            q1ack_2_destruct_r,
                                                                                                                            t1acp_2_destruct_r,
                                                                                                                            sc_0_8_destruct_r,
                                                                                                                            es_3_4_destruct_r}));
  assign lizzieLet25_1Lcall_main_mask_Bool2_r = (& lizzieLet25_1Lcall_main_mask_Bool2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1Lcall_main_mask_Bool2_emitted <= 6'd0;
    else
      lizzieLet25_1Lcall_main_mask_Bool2_emitted <= (lizzieLet25_1Lcall_main_mask_Bool2_r ? 6'd0 :
                                                     lizzieLet25_1Lcall_main_mask_Bool2_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool3) : (lizzieLet25_1Lcall_main_mask_Bool3,CTmain_mask_Bool) > [(sc_0_7_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1acp_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q1ack_1_destruct,Pointer_MaskQTree),
                                                                                                 (t2acq_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q2acl_1_destruct,Pointer_MaskQTree),
                                                                                                 (t3acr_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q3acm_1_destruct,Pointer_MaskQTree)] */
  logic [6:0] lizzieLet25_1Lcall_main_mask_Bool3_emitted;
  logic [6:0] lizzieLet25_1Lcall_main_mask_Bool3_done;
  assign sc_0_7_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[19:4],
                              (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[0]))};
  assign t1acp_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[35:20],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[1]))};
  assign q1ack_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[51:36],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[2]))};
  assign t2acq_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[67:52],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[3]))};
  assign q2acl_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[83:68],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[4]))};
  assign t3acr_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[99:84],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[5]))};
  assign q3acm_1_destruct_d = {lizzieLet25_1Lcall_main_mask_Bool3_d[115:100],
                               (lizzieLet25_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet25_1Lcall_main_mask_Bool3_emitted[6]))};
  assign lizzieLet25_1Lcall_main_mask_Bool3_done = (lizzieLet25_1Lcall_main_mask_Bool3_emitted | ({q3acm_1_destruct_d[0],
                                                                                                   t3acr_1_destruct_d[0],
                                                                                                   q2acl_1_destruct_d[0],
                                                                                                   t2acq_1_destruct_d[0],
                                                                                                   q1ack_1_destruct_d[0],
                                                                                                   t1acp_1_destruct_d[0],
                                                                                                   sc_0_7_destruct_d[0]} & {q3acm_1_destruct_r,
                                                                                                                            t3acr_1_destruct_r,
                                                                                                                            q2acl_1_destruct_r,
                                                                                                                            t2acq_1_destruct_r,
                                                                                                                            q1ack_1_destruct_r,
                                                                                                                            t1acp_1_destruct_r,
                                                                                                                            sc_0_7_destruct_r}));
  assign lizzieLet25_1Lcall_main_mask_Bool3_r = (& lizzieLet25_1Lcall_main_mask_Bool3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1Lcall_main_mask_Bool3_emitted <= 7'd0;
    else
      lizzieLet25_1Lcall_main_mask_Bool3_emitted <= (lizzieLet25_1Lcall_main_mask_Bool3_r ? 7'd0 :
                                                     lizzieLet25_1Lcall_main_mask_Bool3_done);
  
  /* demux (Ty CTmain_mask_Bool,
       Ty CTmain_mask_Bool) : (lizzieLet25_2,CTmain_mask_Bool) (lizzieLet25_1,CTmain_mask_Bool) > [(_24,CTmain_mask_Bool),
                                                                                                   (lizzieLet25_1Lcall_main_mask_Bool3,CTmain_mask_Bool),
                                                                                                   (lizzieLet25_1Lcall_main_mask_Bool2,CTmain_mask_Bool),
                                                                                                   (lizzieLet25_1Lcall_main_mask_Bool1,CTmain_mask_Bool),
                                                                                                   (lizzieLet25_1Lcall_main_mask_Bool0,CTmain_mask_Bool)] */
  logic [4:0] lizzieLet25_1_onehotd;
  always_comb
    if ((lizzieLet25_2_d[0] && lizzieLet25_1_d[0]))
      unique case (lizzieLet25_2_d[3:1])
        3'd0: lizzieLet25_1_onehotd = 5'd1;
        3'd1: lizzieLet25_1_onehotd = 5'd2;
        3'd2: lizzieLet25_1_onehotd = 5'd4;
        3'd3: lizzieLet25_1_onehotd = 5'd8;
        3'd4: lizzieLet25_1_onehotd = 5'd16;
        default: lizzieLet25_1_onehotd = 5'd0;
      endcase
    else lizzieLet25_1_onehotd = 5'd0;
  assign _24_d = {lizzieLet25_1_d[115:1], lizzieLet25_1_onehotd[0]};
  assign lizzieLet25_1Lcall_main_mask_Bool3_d = {lizzieLet25_1_d[115:1],
                                                 lizzieLet25_1_onehotd[1]};
  assign lizzieLet25_1Lcall_main_mask_Bool2_d = {lizzieLet25_1_d[115:1],
                                                 lizzieLet25_1_onehotd[2]};
  assign lizzieLet25_1Lcall_main_mask_Bool1_d = {lizzieLet25_1_d[115:1],
                                                 lizzieLet25_1_onehotd[3]};
  assign lizzieLet25_1Lcall_main_mask_Bool0_d = {lizzieLet25_1_d[115:1],
                                                 lizzieLet25_1_onehotd[4]};
  assign lizzieLet25_1_r = (| (lizzieLet25_1_onehotd & {lizzieLet25_1Lcall_main_mask_Bool0_r,
                                                        lizzieLet25_1Lcall_main_mask_Bool1_r,
                                                        lizzieLet25_1Lcall_main_mask_Bool2_r,
                                                        lizzieLet25_1Lcall_main_mask_Bool3_r,
                                                        _24_r}));
  assign lizzieLet25_2_r = lizzieLet25_1_r;
  
  /* demux (Ty CTmain_mask_Bool,
       Ty Go) : (lizzieLet25_3,CTmain_mask_Bool) (go_11_goMux_data,Go) > [(_23,Go),
                                                                          (lizzieLet25_3Lcall_main_mask_Bool3,Go),
                                                                          (lizzieLet25_3Lcall_main_mask_Bool2,Go),
                                                                          (lizzieLet25_3Lcall_main_mask_Bool1,Go),
                                                                          (lizzieLet25_3Lcall_main_mask_Bool0,Go)] */
  logic [4:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet25_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet25_3_d[3:1])
        3'd0: go_11_goMux_data_onehotd = 5'd1;
        3'd1: go_11_goMux_data_onehotd = 5'd2;
        3'd2: go_11_goMux_data_onehotd = 5'd4;
        3'd3: go_11_goMux_data_onehotd = 5'd8;
        3'd4: go_11_goMux_data_onehotd = 5'd16;
        default: go_11_goMux_data_onehotd = 5'd0;
      endcase
    else go_11_goMux_data_onehotd = 5'd0;
  assign _23_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet25_3Lcall_main_mask_Bool3_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet25_3Lcall_main_mask_Bool2_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet25_3Lcall_main_mask_Bool1_d = go_11_goMux_data_onehotd[3];
  assign lizzieLet25_3Lcall_main_mask_Bool0_d = go_11_goMux_data_onehotd[4];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet25_3Lcall_main_mask_Bool0_r,
                                                              lizzieLet25_3Lcall_main_mask_Bool1_r,
                                                              lizzieLet25_3Lcall_main_mask_Bool2_r,
                                                              lizzieLet25_3Lcall_main_mask_Bool3_r,
                                                              _23_r}));
  assign lizzieLet25_3_r = go_11_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_main_mask_Bool0,Go) > (lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d;
  logic lizzieLet25_3Lcall_main_mask_Bool0_bufchan_r;
  assign lizzieLet25_3Lcall_main_mask_Bool0_r = ((! lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d[0]) || lizzieLet25_3Lcall_main_mask_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_main_mask_Bool0_r)
        lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d <= lizzieLet25_3Lcall_main_mask_Bool0_d;
  Go_t lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf;
  assign lizzieLet25_3Lcall_main_mask_Bool0_bufchan_r = (! lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_d = (lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf[0] ? lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf :
                                                          lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_r && lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf[0]))
        lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_r) && (! lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf[0])))
        lizzieLet25_3Lcall_main_mask_Bool0_bufchan_buf <= lizzieLet25_3Lcall_main_mask_Bool0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_main_mask_Bool1,Go) > (lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d;
  logic lizzieLet25_3Lcall_main_mask_Bool1_bufchan_r;
  assign lizzieLet25_3Lcall_main_mask_Bool1_r = ((! lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d[0]) || lizzieLet25_3Lcall_main_mask_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_main_mask_Bool1_r)
        lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d <= lizzieLet25_3Lcall_main_mask_Bool1_d;
  Go_t lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf;
  assign lizzieLet25_3Lcall_main_mask_Bool1_bufchan_r = (! lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_d = (lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf[0] ? lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf :
                                                          lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_r && lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf[0]))
        lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_main_mask_Bool1_1_argbuf_r) && (! lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf[0])))
        lizzieLet25_3Lcall_main_mask_Bool1_bufchan_buf <= lizzieLet25_3Lcall_main_mask_Bool1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_main_mask_Bool2,Go) > (lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d;
  logic lizzieLet25_3Lcall_main_mask_Bool2_bufchan_r;
  assign lizzieLet25_3Lcall_main_mask_Bool2_r = ((! lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d[0]) || lizzieLet25_3Lcall_main_mask_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_main_mask_Bool2_r)
        lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d <= lizzieLet25_3Lcall_main_mask_Bool2_d;
  Go_t lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf;
  assign lizzieLet25_3Lcall_main_mask_Bool2_bufchan_r = (! lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_d = (lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf[0] ? lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf :
                                                          lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_r && lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf[0]))
        lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_main_mask_Bool2_1_argbuf_r) && (! lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf[0])))
        lizzieLet25_3Lcall_main_mask_Bool2_bufchan_buf <= lizzieLet25_3Lcall_main_mask_Bool2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_3Lcall_main_mask_Bool3,Go) > (lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf,Go) */
  Go_t lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d;
  logic lizzieLet25_3Lcall_main_mask_Bool3_bufchan_r;
  assign lizzieLet25_3Lcall_main_mask_Bool3_r = ((! lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d[0]) || lizzieLet25_3Lcall_main_mask_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_3Lcall_main_mask_Bool3_r)
        lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d <= lizzieLet25_3Lcall_main_mask_Bool3_d;
  Go_t lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf;
  assign lizzieLet25_3Lcall_main_mask_Bool3_bufchan_r = (! lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf[0]);
  assign lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_d = (lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf[0] ? lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf :
                                                          lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_r && lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf[0]))
        lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_3Lcall_main_mask_Bool3_1_argbuf_r) && (! lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf[0])))
        lizzieLet25_3Lcall_main_mask_Bool3_bufchan_buf <= lizzieLet25_3Lcall_main_mask_Bool3_bufchan_d;
  
  /* demux (Ty CTmain_mask_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet25_4,CTmain_mask_Bool) (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet25_4Lmain_mask_Boolsbos,Pointer_QTree_Bool),
                                                                                                              (lizzieLet25_4Lcall_main_mask_Bool3,Pointer_QTree_Bool),
                                                                                                              (lizzieLet25_4Lcall_main_mask_Bool2,Pointer_QTree_Bool),
                                                                                                              (lizzieLet25_4Lcall_main_mask_Bool1,Pointer_QTree_Bool),
                                                                                                              (lizzieLet25_4Lcall_main_mask_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet25_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet25_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet25_4Lmain_mask_Boolsbos_d = {srtarg_0_1_goMux_mux_d[16:1],
                                               srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet25_4Lcall_main_mask_Bool3_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet25_4Lcall_main_mask_Bool2_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet25_4Lcall_main_mask_Bool1_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet25_4Lcall_main_mask_Bool0_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet25_4Lcall_main_mask_Bool0_r,
                                                                      lizzieLet25_4Lcall_main_mask_Bool1_r,
                                                                      lizzieLet25_4Lcall_main_mask_Bool2_r,
                                                                      lizzieLet25_4Lcall_main_mask_Bool3_r,
                                                                      lizzieLet25_4Lmain_mask_Boolsbos_r}));
  assign lizzieLet25_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet25_4Lcall_main_mask_Bool0,Pointer_QTree_Bool),
                          (es_1_1_destruct,Pointer_QTree_Bool),
                          (es_2_4_destruct,Pointer_QTree_Bool),
                          (es_3_6_destruct,Pointer_QTree_Bool)] > (lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool,QTree_Bool) */
  assign lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet25_4Lcall_main_mask_Bool0_d[0],
                                                                                                      es_1_1_destruct_d[0],
                                                                                                      es_2_4_destruct_d[0],
                                                                                                      es_3_6_destruct_d[0]}), lizzieLet25_4Lcall_main_mask_Bool0_d, es_1_1_destruct_d, es_2_4_destruct_d, es_3_6_destruct_d);
  assign {lizzieLet25_4Lcall_main_mask_Bool0_r,
          es_1_1_destruct_r,
          es_2_4_destruct_r,
          es_3_6_destruct_r} = {4 {(lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_r && lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool,QTree_Bool) > (lizzieLet29_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d;
  logic lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r;
  assign lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_r = ((! lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d[0]) || lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                           1'd0};
    else
      if (lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_r)
        lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d <= lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_d;
  QTree_Bool_t lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf;
  assign lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_r = (! lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf[0] ? lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf :
                                   lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                             1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf[0]))
        lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                               1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf[0])))
        lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_buf <= lizzieLet25_4Lcall_main_mask_Bool0_1es_1_1_1es_2_4_1es_3_6_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool0) : [(lizzieLet25_4Lcall_main_mask_Bool1,Pointer_QTree_Bool),
                                     (es_2_3_destruct,Pointer_QTree_Bool),
                                     (es_3_5_destruct,Pointer_QTree_Bool),
                                     (sc_0_9_destruct,Pointer_CTmain_mask_Bool)] > (lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0,CTmain_mask_Bool) */
  assign lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_d = Lcall_main_mask_Bool0_dc((& {lizzieLet25_4Lcall_main_mask_Bool1_d[0],
                                                                                                                            es_2_3_destruct_d[0],
                                                                                                                            es_3_5_destruct_d[0],
                                                                                                                            sc_0_9_destruct_d[0]}), lizzieLet25_4Lcall_main_mask_Bool1_d, es_2_3_destruct_d, es_3_5_destruct_d, sc_0_9_destruct_d);
  assign {lizzieLet25_4Lcall_main_mask_Bool1_r,
          es_2_3_destruct_r,
          es_3_5_destruct_r,
          sc_0_9_destruct_r} = {4 {(lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_r && lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0,CTmain_mask_Bool) > (lizzieLet28_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d;
  logic lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_r;
  assign lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_r = ((! lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d[0]) || lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d <= {115'd0,
                                                                                                      1'd0};
    else
      if (lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_r)
        lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d <= lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_d;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf;
  assign lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_r = (! lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf[0] ? lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf :
                                   lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf <= {115'd0,
                                                                                                        1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf[0]))
        lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf <= {115'd0,
                                                                                                          1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf[0])))
        lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_buf <= lizzieLet25_4Lcall_main_mask_Bool1_1es_2_3_1es_3_5_1sc_0_9_1Lcall_main_mask_Bool0_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool1) : [(lizzieLet25_4Lcall_main_mask_Bool2,Pointer_QTree_Bool),
                                     (es_3_4_destruct,Pointer_QTree_Bool),
                                     (sc_0_8_destruct,Pointer_CTmain_mask_Bool),
                                     (t1acp_2_destruct,Pointer_QTree_Bool),
                                     (q1ack_2_destruct,Pointer_MaskQTree)] > (lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1,CTmain_mask_Bool) */
  assign lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_d = Lcall_main_mask_Bool1_dc((& {lizzieLet25_4Lcall_main_mask_Bool2_d[0],
                                                                                                                                      es_3_4_destruct_d[0],
                                                                                                                                      sc_0_8_destruct_d[0],
                                                                                                                                      t1acp_2_destruct_d[0],
                                                                                                                                      q1ack_2_destruct_d[0]}), lizzieLet25_4Lcall_main_mask_Bool2_d, es_3_4_destruct_d, sc_0_8_destruct_d, t1acp_2_destruct_d, q1ack_2_destruct_d);
  assign {lizzieLet25_4Lcall_main_mask_Bool2_r,
          es_3_4_destruct_r,
          sc_0_8_destruct_r,
          t1acp_2_destruct_r,
          q1ack_2_destruct_r} = {5 {(lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_r && lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1,CTmain_mask_Bool) > (lizzieLet27_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d;
  logic lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_r;
  assign lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_r = ((! lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d[0]) || lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d <= {115'd0,
                                                                                                                1'd0};
    else
      if (lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_r)
        lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d <= lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_d;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf;
  assign lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_r = (! lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf[0] ? lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf :
                                   lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf <= {115'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf[0]))
        lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf <= {115'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf[0])))
        lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_buf <= lizzieLet25_4Lcall_main_mask_Bool2_1es_3_4_1sc_0_8_1t1acp_2_1q1ack_2_1Lcall_main_mask_Bool1_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool2) : [(lizzieLet25_4Lcall_main_mask_Bool3,Pointer_QTree_Bool),
                                     (sc_0_7_destruct,Pointer_CTmain_mask_Bool),
                                     (t1acp_1_destruct,Pointer_QTree_Bool),
                                     (q1ack_1_destruct,Pointer_MaskQTree),
                                     (t2acq_1_destruct,Pointer_QTree_Bool),
                                     (q2acl_1_destruct,Pointer_MaskQTree)] > (lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2,CTmain_mask_Bool) */
  assign lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_d = Lcall_main_mask_Bool2_dc((& {lizzieLet25_4Lcall_main_mask_Bool3_d[0],
                                                                                                                                                sc_0_7_destruct_d[0],
                                                                                                                                                t1acp_1_destruct_d[0],
                                                                                                                                                q1ack_1_destruct_d[0],
                                                                                                                                                t2acq_1_destruct_d[0],
                                                                                                                                                q2acl_1_destruct_d[0]}), lizzieLet25_4Lcall_main_mask_Bool3_d, sc_0_7_destruct_d, t1acp_1_destruct_d, q1ack_1_destruct_d, t2acq_1_destruct_d, q2acl_1_destruct_d);
  assign {lizzieLet25_4Lcall_main_mask_Bool3_r,
          sc_0_7_destruct_r,
          t1acp_1_destruct_r,
          q1ack_1_destruct_r,
          t2acq_1_destruct_r,
          q2acl_1_destruct_r} = {6 {(lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_r && lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2,CTmain_mask_Bool) > (lizzieLet26_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d;
  logic lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_r;
  assign lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_r = ((! lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d[0]) || lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d <= {115'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_r)
        lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d <= lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_d;
  CTmain_mask_Bool_t lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf;
  assign lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_r = (! lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf[0] ? lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf :
                                   lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf <= {115'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf[0]))
        lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf <= {115'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf[0])))
        lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_buf <= lizzieLet25_4Lcall_main_mask_Bool3_1sc_0_7_1t1acp_1_1q1ack_1_1t2acq_1_1q2acl_1_1Lcall_main_mask_Bool2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet25_4Lmain_mask_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                        (lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet25_4Lmain_mask_Boolsbos_emitted;
  logic [1:0] lizzieLet25_4Lmain_mask_Boolsbos_done;
  assign lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d = {lizzieLet25_4Lmain_mask_Boolsbos_d[16:1],
                                                                    (lizzieLet25_4Lmain_mask_Boolsbos_d[0] && (! lizzieLet25_4Lmain_mask_Boolsbos_emitted[0]))};
  assign lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d = {lizzieLet25_4Lmain_mask_Boolsbos_d[16:1],
                                                                    (lizzieLet25_4Lmain_mask_Boolsbos_d[0] && (! lizzieLet25_4Lmain_mask_Boolsbos_emitted[1]))};
  assign lizzieLet25_4Lmain_mask_Boolsbos_done = (lizzieLet25_4Lmain_mask_Boolsbos_emitted | ({lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d[0],
                                                                                               lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r,
                                                                                                                                                              lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet25_4Lmain_mask_Boolsbos_r = (& lizzieLet25_4Lmain_mask_Boolsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lmain_mask_Boolsbos_emitted <= 2'd0;
    else
      lizzieLet25_4Lmain_mask_Boolsbos_emitted <= (lizzieLet25_4Lmain_mask_Boolsbos_r ? 2'd0 :
                                                   lizzieLet25_4Lmain_mask_Boolsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_main_mask_Bool_goConst,Go) */
  assign call_main_mask_Bool_goConst_d = lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r = call_main_mask_Bool_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (main_mask_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r = ((! lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                          1'd0};
    else
      if (lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r)
        lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign main_mask_Bool_resbuf_d = (lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf :
                                    lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                            1'd0};
    else
      if ((main_mask_Bool_resbuf_r && lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                              1'd0};
      else if (((! main_mask_Bool_resbuf_r) && (! lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet25_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool0) : (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) > [(es_2_5_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_3_8_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_4_2_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_14_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted ;
  logic [3:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_done ;
  assign es_2_5_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [19:4],
                              (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [0]))};
  assign es_3_8_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [35:20],
                              (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [1]))};
  assign es_4_2_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [51:36],
                              (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [2]))};
  assign sc_0_14_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [67:52],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [3]))};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_done  = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  | ({sc_0_14_destruct_d[0],
                                                                                                                               es_4_2_destruct_d[0],
                                                                                                                               es_3_8_destruct_d[0],
                                                                                                                               es_2_5_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                                                        es_4_2_destruct_r,
                                                                                                                                                        es_3_8_destruct_r,
                                                                                                                                                        es_2_5_destruct_r}));
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_r  = (& \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  <= 4'd0;
    else
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  <= (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_r  ? 4'd0 :
                                                                   \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool1) : (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) > [(es_3_7_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_4_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_13_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacA_4_destruct,MyDTBool_Bool),
                                                                                                                                     (gacB_4_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'acC_4_destruct,MyBool),
                                                                                                                                     (q1acF_3_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted ;
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_done ;
  assign es_3_7_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [19:4],
                              (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [0]))};
  assign es_4_1_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [35:20],
                              (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [1]))};
  assign sc_0_13_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [51:36],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [2]))};
  assign isZacA_4_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [3]));
  assign gacB_4_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [4]));
  assign \v'acC_4_destruct_d  = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [52:52],
                                 (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [5]))};
  assign q1acF_3_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [68:53],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [6]))};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_done  = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  | ({q1acF_3_destruct_d[0],
                                                                                                                               \v'acC_4_destruct_d [0],
                                                                                                                               gacB_4_destruct_d[0],
                                                                                                                               isZacA_4_destruct_d[0],
                                                                                                                               sc_0_13_destruct_d[0],
                                                                                                                               es_4_1_destruct_d[0],
                                                                                                                               es_3_7_destruct_d[0]} & {q1acF_3_destruct_r,
                                                                                                                                                        \v'acC_4_destruct_r ,
                                                                                                                                                        gacB_4_destruct_r,
                                                                                                                                                        isZacA_4_destruct_r,
                                                                                                                                                        sc_0_13_destruct_r,
                                                                                                                                                        es_4_1_destruct_r,
                                                                                                                                                        es_3_7_destruct_r}));
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_r  = (& \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  <= 7'd0;
    else
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  <= (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_r  ? 7'd0 :
                                                                   \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool2) : (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) > [(es_4_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_12_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacA_3_destruct,MyDTBool_Bool),
                                                                                                                                     (gacB_3_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'acC_3_destruct,MyBool),
                                                                                                                                     (q1acF_2_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2acG_2_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted ;
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_done ;
  assign es_4_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [19:4],
                            (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [0]))};
  assign sc_0_12_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [35:20],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [1]))};
  assign isZacA_3_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [2]));
  assign gacB_3_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [3]));
  assign \v'acC_3_destruct_d  = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [36:36],
                                 (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [4]))};
  assign q1acF_2_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [52:37],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [5]))};
  assign q2acG_2_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [68:53],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [6]))};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_done  = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  | ({q2acG_2_destruct_d[0],
                                                                                                                               q1acF_2_destruct_d[0],
                                                                                                                               \v'acC_3_destruct_d [0],
                                                                                                                               gacB_3_destruct_d[0],
                                                                                                                               isZacA_3_destruct_d[0],
                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                               es_4_destruct_d[0]} & {q2acG_2_destruct_r,
                                                                                                                                                      q1acF_2_destruct_r,
                                                                                                                                                      \v'acC_3_destruct_r ,
                                                                                                                                                      gacB_3_destruct_r,
                                                                                                                                                      isZacA_3_destruct_r,
                                                                                                                                                      sc_0_12_destruct_r,
                                                                                                                                                      es_4_destruct_r}));
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_r  = (& \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  <= 7'd0;
    else
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  <= (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_r  ? 7'd0 :
                                                                   \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool3) : (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) > [(sc_0_11_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacA_2_destruct,MyDTBool_Bool),
                                                                                                                                     (gacB_2_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'acC_2_destruct,MyBool),
                                                                                                                                     (q1acF_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2acG_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q3acH_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted ;
  logic [6:0] \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_done ;
  assign sc_0_11_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [19:4],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [0]))};
  assign isZacA_2_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [1]));
  assign gacB_2_destruct_d = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [2]));
  assign \v'acC_2_destruct_d  = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [20:20],
                                 (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [3]))};
  assign q1acF_1_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [36:21],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [4]))};
  assign q2acG_1_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [52:37],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [5]))};
  assign q3acH_1_destruct_d = {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [68:53],
                               (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [6]))};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_done  = (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  | ({q3acH_1_destruct_d[0],
                                                                                                                               q2acG_1_destruct_d[0],
                                                                                                                               q1acF_1_destruct_d[0],
                                                                                                                               \v'acC_2_destruct_d [0],
                                                                                                                               gacB_2_destruct_d[0],
                                                                                                                               isZacA_2_destruct_d[0],
                                                                                                                               sc_0_11_destruct_d[0]} & {q3acH_1_destruct_r,
                                                                                                                                                         q2acG_1_destruct_r,
                                                                                                                                                         q1acF_1_destruct_r,
                                                                                                                                                         \v'acC_2_destruct_r ,
                                                                                                                                                         gacB_2_destruct_r,
                                                                                                                                                         isZacA_2_destruct_r,
                                                                                                                                                         sc_0_11_destruct_r}));
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_r  = (& \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  <= 7'd0;
    else
      \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  <= (\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_r  ? 7'd0 :
                                                                   \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_done );
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet30_2,CTmap''_map''_Bool_Bool_Bool) (lizzieLet30_1,CTmap''_map''_Bool_Bool_Bool) > [(_22,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool)] */
  logic [4:0] lizzieLet30_1_onehotd;
  always_comb
    if ((lizzieLet30_2_d[0] && lizzieLet30_1_d[0]))
      unique case (lizzieLet30_2_d[3:1])
        3'd0: lizzieLet30_1_onehotd = 5'd1;
        3'd1: lizzieLet30_1_onehotd = 5'd2;
        3'd2: lizzieLet30_1_onehotd = 5'd4;
        3'd3: lizzieLet30_1_onehotd = 5'd8;
        3'd4: lizzieLet30_1_onehotd = 5'd16;
        default: lizzieLet30_1_onehotd = 5'd0;
      endcase
    else lizzieLet30_1_onehotd = 5'd0;
  assign _22_d = {lizzieLet30_1_d[68:1], lizzieLet30_1_onehotd[0]};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_d  = {lizzieLet30_1_d[68:1],
                                                               lizzieLet30_1_onehotd[1]};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_d  = {lizzieLet30_1_d[68:1],
                                                               lizzieLet30_1_onehotd[2]};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_d  = {lizzieLet30_1_d[68:1],
                                                               lizzieLet30_1_onehotd[3]};
  assign \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_d  = {lizzieLet30_1_d[68:1],
                                                               lizzieLet30_1_onehotd[4]};
  assign lizzieLet30_1_r = (| (lizzieLet30_1_onehotd & {\lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                        \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                        \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                        \lizzieLet30_1Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                        _22_r}));
  assign lizzieLet30_2_r = lizzieLet30_1_r;
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty Go) : (lizzieLet30_3,CTmap''_map''_Bool_Bool_Bool) (go_12_goMux_data,Go) > [(_21,Go),
                                                                                      (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3,Go),
                                                                                      (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2,Go),
                                                                                      (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1,Go),
                                                                                      (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0,Go)] */
  logic [4:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet30_3_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet30_3_d[3:1])
        3'd0: go_12_goMux_data_onehotd = 5'd1;
        3'd1: go_12_goMux_data_onehotd = 5'd2;
        3'd2: go_12_goMux_data_onehotd = 5'd4;
        3'd3: go_12_goMux_data_onehotd = 5'd8;
        3'd4: go_12_goMux_data_onehotd = 5'd16;
        default: go_12_goMux_data_onehotd = 5'd0;
      endcase
    else go_12_goMux_data_onehotd = 5'd0;
  assign _21_d = go_12_goMux_data_onehotd[0];
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_d  = go_12_goMux_data_onehotd[1];
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_d  = go_12_goMux_data_onehotd[2];
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_d  = go_12_goMux_data_onehotd[3];
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_d  = go_12_goMux_data_onehotd[4];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                              \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                              \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                              \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                              _21_r}));
  assign lizzieLet30_3_r = go_12_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0,Go) > (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf,Go) */
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_r  = ((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d [0]) || \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_r )
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_d ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r  = (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]);
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d  = (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0] ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  :
                                                                        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r  && \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ) && (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0])))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1,Go) > (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf,Go) */
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_r  = ((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d [0]) || \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_r )
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_d ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r  = (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]);
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d  = (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0] ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  :
                                                                        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r  && \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ) && (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0])))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2,Go) > (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf,Go) */
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_r  = ((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d [0]) || \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_r )
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_d ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r  = (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]);
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d  = (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0] ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  :
                                                                        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r  && \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ) && (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0])))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3,Go) > (lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf,Go) */
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  logic \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_r  = ((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d [0]) || \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_r )
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_d ;
  Go_t \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf ;
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r  = (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]);
  assign \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d  = (\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0] ? \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  :
                                                                        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r  && \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ) && (! \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0])))
        \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= \lizzieLet30_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet30_4,CTmap''_map''_Bool_Bool_Bool) (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet30_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet30_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                             srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                                      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                                      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                                      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                                      \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_r }));
  assign lizzieLet30_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0,Pointer_QTree_Bool),
                          (es_2_5_destruct,Pointer_QTree_Bool),
                          (es_3_8_destruct,Pointer_QTree_Bool),
                          (es_4_2_destruct,Pointer_QTree_Bool)] > (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_d [0],
                                                                                                                    es_2_5_destruct_d[0],
                                                                                                                    es_3_8_destruct_d[0],
                                                                                                                    es_4_2_destruct_d[0]}), \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_d , es_2_5_destruct_d, es_3_8_destruct_d, es_4_2_destruct_d);
  assign {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_r ,
          es_2_5_destruct_r,
          es_3_8_destruct_r,
          es_4_2_destruct_r} = {4 {(\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_r  && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool,QTree_Bool) > (lizzieLet34_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_r ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_r  = ((! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d [0]) || \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                                         1'd0};
    else
      if (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_r )
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_r  = (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet34_1_argbuf_d = (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf [0] ? \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                           1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                             1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_buf  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_5_1es_3_8_1es_4_2_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool0) : [(lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                 (es_3_7_destruct,Pointer_QTree_Bool),
                                                 (es_4_1_destruct,Pointer_QTree_Bool),
                                                 (sc_0_13_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d  = \Lcall_map''_map''_Bool_Bool_Bool0_dc ((& {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_d [0],
                                                                                                                                                                     es_3_7_destruct_d[0],
                                                                                                                                                                     es_4_1_destruct_d[0],
                                                                                                                                                                     sc_0_13_destruct_d[0]}), \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_d , es_3_7_destruct_d, es_4_1_destruct_d, sc_0_13_destruct_d);
  assign {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_r ,
          es_3_7_destruct_r,
          es_4_1_destruct_r,
          sc_0_13_destruct_r} = {4 {(\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r  && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet33_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r  = ((! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d [0]) || \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= {68'd0,
                                                                                                                                 1'd0};
    else
      if (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r )
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r  = (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]);
  assign lizzieLet33_1_argbuf_d = (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0] ? \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  :
                                   \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= {68'd0,
                                                                                                                                   1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= {68'd0,
                                                                                                                                     1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0])))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_7_1es_4_1_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool1) : [(lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                 (es_4_destruct,Pointer_QTree_Bool),
                                                 (sc_0_12_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (isZacA_3_1,MyDTBool_Bool),
                                                 (gacB_3_1,MyDTBool_Bool_Bool),
                                                 (v'acC_3_1,MyBool),
                                                 (q1acF_2_destruct,Pointer_QTree_Bool)] > (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_d  = \Lcall_map''_map''_Bool_Bool_Bool1_dc ((& {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_d [0],
                                                                                                                                                                                               es_4_destruct_d[0],
                                                                                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                                                                                               isZacA_3_1_d[0],
                                                                                                                                                                                               gacB_3_1_d[0],
                                                                                                                                                                                               \v'acC_3_1_d [0],
                                                                                                                                                                                               q1acF_2_destruct_d[0]}), \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_d , es_4_destruct_d, sc_0_12_destruct_d, isZacA_3_1_d, gacB_3_1_d, \v'acC_3_1_d , q1acF_2_destruct_d);
  assign {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_r ,
          es_4_destruct_r,
          sc_0_12_destruct_r,
          isZacA_3_1_r,
          gacB_3_1_r,
          \v'acC_3_1_r ,
          q1acF_2_destruct_r} = {7 {(\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_r  && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet32_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_r  = ((! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d [0]) || \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= {68'd0,
                                                                                                                                                           1'd0};
    else
      if (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_r )
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r  = (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]);
  assign lizzieLet32_1_argbuf_d = (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0] ? \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  :
                                   \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= {68'd0,
                                                                                                                                                             1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= {68'd0,
                                                                                                                                                               1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0])))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_1sc_0_12_1isZacA_3_1gacB_3_1v'acC_3_1q1acF_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool2) : [(lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                 (sc_0_11_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (isZacA_2_1,MyDTBool_Bool),
                                                 (gacB_2_1,MyDTBool_Bool_Bool),
                                                 (v'acC_2_1,MyBool),
                                                 (q1acF_1_destruct,Pointer_QTree_Bool),
                                                 (q2acG_1_destruct,Pointer_QTree_Bool)] > (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_d  = \Lcall_map''_map''_Bool_Bool_Bool2_dc ((& {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_d [0],
                                                                                                                                                                                                  sc_0_11_destruct_d[0],
                                                                                                                                                                                                  isZacA_2_1_d[0],
                                                                                                                                                                                                  gacB_2_1_d[0],
                                                                                                                                                                                                  \v'acC_2_1_d [0],
                                                                                                                                                                                                  q1acF_1_destruct_d[0],
                                                                                                                                                                                                  q2acG_1_destruct_d[0]}), \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_d , sc_0_11_destruct_d, isZacA_2_1_d, gacB_2_1_d, \v'acC_2_1_d , q1acF_1_destruct_d, q2acG_1_destruct_d);
  assign {\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_r ,
          sc_0_11_destruct_r,
          isZacA_2_1_r,
          gacB_2_1_r,
          \v'acC_2_1_r ,
          q1acF_1_destruct_r,
          q2acG_1_destruct_r} = {7 {(\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_r  && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet31_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  logic \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_r  = ((! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d [0]) || \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= {68'd0,
                                                                                                                                                              1'd0};
    else
      if (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_r )
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf ;
  assign \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r  = (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]);
  assign lizzieLet31_1_argbuf_d = (\lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0] ? \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  :
                                   \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= {68'd0,
                                                                                                                                                                1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= {68'd0,
                                                                                                                                                                  1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0])))
        \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= \lizzieLet30_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacA_2_1gacB_2_1v'acC_2_1q1acF_1_1q2acG_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                                    (lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted ;
  logic [1:0] \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_done ;
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d  = {\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d [16:1],
                                                                                  (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d [0] && (! \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted [0]))};
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d  = {\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d [16:1],
                                                                                  (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_d [0] && (! \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted [1]))};
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_done  = (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  | ({\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d [0],
                                                                                                                           \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                        \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_r  = (& \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  <= 2'd0;
    else
      \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  <= (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_r  ? 2'd0 :
                                                                 \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_map''_map''_Bool_Bool_Bool_goConst,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_goConst_d  = \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r  = \call_map''_map''_Bool_Bool_Bool_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (map''_map''_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                        1'd0};
    else
      if (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r )
        \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Bool_t \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \map''_map''_Bool_Bool_Bool_resbuf_d  = (\lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  :
                                                  \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                          1'd0};
    else
      if ((\map''_map''_Bool_Bool_Bool_resbuf_r  && \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                            1'd0};
      else if (((! \map''_map''_Bool_Bool_Bool_resbuf_r ) && (! \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet30_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet4_1MQNode,MaskQTree) > [(q1ack_destruct,Pointer_MaskQTree),
                                                           (q2acl_destruct,Pointer_MaskQTree),
                                                           (q3acm_destruct,Pointer_MaskQTree),
                                                           (q4acn_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet4_1MQNode_emitted;
  logic [3:0] lizzieLet4_1MQNode_done;
  assign q1ack_destruct_d = {lizzieLet4_1MQNode_d[18:3],
                             (lizzieLet4_1MQNode_d[0] && (! lizzieLet4_1MQNode_emitted[0]))};
  assign q2acl_destruct_d = {lizzieLet4_1MQNode_d[34:19],
                             (lizzieLet4_1MQNode_d[0] && (! lizzieLet4_1MQNode_emitted[1]))};
  assign q3acm_destruct_d = {lizzieLet4_1MQNode_d[50:35],
                             (lizzieLet4_1MQNode_d[0] && (! lizzieLet4_1MQNode_emitted[2]))};
  assign q4acn_destruct_d = {lizzieLet4_1MQNode_d[66:51],
                             (lizzieLet4_1MQNode_d[0] && (! lizzieLet4_1MQNode_emitted[3]))};
  assign lizzieLet4_1MQNode_done = (lizzieLet4_1MQNode_emitted | ({q4acn_destruct_d[0],
                                                                   q3acm_destruct_d[0],
                                                                   q2acl_destruct_d[0],
                                                                   q1ack_destruct_d[0]} & {q4acn_destruct_r,
                                                                                           q3acm_destruct_r,
                                                                                           q2acl_destruct_r,
                                                                                           q1ack_destruct_r}));
  assign lizzieLet4_1MQNode_r = (& lizzieLet4_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1MQNode_emitted <= 4'd0;
    else
      lizzieLet4_1MQNode_emitted <= (lizzieLet4_1MQNode_r ? 4'd0 :
                                     lizzieLet4_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet4_2,MaskQTree) (lizzieLet4_1,MaskQTree) > [(_20,MaskQTree),
                                                                            (_19,MaskQTree),
                                                                            (lizzieLet4_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 3'd1;
        2'd1: lizzieLet4_1_onehotd = 3'd2;
        2'd2: lizzieLet4_1_onehotd = 3'd4;
        default: lizzieLet4_1_onehotd = 3'd0;
      endcase
    else lizzieLet4_1_onehotd = 3'd0;
  assign _20_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _19_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1MQNode_d = {lizzieLet4_1_d[66:1],
                                 lizzieLet4_1_onehotd[2]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {lizzieLet4_1MQNode_r,
                                                      _19_r,
                                                      _20_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet4_3,MaskQTree) (go_5_goMux_data,Go) > [(lizzieLet4_3MQNone,Go),
                                                                 (lizzieLet4_3MQVal,Go),
                                                                 (lizzieLet4_3MQNode,Go)] */
  logic [2:0] go_5_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_5_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_5_goMux_data_onehotd = 3'd1;
        2'd1: go_5_goMux_data_onehotd = 3'd2;
        2'd2: go_5_goMux_data_onehotd = 3'd4;
        default: go_5_goMux_data_onehotd = 3'd0;
      endcase
    else go_5_goMux_data_onehotd = 3'd0;
  assign lizzieLet4_3MQNone_d = go_5_goMux_data_onehotd[0];
  assign lizzieLet4_3MQVal_d = go_5_goMux_data_onehotd[1];
  assign lizzieLet4_3MQNode_d = go_5_goMux_data_onehotd[2];
  assign go_5_goMux_data_r = (| (go_5_goMux_data_onehotd & {lizzieLet4_3MQNode_r,
                                                            lizzieLet4_3MQVal_r,
                                                            lizzieLet4_3MQNone_r}));
  assign lizzieLet4_3_r = go_5_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3MQNone,Go) > [(lizzieLet4_3MQNone_1,Go),
                                          (lizzieLet4_3MQNone_2,Go)] */
  logic [1:0] lizzieLet4_3MQNone_emitted;
  logic [1:0] lizzieLet4_3MQNone_done;
  assign lizzieLet4_3MQNone_1_d = (lizzieLet4_3MQNone_d[0] && (! lizzieLet4_3MQNone_emitted[0]));
  assign lizzieLet4_3MQNone_2_d = (lizzieLet4_3MQNone_d[0] && (! lizzieLet4_3MQNone_emitted[1]));
  assign lizzieLet4_3MQNone_done = (lizzieLet4_3MQNone_emitted | ({lizzieLet4_3MQNone_2_d[0],
                                                                   lizzieLet4_3MQNone_1_d[0]} & {lizzieLet4_3MQNone_2_r,
                                                                                                 lizzieLet4_3MQNone_1_r}));
  assign lizzieLet4_3MQNone_r = (& lizzieLet4_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQNone_emitted <= 2'd0;
    else
      lizzieLet4_3MQNone_emitted <= (lizzieLet4_3MQNone_r ? 2'd0 :
                                     lizzieLet4_3MQNone_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet4_3MQNone_1,Go)] > (lizzieLet4_3MQNone_1QNone_Bool,QTree_Bool) */
  assign lizzieLet4_3MQNone_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet4_3MQNone_1_d[0]}), lizzieLet4_3MQNone_1_d);
  assign {lizzieLet4_3MQNone_1_r} = {1 {(lizzieLet4_3MQNone_1QNone_Bool_r && lizzieLet4_3MQNone_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet4_3MQNone_1QNone_Bool,QTree_Bool) > (lizzieLet5_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet4_3MQNone_1QNone_Bool_bufchan_d;
  logic lizzieLet4_3MQNone_1QNone_Bool_bufchan_r;
  assign lizzieLet4_3MQNone_1QNone_Bool_r = ((! lizzieLet4_3MQNone_1QNone_Bool_bufchan_d[0]) || lizzieLet4_3MQNone_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3MQNone_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet4_3MQNone_1QNone_Bool_r)
        lizzieLet4_3MQNone_1QNone_Bool_bufchan_d <= lizzieLet4_3MQNone_1QNone_Bool_d;
  QTree_Bool_t lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf;
  assign lizzieLet4_3MQNone_1QNone_Bool_bufchan_r = (! lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf[0] ? lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf :
                                  lizzieLet4_3MQNone_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf[0]))
        lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf[0])))
        lizzieLet4_3MQNone_1QNone_Bool_bufchan_buf <= lizzieLet4_3MQNone_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3MQNone_2,Go) > (lizzieLet4_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet4_3MQNone_2_bufchan_d;
  logic lizzieLet4_3MQNone_2_bufchan_r;
  assign lizzieLet4_3MQNone_2_r = ((! lizzieLet4_3MQNone_2_bufchan_d[0]) || lizzieLet4_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3MQNone_2_r)
        lizzieLet4_3MQNone_2_bufchan_d <= lizzieLet4_3MQNone_2_d;
  Go_t lizzieLet4_3MQNone_2_bufchan_buf;
  assign lizzieLet4_3MQNone_2_bufchan_r = (! lizzieLet4_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet4_3MQNone_2_argbuf_d = (lizzieLet4_3MQNone_2_bufchan_buf[0] ? lizzieLet4_3MQNone_2_bufchan_buf :
                                          lizzieLet4_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3MQNone_2_argbuf_r && lizzieLet4_3MQNone_2_bufchan_buf[0]))
        lizzieLet4_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3MQNone_2_argbuf_r) && (! lizzieLet4_3MQNone_2_bufchan_buf[0])))
        lizzieLet4_3MQNone_2_bufchan_buf <= lizzieLet4_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet4_3MQNone_2_argbuf,Go),
                           (lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf,Go),
                           (lizzieLet4_3MQVal_1_argbuf,Go),
                           (lizzieLet4_4MQNode_3QNone_Bool_2_argbuf,Go),
                           (lizzieLet4_4MQNode_3QVal_Bool_2_argbuf,Go),
                           (lizzieLet4_4MQNode_3QError_Bool_2_argbuf,Go)] > (go_11_goMux_choice,C6) (go_11_goMux_data,Go) */
  logic [5:0] lizzieLet4_3MQNone_2_argbuf_select_d;
  assign lizzieLet4_3MQNone_2_argbuf_select_d = ((| lizzieLet4_3MQNone_2_argbuf_select_q) ? lizzieLet4_3MQNone_2_argbuf_select_q :
                                                 (lizzieLet4_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                  (lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_d[0] ? 6'd2 :
                                                   (lizzieLet4_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                    (lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_d[0] ? 6'd8 :
                                                     (lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_d[0] ? 6'd16 :
                                                      (lizzieLet4_4MQNode_3QError_Bool_2_argbuf_d[0] ? 6'd32 :
                                                       6'd0)))))));
  logic [5:0] lizzieLet4_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet4_3MQNone_2_argbuf_select_q <= (lizzieLet4_3MQNone_2_argbuf_done ? 6'd0 :
                                               lizzieLet4_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3MQNone_2_argbuf_emit_q <= (lizzieLet4_3MQNone_2_argbuf_done ? 2'd0 :
                                             lizzieLet4_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3MQNone_2_argbuf_emit_d;
  assign lizzieLet4_3MQNone_2_argbuf_emit_d = (lizzieLet4_3MQNone_2_argbuf_emit_q | ({go_11_goMux_choice_d[0],
                                                                                      go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                go_11_goMux_data_r}));
  logic lizzieLet4_3MQNone_2_argbuf_done;
  assign lizzieLet4_3MQNone_2_argbuf_done = (& lizzieLet4_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet4_4MQNode_3QError_Bool_2_argbuf_r,
          lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_r,
          lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_r,
          lizzieLet4_3MQVal_1_argbuf_r,
          lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_r,
          lizzieLet4_3MQNone_2_argbuf_r} = (lizzieLet4_3MQNone_2_argbuf_done ? lizzieLet4_3MQNone_2_argbuf_select_d :
                                            6'd0);
  assign go_11_goMux_data_d = ((lizzieLet4_3MQNone_2_argbuf_select_d[0] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet4_3MQNone_2_argbuf_d :
                               ((lizzieLet4_3MQNone_2_argbuf_select_d[1] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet25_3Lcall_main_mask_Bool0_1_argbuf_d :
                                ((lizzieLet4_3MQNone_2_argbuf_select_d[2] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet4_3MQVal_1_argbuf_d :
                                 ((lizzieLet4_3MQNone_2_argbuf_select_d[3] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_d :
                                  ((lizzieLet4_3MQNone_2_argbuf_select_d[4] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_d :
                                   ((lizzieLet4_3MQNone_2_argbuf_select_d[5] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet4_4MQNode_3QError_Bool_2_argbuf_d :
                                    1'd0))))));
  assign go_11_goMux_choice_d = ((lizzieLet4_3MQNone_2_argbuf_select_d[0] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet4_3MQNone_2_argbuf_select_d[1] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet4_3MQNone_2_argbuf_select_d[2] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet4_3MQNone_2_argbuf_select_d[3] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet4_3MQNone_2_argbuf_select_d[4] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet4_3MQNone_2_argbuf_select_d[5] && (! lizzieLet4_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet4_3MQVal,Go) > (lizzieLet4_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet4_3MQVal_bufchan_d;
  logic lizzieLet4_3MQVal_bufchan_r;
  assign lizzieLet4_3MQVal_r = ((! lizzieLet4_3MQVal_bufchan_d[0]) || lizzieLet4_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3MQVal_r)
        lizzieLet4_3MQVal_bufchan_d <= lizzieLet4_3MQVal_d;
  Go_t lizzieLet4_3MQVal_bufchan_buf;
  assign lizzieLet4_3MQVal_bufchan_r = (! lizzieLet4_3MQVal_bufchan_buf[0]);
  assign lizzieLet4_3MQVal_1_argbuf_d = (lizzieLet4_3MQVal_bufchan_buf[0] ? lizzieLet4_3MQVal_bufchan_buf :
                                         lizzieLet4_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3MQVal_1_argbuf_r && lizzieLet4_3MQVal_bufchan_buf[0]))
        lizzieLet4_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3MQVal_1_argbuf_r) && (! lizzieLet4_3MQVal_bufchan_buf[0])))
        lizzieLet4_3MQVal_bufchan_buf <= lizzieLet4_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Bool) : (lizzieLet4_4,MaskQTree) (readPointer_QTree_Boolmaci_1_argbuf_rwb,QTree_Bool) > [(_18,QTree_Bool),
                                                                                                         (_17,QTree_Bool),
                                                                                                         (lizzieLet4_4MQNode,QTree_Bool)] */
  logic [2:0] readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && readPointer_QTree_Boolmaci_1_argbuf_rwb_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd = 3'd0;
  assign _18_d = {readPointer_QTree_Boolmaci_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd[0]};
  assign _17_d = {readPointer_QTree_Boolmaci_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet4_4MQNode_d = {readPointer_QTree_Boolmaci_1_argbuf_rwb_d[66:1],
                                 readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Boolmaci_1_argbuf_rwb_r = (| (readPointer_QTree_Boolmaci_1_argbuf_rwb_onehotd & {lizzieLet4_4MQNode_r,
                                                                                                            _17_r,
                                                                                                            _18_r}));
  assign lizzieLet4_4_r = readPointer_QTree_Boolmaci_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet4_4MQNode,QTree_Bool) > [(lizzieLet4_4MQNode_1,QTree_Bool),
                                                          (lizzieLet4_4MQNode_2,QTree_Bool),
                                                          (lizzieLet4_4MQNode_3,QTree_Bool),
                                                          (lizzieLet4_4MQNode_4,QTree_Bool),
                                                          (lizzieLet4_4MQNode_5,QTree_Bool),
                                                          (lizzieLet4_4MQNode_6,QTree_Bool),
                                                          (lizzieLet4_4MQNode_7,QTree_Bool),
                                                          (lizzieLet4_4MQNode_8,QTree_Bool)] */
  logic [7:0] lizzieLet4_4MQNode_emitted;
  logic [7:0] lizzieLet4_4MQNode_done;
  assign lizzieLet4_4MQNode_1_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[0]))};
  assign lizzieLet4_4MQNode_2_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[1]))};
  assign lizzieLet4_4MQNode_3_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[2]))};
  assign lizzieLet4_4MQNode_4_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[3]))};
  assign lizzieLet4_4MQNode_5_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[4]))};
  assign lizzieLet4_4MQNode_6_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[5]))};
  assign lizzieLet4_4MQNode_7_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[6]))};
  assign lizzieLet4_4MQNode_8_d = {lizzieLet4_4MQNode_d[66:1],
                                   (lizzieLet4_4MQNode_d[0] && (! lizzieLet4_4MQNode_emitted[7]))};
  assign lizzieLet4_4MQNode_done = (lizzieLet4_4MQNode_emitted | ({lizzieLet4_4MQNode_8_d[0],
                                                                   lizzieLet4_4MQNode_7_d[0],
                                                                   lizzieLet4_4MQNode_6_d[0],
                                                                   lizzieLet4_4MQNode_5_d[0],
                                                                   lizzieLet4_4MQNode_4_d[0],
                                                                   lizzieLet4_4MQNode_3_d[0],
                                                                   lizzieLet4_4MQNode_2_d[0],
                                                                   lizzieLet4_4MQNode_1_d[0]} & {lizzieLet4_4MQNode_8_r,
                                                                                                 lizzieLet4_4MQNode_7_r,
                                                                                                 lizzieLet4_4MQNode_6_r,
                                                                                                 lizzieLet4_4MQNode_5_r,
                                                                                                 lizzieLet4_4MQNode_4_r,
                                                                                                 lizzieLet4_4MQNode_3_r,
                                                                                                 lizzieLet4_4MQNode_2_r,
                                                                                                 lizzieLet4_4MQNode_1_r}));
  assign lizzieLet4_4MQNode_r = (& lizzieLet4_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_4MQNode_emitted <= 8'd0;
    else
      lizzieLet4_4MQNode_emitted <= (lizzieLet4_4MQNode_r ? 8'd0 :
                                     lizzieLet4_4MQNode_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet4_4MQNode_1QNode_Bool,QTree_Bool) > [(t1acp_destruct,Pointer_QTree_Bool),
                                                                            (t2acq_destruct,Pointer_QTree_Bool),
                                                                            (t3acr_destruct,Pointer_QTree_Bool),
                                                                            (t4acs_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet4_4MQNode_1QNode_Bool_emitted;
  logic [3:0] lizzieLet4_4MQNode_1QNode_Bool_done;
  assign t1acp_destruct_d = {lizzieLet4_4MQNode_1QNode_Bool_d[18:3],
                             (lizzieLet4_4MQNode_1QNode_Bool_d[0] && (! lizzieLet4_4MQNode_1QNode_Bool_emitted[0]))};
  assign t2acq_destruct_d = {lizzieLet4_4MQNode_1QNode_Bool_d[34:19],
                             (lizzieLet4_4MQNode_1QNode_Bool_d[0] && (! lizzieLet4_4MQNode_1QNode_Bool_emitted[1]))};
  assign t3acr_destruct_d = {lizzieLet4_4MQNode_1QNode_Bool_d[50:35],
                             (lizzieLet4_4MQNode_1QNode_Bool_d[0] && (! lizzieLet4_4MQNode_1QNode_Bool_emitted[2]))};
  assign t4acs_destruct_d = {lizzieLet4_4MQNode_1QNode_Bool_d[66:51],
                             (lizzieLet4_4MQNode_1QNode_Bool_d[0] && (! lizzieLet4_4MQNode_1QNode_Bool_emitted[3]))};
  assign lizzieLet4_4MQNode_1QNode_Bool_done = (lizzieLet4_4MQNode_1QNode_Bool_emitted | ({t4acs_destruct_d[0],
                                                                                           t3acr_destruct_d[0],
                                                                                           t2acq_destruct_d[0],
                                                                                           t1acp_destruct_d[0]} & {t4acs_destruct_r,
                                                                                                                   t3acr_destruct_r,
                                                                                                                   t2acq_destruct_r,
                                                                                                                   t1acp_destruct_r}));
  assign lizzieLet4_4MQNode_1QNode_Bool_r = (& lizzieLet4_4MQNode_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet4_4MQNode_1QNode_Bool_emitted <= (lizzieLet4_4MQNode_1QNode_Bool_r ? 4'd0 :
                                                 lizzieLet4_4MQNode_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet4_4MQNode_2,QTree_Bool) (lizzieLet4_4MQNode_1,QTree_Bool) > [(_16,QTree_Bool),
                                                                                               (_15,QTree_Bool),
                                                                                               (lizzieLet4_4MQNode_1QNode_Bool,QTree_Bool),
                                                                                               (_14,QTree_Bool)] */
  logic [3:0] lizzieLet4_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_2_d[0] && lizzieLet4_4MQNode_1_d[0]))
      unique case (lizzieLet4_4MQNode_2_d[2:1])
        2'd0: lizzieLet4_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet4_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet4_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet4_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet4_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_4MQNode_1_onehotd = 4'd0;
  assign _16_d = {lizzieLet4_4MQNode_1_d[66:1],
                  lizzieLet4_4MQNode_1_onehotd[0]};
  assign _15_d = {lizzieLet4_4MQNode_1_d[66:1],
                  lizzieLet4_4MQNode_1_onehotd[1]};
  assign lizzieLet4_4MQNode_1QNode_Bool_d = {lizzieLet4_4MQNode_1_d[66:1],
                                             lizzieLet4_4MQNode_1_onehotd[2]};
  assign _14_d = {lizzieLet4_4MQNode_1_d[66:1],
                  lizzieLet4_4MQNode_1_onehotd[3]};
  assign lizzieLet4_4MQNode_1_r = (| (lizzieLet4_4MQNode_1_onehotd & {_14_r,
                                                                      lizzieLet4_4MQNode_1QNode_Bool_r,
                                                                      _15_r,
                                                                      _16_r}));
  assign lizzieLet4_4MQNode_2_r = lizzieLet4_4MQNode_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet4_4MQNode_3,QTree_Bool) (lizzieLet4_3MQNode,Go) > [(lizzieLet4_4MQNode_3QNone_Bool,Go),
                                                                             (lizzieLet4_4MQNode_3QVal_Bool,Go),
                                                                             (lizzieLet4_4MQNode_3QNode_Bool,Go),
                                                                             (lizzieLet4_4MQNode_3QError_Bool,Go)] */
  logic [3:0] lizzieLet4_3MQNode_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_3_d[0] && lizzieLet4_3MQNode_d[0]))
      unique case (lizzieLet4_4MQNode_3_d[2:1])
        2'd0: lizzieLet4_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet4_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet4_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet4_3MQNode_onehotd = 4'd8;
        default: lizzieLet4_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet4_3MQNode_onehotd = 4'd0;
  assign lizzieLet4_4MQNode_3QNone_Bool_d = lizzieLet4_3MQNode_onehotd[0];
  assign lizzieLet4_4MQNode_3QVal_Bool_d = lizzieLet4_3MQNode_onehotd[1];
  assign lizzieLet4_4MQNode_3QNode_Bool_d = lizzieLet4_3MQNode_onehotd[2];
  assign lizzieLet4_4MQNode_3QError_Bool_d = lizzieLet4_3MQNode_onehotd[3];
  assign lizzieLet4_3MQNode_r = (| (lizzieLet4_3MQNode_onehotd & {lizzieLet4_4MQNode_3QError_Bool_r,
                                                                  lizzieLet4_4MQNode_3QNode_Bool_r,
                                                                  lizzieLet4_4MQNode_3QVal_Bool_r,
                                                                  lizzieLet4_4MQNode_3QNone_Bool_r}));
  assign lizzieLet4_4MQNode_3_r = lizzieLet4_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet4_4MQNode_3QError_Bool,Go) > [(lizzieLet4_4MQNode_3QError_Bool_1,Go),
                                                       (lizzieLet4_4MQNode_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet4_4MQNode_3QError_Bool_emitted;
  logic [1:0] lizzieLet4_4MQNode_3QError_Bool_done;
  assign lizzieLet4_4MQNode_3QError_Bool_1_d = (lizzieLet4_4MQNode_3QError_Bool_d[0] && (! lizzieLet4_4MQNode_3QError_Bool_emitted[0]));
  assign lizzieLet4_4MQNode_3QError_Bool_2_d = (lizzieLet4_4MQNode_3QError_Bool_d[0] && (! lizzieLet4_4MQNode_3QError_Bool_emitted[1]));
  assign lizzieLet4_4MQNode_3QError_Bool_done = (lizzieLet4_4MQNode_3QError_Bool_emitted | ({lizzieLet4_4MQNode_3QError_Bool_2_d[0],
                                                                                             lizzieLet4_4MQNode_3QError_Bool_1_d[0]} & {lizzieLet4_4MQNode_3QError_Bool_2_r,
                                                                                                                                        lizzieLet4_4MQNode_3QError_Bool_1_r}));
  assign lizzieLet4_4MQNode_3QError_Bool_r = (& lizzieLet4_4MQNode_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet4_4MQNode_3QError_Bool_emitted <= (lizzieLet4_4MQNode_3QError_Bool_r ? 2'd0 :
                                                  lizzieLet4_4MQNode_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet4_4MQNode_3QError_Bool_1,Go)] > (lizzieLet4_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet4_4MQNode_3QError_Bool_1_d[0]}), lizzieLet4_4MQNode_3QError_Bool_1_d);
  assign {lizzieLet4_4MQNode_3QError_Bool_1_r} = {1 {(lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_r && lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet4_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet10_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_r = ((! lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_r)
        lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet4_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_4MQNode_3QError_Bool_2,Go) > (lizzieLet4_4MQNode_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d;
  logic lizzieLet4_4MQNode_3QError_Bool_2_bufchan_r;
  assign lizzieLet4_4MQNode_3QError_Bool_2_r = ((! lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d[0]) || lizzieLet4_4MQNode_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_4MQNode_3QError_Bool_2_r)
        lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d <= lizzieLet4_4MQNode_3QError_Bool_2_d;
  Go_t lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf;
  assign lizzieLet4_4MQNode_3QError_Bool_2_bufchan_r = (! lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_3QError_Bool_2_argbuf_d = (lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf[0] ? lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf :
                                                       lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_4MQNode_3QError_Bool_2_argbuf_r && lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_4MQNode_3QError_Bool_2_argbuf_r) && (! lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QError_Bool_2_bufchan_buf <= lizzieLet4_4MQNode_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_4MQNode_3QNode_Bool,Go) > (lizzieLet4_4MQNode_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet4_4MQNode_3QNode_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_3QNode_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_3QNode_Bool_r = ((! lizzieLet4_4MQNode_3QNode_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_4MQNode_3QNode_Bool_r)
        lizzieLet4_4MQNode_3QNode_Bool_bufchan_d <= lizzieLet4_4MQNode_3QNode_Bool_d;
  Go_t lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_3QNode_Bool_bufchan_r = (! lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_d = (lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf :
                                                      lizzieLet4_4MQNode_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_r && lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_4MQNode_3QNode_Bool_1_argbuf_r) && (! lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QNode_Bool_bufchan_buf <= lizzieLet4_4MQNode_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_4MQNode_3QNone_Bool,Go) > [(lizzieLet4_4MQNode_3QNone_Bool_1,Go),
                                                      (lizzieLet4_4MQNode_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet4_4MQNode_3QNone_Bool_emitted;
  logic [1:0] lizzieLet4_4MQNode_3QNone_Bool_done;
  assign lizzieLet4_4MQNode_3QNone_Bool_1_d = (lizzieLet4_4MQNode_3QNone_Bool_d[0] && (! lizzieLet4_4MQNode_3QNone_Bool_emitted[0]));
  assign lizzieLet4_4MQNode_3QNone_Bool_2_d = (lizzieLet4_4MQNode_3QNone_Bool_d[0] && (! lizzieLet4_4MQNode_3QNone_Bool_emitted[1]));
  assign lizzieLet4_4MQNode_3QNone_Bool_done = (lizzieLet4_4MQNode_3QNone_Bool_emitted | ({lizzieLet4_4MQNode_3QNone_Bool_2_d[0],
                                                                                           lizzieLet4_4MQNode_3QNone_Bool_1_d[0]} & {lizzieLet4_4MQNode_3QNone_Bool_2_r,
                                                                                                                                     lizzieLet4_4MQNode_3QNone_Bool_1_r}));
  assign lizzieLet4_4MQNode_3QNone_Bool_r = (& lizzieLet4_4MQNode_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet4_4MQNode_3QNone_Bool_emitted <= (lizzieLet4_4MQNode_3QNone_Bool_r ? 2'd0 :
                                                 lizzieLet4_4MQNode_3QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet4_4MQNode_3QNone_Bool_1,Go)] > (lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet4_4MQNode_3QNone_Bool_1_d[0]}), lizzieLet4_4MQNode_3QNone_Bool_1_d);
  assign {lizzieLet4_4MQNode_3QNone_Bool_1_r} = {1 {(lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_r && lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet7_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_r = ((! lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0,
                                                               1'd0};
    else
      if (lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_r)
        lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf :
                                  lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                   1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet4_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_4MQNode_3QNone_Bool_2,Go) > (lizzieLet4_4MQNode_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d;
  logic lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_r;
  assign lizzieLet4_4MQNode_3QNone_Bool_2_r = ((! lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d[0]) || lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_4MQNode_3QNone_Bool_2_r)
        lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d <= lizzieLet4_4MQNode_3QNone_Bool_2_d;
  Go_t lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_r = (! lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_d = (lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf :
                                                      lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_r && lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_4MQNode_3QNone_Bool_2_argbuf_r) && (! lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_buf <= lizzieLet4_4MQNode_3QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_4MQNode_3QVal_Bool,Go) > [(lizzieLet4_4MQNode_3QVal_Bool_1,Go),
                                                     (lizzieLet4_4MQNode_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet4_4MQNode_3QVal_Bool_emitted;
  logic [1:0] lizzieLet4_4MQNode_3QVal_Bool_done;
  assign lizzieLet4_4MQNode_3QVal_Bool_1_d = (lizzieLet4_4MQNode_3QVal_Bool_d[0] && (! lizzieLet4_4MQNode_3QVal_Bool_emitted[0]));
  assign lizzieLet4_4MQNode_3QVal_Bool_2_d = (lizzieLet4_4MQNode_3QVal_Bool_d[0] && (! lizzieLet4_4MQNode_3QVal_Bool_emitted[1]));
  assign lizzieLet4_4MQNode_3QVal_Bool_done = (lizzieLet4_4MQNode_3QVal_Bool_emitted | ({lizzieLet4_4MQNode_3QVal_Bool_2_d[0],
                                                                                         lizzieLet4_4MQNode_3QVal_Bool_1_d[0]} & {lizzieLet4_4MQNode_3QVal_Bool_2_r,
                                                                                                                                  lizzieLet4_4MQNode_3QVal_Bool_1_r}));
  assign lizzieLet4_4MQNode_3QVal_Bool_r = (& lizzieLet4_4MQNode_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_4MQNode_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet4_4MQNode_3QVal_Bool_emitted <= (lizzieLet4_4MQNode_3QVal_Bool_r ? 2'd0 :
                                                lizzieLet4_4MQNode_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet4_4MQNode_3QVal_Bool_1,Go)] > (lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet4_4MQNode_3QVal_Bool_1_d[0]}), lizzieLet4_4MQNode_3QVal_Bool_1_d);
  assign {lizzieLet4_4MQNode_3QVal_Bool_1_r} = {1 {(lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_r && lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet8_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_r = ((! lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                               1'd0};
    else
      if (lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_r)
        lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                   1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet4_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_4MQNode_3QVal_Bool_2,Go) > (lizzieLet4_4MQNode_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d;
  logic lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_r;
  assign lizzieLet4_4MQNode_3QVal_Bool_2_r = ((! lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d[0]) || lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_4MQNode_3QVal_Bool_2_r)
        lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d <= lizzieLet4_4MQNode_3QVal_Bool_2_d;
  Go_t lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_r = (! lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_d = (lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf :
                                                     lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_r && lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_4MQNode_3QVal_Bool_2_argbuf_r) && (! lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_buf <= lizzieLet4_4MQNode_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_4MQNode_4,QTree_Bool) (lizzieLet4_6MQNode,Pointer_CTmain_mask_Bool) > [(lizzieLet4_4MQNode_4QNone_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                         (lizzieLet4_4MQNode_4QVal_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                         (lizzieLet4_4MQNode_4QNode_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                         (lizzieLet4_4MQNode_4QError_Bool,Pointer_CTmain_mask_Bool)] */
  logic [3:0] lizzieLet4_6MQNode_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_4_d[0] && lizzieLet4_6MQNode_d[0]))
      unique case (lizzieLet4_4MQNode_4_d[2:1])
        2'd0: lizzieLet4_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet4_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet4_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet4_6MQNode_onehotd = 4'd8;
        default: lizzieLet4_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet4_6MQNode_onehotd = 4'd0;
  assign lizzieLet4_4MQNode_4QNone_Bool_d = {lizzieLet4_6MQNode_d[16:1],
                                             lizzieLet4_6MQNode_onehotd[0]};
  assign lizzieLet4_4MQNode_4QVal_Bool_d = {lizzieLet4_6MQNode_d[16:1],
                                            lizzieLet4_6MQNode_onehotd[1]};
  assign lizzieLet4_4MQNode_4QNode_Bool_d = {lizzieLet4_6MQNode_d[16:1],
                                             lizzieLet4_6MQNode_onehotd[2]};
  assign lizzieLet4_4MQNode_4QError_Bool_d = {lizzieLet4_6MQNode_d[16:1],
                                              lizzieLet4_6MQNode_onehotd[3]};
  assign lizzieLet4_6MQNode_r = (| (lizzieLet4_6MQNode_onehotd & {lizzieLet4_4MQNode_4QError_Bool_r,
                                                                  lizzieLet4_4MQNode_4QNode_Bool_r,
                                                                  lizzieLet4_4MQNode_4QVal_Bool_r,
                                                                  lizzieLet4_4MQNode_4QNone_Bool_r}));
  assign lizzieLet4_4MQNode_4_r = lizzieLet4_6MQNode_r;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_4MQNode_4QError_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet4_4MQNode_4QError_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QError_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_4QError_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_4QError_Bool_r = ((! lizzieLet4_4MQNode_4QError_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4MQNode_4QError_Bool_r)
        lizzieLet4_4MQNode_4QError_Bool_bufchan_d <= lizzieLet4_4MQNode_4QError_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QError_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_4QError_Bool_bufchan_r = (! lizzieLet4_4MQNode_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_4QError_Bool_1_argbuf_d = (lizzieLet4_4MQNode_4QError_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_4QError_Bool_bufchan_buf :
                                                       lizzieLet4_4MQNode_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4MQNode_4QError_Bool_1_argbuf_r && lizzieLet4_4MQNode_4QError_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4MQNode_4QError_Bool_1_argbuf_r) && (! lizzieLet4_4MQNode_4QError_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_4QError_Bool_bufchan_buf <= lizzieLet4_4MQNode_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool3) : [(lizzieLet4_4MQNode_4QNode_Bool,Pointer_CTmain_mask_Bool),
                                     (t1acp_destruct,Pointer_QTree_Bool),
                                     (lizzieLet4_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                     (t2acq_destruct,Pointer_QTree_Bool),
                                     (lizzieLet4_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                     (t3acr_destruct,Pointer_QTree_Bool),
                                     (lizzieLet4_4MQNode_7QNode_Bool,Pointer_MaskQTree)] > (lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3,CTmain_mask_Bool) */
  assign lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d = Lcall_main_mask_Bool3_dc((& {lizzieLet4_4MQNode_4QNode_Bool_d[0],
                                                                                                                                                                                                                     t1acp_destruct_d[0],
                                                                                                                                                                                                                     lizzieLet4_4MQNode_5QNode_Bool_d[0],
                                                                                                                                                                                                                     t2acq_destruct_d[0],
                                                                                                                                                                                                                     lizzieLet4_4MQNode_6QNode_Bool_d[0],
                                                                                                                                                                                                                     t3acr_destruct_d[0],
                                                                                                                                                                                                                     lizzieLet4_4MQNode_7QNode_Bool_d[0]}), lizzieLet4_4MQNode_4QNode_Bool_d, t1acp_destruct_d, lizzieLet4_4MQNode_5QNode_Bool_d, t2acq_destruct_d, lizzieLet4_4MQNode_6QNode_Bool_d, t3acr_destruct_d, lizzieLet4_4MQNode_7QNode_Bool_d);
  assign {lizzieLet4_4MQNode_4QNode_Bool_r,
          t1acp_destruct_r,
          lizzieLet4_4MQNode_5QNode_Bool_r,
          t2acq_destruct_r,
          lizzieLet4_4MQNode_6QNode_Bool_r,
          t3acr_destruct_r,
          lizzieLet4_4MQNode_7QNode_Bool_r} = {7 {(lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r && lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3,CTmain_mask_Bool) > (lizzieLet9_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d;
  logic lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r;
  assign lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r = ((! lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d[0]) || lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d <= {115'd0,
                                                                                                                                                                                               1'd0};
    else
      if (lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r)
        lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d <= lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d;
  CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf;
  assign lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r = (! lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0] ? lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf :
                                  lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0]))
        lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                   1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0])))
        lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= lizzieLet4_4MQNode_4QNode_Bool_1t1acp_1lizzieLet4_4MQNode_5QNode_Bool_1t2acq_1lizzieLet4_4MQNode_6QNode_Bool_1t3acr_1lizzieLet4_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_4MQNode_4QNone_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet4_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNone_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_4QNone_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_4QNone_Bool_r = ((! lizzieLet4_4MQNode_4QNone_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4MQNode_4QNone_Bool_r)
        lizzieLet4_4MQNode_4QNone_Bool_bufchan_d <= lizzieLet4_4MQNode_4QNone_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_4QNone_Bool_bufchan_r = (! lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_d = (lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf :
                                                      lizzieLet4_4MQNode_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_r && lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4MQNode_4QNone_Bool_1_argbuf_r) && (! lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_4QNone_Bool_bufchan_buf <= lizzieLet4_4MQNode_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_4MQNode_4QVal_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet4_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QVal_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_4QVal_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_4QVal_Bool_r = ((! lizzieLet4_4MQNode_4QVal_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4MQNode_4QVal_Bool_r)
        lizzieLet4_4MQNode_4QVal_Bool_bufchan_d <= lizzieLet4_4MQNode_4QVal_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_4QVal_Bool_bufchan_r = (! lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_d = (lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf :
                                                     lizzieLet4_4MQNode_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_r && lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4MQNode_4QVal_Bool_1_argbuf_r) && (! lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_4QVal_Bool_bufchan_buf <= lizzieLet4_4MQNode_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet4_4MQNode_5,QTree_Bool) (q1ack_destruct,Pointer_MaskQTree) > [(_13,Pointer_MaskQTree),
                                                                                                       (_12,Pointer_MaskQTree),
                                                                                                       (lizzieLet4_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_11,Pointer_MaskQTree)] */
  logic [3:0] q1ack_destruct_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_5_d[0] && q1ack_destruct_d[0]))
      unique case (lizzieLet4_4MQNode_5_d[2:1])
        2'd0: q1ack_destruct_onehotd = 4'd1;
        2'd1: q1ack_destruct_onehotd = 4'd2;
        2'd2: q1ack_destruct_onehotd = 4'd4;
        2'd3: q1ack_destruct_onehotd = 4'd8;
        default: q1ack_destruct_onehotd = 4'd0;
      endcase
    else q1ack_destruct_onehotd = 4'd0;
  assign _13_d = {q1ack_destruct_d[16:1], q1ack_destruct_onehotd[0]};
  assign _12_d = {q1ack_destruct_d[16:1], q1ack_destruct_onehotd[1]};
  assign lizzieLet4_4MQNode_5QNode_Bool_d = {q1ack_destruct_d[16:1],
                                             q1ack_destruct_onehotd[2]};
  assign _11_d = {q1ack_destruct_d[16:1], q1ack_destruct_onehotd[3]};
  assign q1ack_destruct_r = (| (q1ack_destruct_onehotd & {_11_r,
                                                          lizzieLet4_4MQNode_5QNode_Bool_r,
                                                          _12_r,
                                                          _13_r}));
  assign lizzieLet4_4MQNode_5_r = q1ack_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet4_4MQNode_6,QTree_Bool) (q2acl_destruct,Pointer_MaskQTree) > [(_10,Pointer_MaskQTree),
                                                                                                       (_9,Pointer_MaskQTree),
                                                                                                       (lizzieLet4_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_8,Pointer_MaskQTree)] */
  logic [3:0] q2acl_destruct_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_6_d[0] && q2acl_destruct_d[0]))
      unique case (lizzieLet4_4MQNode_6_d[2:1])
        2'd0: q2acl_destruct_onehotd = 4'd1;
        2'd1: q2acl_destruct_onehotd = 4'd2;
        2'd2: q2acl_destruct_onehotd = 4'd4;
        2'd3: q2acl_destruct_onehotd = 4'd8;
        default: q2acl_destruct_onehotd = 4'd0;
      endcase
    else q2acl_destruct_onehotd = 4'd0;
  assign _10_d = {q2acl_destruct_d[16:1], q2acl_destruct_onehotd[0]};
  assign _9_d = {q2acl_destruct_d[16:1], q2acl_destruct_onehotd[1]};
  assign lizzieLet4_4MQNode_6QNode_Bool_d = {q2acl_destruct_d[16:1],
                                             q2acl_destruct_onehotd[2]};
  assign _8_d = {q2acl_destruct_d[16:1], q2acl_destruct_onehotd[3]};
  assign q2acl_destruct_r = (| (q2acl_destruct_onehotd & {_8_r,
                                                          lizzieLet4_4MQNode_6QNode_Bool_r,
                                                          _9_r,
                                                          _10_r}));
  assign lizzieLet4_4MQNode_6_r = q2acl_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet4_4MQNode_7,QTree_Bool) (q3acm_destruct,Pointer_MaskQTree) > [(_7,Pointer_MaskQTree),
                                                                                                       (_6,Pointer_MaskQTree),
                                                                                                       (lizzieLet4_4MQNode_7QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_5,Pointer_MaskQTree)] */
  logic [3:0] q3acm_destruct_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_7_d[0] && q3acm_destruct_d[0]))
      unique case (lizzieLet4_4MQNode_7_d[2:1])
        2'd0: q3acm_destruct_onehotd = 4'd1;
        2'd1: q3acm_destruct_onehotd = 4'd2;
        2'd2: q3acm_destruct_onehotd = 4'd4;
        2'd3: q3acm_destruct_onehotd = 4'd8;
        default: q3acm_destruct_onehotd = 4'd0;
      endcase
    else q3acm_destruct_onehotd = 4'd0;
  assign _7_d = {q3acm_destruct_d[16:1], q3acm_destruct_onehotd[0]};
  assign _6_d = {q3acm_destruct_d[16:1], q3acm_destruct_onehotd[1]};
  assign lizzieLet4_4MQNode_7QNode_Bool_d = {q3acm_destruct_d[16:1],
                                             q3acm_destruct_onehotd[2]};
  assign _5_d = {q3acm_destruct_d[16:1], q3acm_destruct_onehotd[3]};
  assign q3acm_destruct_r = (| (q3acm_destruct_onehotd & {_5_r,
                                                          lizzieLet4_4MQNode_7QNode_Bool_r,
                                                          _6_r,
                                                          _7_r}));
  assign lizzieLet4_4MQNode_7_r = q3acm_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet4_4MQNode_8,QTree_Bool) (q4acn_destruct,Pointer_MaskQTree) > [(_4,Pointer_MaskQTree),
                                                                                                       (_3,Pointer_MaskQTree),
                                                                                                       (lizzieLet4_4MQNode_8QNode_Bool,Pointer_MaskQTree),
                                                                                                       (_2,Pointer_MaskQTree)] */
  logic [3:0] q4acn_destruct_onehotd;
  always_comb
    if ((lizzieLet4_4MQNode_8_d[0] && q4acn_destruct_d[0]))
      unique case (lizzieLet4_4MQNode_8_d[2:1])
        2'd0: q4acn_destruct_onehotd = 4'd1;
        2'd1: q4acn_destruct_onehotd = 4'd2;
        2'd2: q4acn_destruct_onehotd = 4'd4;
        2'd3: q4acn_destruct_onehotd = 4'd8;
        default: q4acn_destruct_onehotd = 4'd0;
      endcase
    else q4acn_destruct_onehotd = 4'd0;
  assign _4_d = {q4acn_destruct_d[16:1], q4acn_destruct_onehotd[0]};
  assign _3_d = {q4acn_destruct_d[16:1], q4acn_destruct_onehotd[1]};
  assign lizzieLet4_4MQNode_8QNode_Bool_d = {q4acn_destruct_d[16:1],
                                             q4acn_destruct_onehotd[2]};
  assign _2_d = {q4acn_destruct_d[16:1], q4acn_destruct_onehotd[3]};
  assign q4acn_destruct_r = (| (q4acn_destruct_onehotd & {_2_r,
                                                          lizzieLet4_4MQNode_8QNode_Bool_r,
                                                          _3_r,
                                                          _4_r}));
  assign lizzieLet4_4MQNode_8_r = q4acn_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet4_4MQNode_8QNode_Bool,Pointer_MaskQTree) > (lizzieLet4_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet4_4MQNode_8QNode_Bool_bufchan_d;
  logic lizzieLet4_4MQNode_8QNode_Bool_bufchan_r;
  assign lizzieLet4_4MQNode_8QNode_Bool_r = ((! lizzieLet4_4MQNode_8QNode_Bool_bufchan_d[0]) || lizzieLet4_4MQNode_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_8QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4MQNode_8QNode_Bool_r)
        lizzieLet4_4MQNode_8QNode_Bool_bufchan_d <= lizzieLet4_4MQNode_8QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf;
  assign lizzieLet4_4MQNode_8QNode_Bool_bufchan_r = (! lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_d = (lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf[0] ? lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf :
                                                      lizzieLet4_4MQNode_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_r && lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf[0]))
        lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4MQNode_8QNode_Bool_1_argbuf_r) && (! lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf[0])))
        lizzieLet4_4MQNode_8QNode_Bool_bufchan_buf <= lizzieLet4_4MQNode_8QNode_Bool_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Bool) : (lizzieLet4_5,MaskQTree) (maci_2,Pointer_QTree_Bool) > [(_1,Pointer_QTree_Bool),
                                                                                        (lizzieLet4_5MQVal,Pointer_QTree_Bool),
                                                                                        (_0,Pointer_QTree_Bool)] */
  logic [2:0] maci_2_onehotd;
  always_comb
    if ((lizzieLet4_5_d[0] && maci_2_d[0]))
      unique case (lizzieLet4_5_d[2:1])
        2'd0: maci_2_onehotd = 3'd1;
        2'd1: maci_2_onehotd = 3'd2;
        2'd2: maci_2_onehotd = 3'd4;
        default: maci_2_onehotd = 3'd0;
      endcase
    else maci_2_onehotd = 3'd0;
  assign _1_d = {maci_2_d[16:1], maci_2_onehotd[0]};
  assign lizzieLet4_5MQVal_d = {maci_2_d[16:1], maci_2_onehotd[1]};
  assign _0_d = {maci_2_d[16:1], maci_2_onehotd[2]};
  assign maci_2_r = (| (maci_2_onehotd & {_0_r,
                                          lizzieLet4_5MQVal_r,
                                          _1_r}));
  assign lizzieLet4_5_r = maci_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet4_5MQVal,Pointer_QTree_Bool) > (lizzieLet4_5MQVal_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet4_5MQVal_bufchan_d;
  logic lizzieLet4_5MQVal_bufchan_r;
  assign lizzieLet4_5MQVal_r = ((! lizzieLet4_5MQVal_bufchan_d[0]) || lizzieLet4_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_5MQVal_r)
        lizzieLet4_5MQVal_bufchan_d <= lizzieLet4_5MQVal_d;
  Pointer_QTree_Bool_t lizzieLet4_5MQVal_bufchan_buf;
  assign lizzieLet4_5MQVal_bufchan_r = (! lizzieLet4_5MQVal_bufchan_buf[0]);
  assign lizzieLet4_5MQVal_1_argbuf_d = (lizzieLet4_5MQVal_bufchan_buf[0] ? lizzieLet4_5MQVal_bufchan_buf :
                                         lizzieLet4_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_5MQVal_1_argbuf_r && lizzieLet4_5MQVal_bufchan_buf[0]))
        lizzieLet4_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_5MQVal_1_argbuf_r) && (! lizzieLet4_5MQVal_bufchan_buf[0])))
        lizzieLet4_5MQVal_bufchan_buf <= lizzieLet4_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_6,MaskQTree) (sc_0_1_goMux_mux,Pointer_CTmain_mask_Bool) > [(lizzieLet4_6MQNone,Pointer_CTmain_mask_Bool),
                                                                                                              (lizzieLet4_6MQVal,Pointer_CTmain_mask_Bool),
                                                                                                              (lizzieLet4_6MQNode,Pointer_CTmain_mask_Bool)] */
  logic [2:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet4_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 3'd4;
        default: sc_0_1_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 3'd0;
  assign lizzieLet4_6MQNone_d = {sc_0_1_goMux_mux_d[16:1],
                                 sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet4_6MQVal_d = {sc_0_1_goMux_mux_d[16:1],
                                sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet4_6MQNode_d = {sc_0_1_goMux_mux_d[16:1],
                                 sc_0_1_goMux_mux_onehotd[2]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet4_6MQNode_r,
                                                              lizzieLet4_6MQVal_r,
                                                              lizzieLet4_6MQNone_r}));
  assign lizzieLet4_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_6MQNone,Pointer_CTmain_mask_Bool) > (lizzieLet4_6MQNone_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQNone_bufchan_d;
  logic lizzieLet4_6MQNone_bufchan_r;
  assign lizzieLet4_6MQNone_r = ((! lizzieLet4_6MQNone_bufchan_d[0]) || lizzieLet4_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_6MQNone_r)
        lizzieLet4_6MQNone_bufchan_d <= lizzieLet4_6MQNone_d;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQNone_bufchan_buf;
  assign lizzieLet4_6MQNone_bufchan_r = (! lizzieLet4_6MQNone_bufchan_buf[0]);
  assign lizzieLet4_6MQNone_1_argbuf_d = (lizzieLet4_6MQNone_bufchan_buf[0] ? lizzieLet4_6MQNone_bufchan_buf :
                                          lizzieLet4_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_6MQNone_1_argbuf_r && lizzieLet4_6MQNone_bufchan_buf[0]))
        lizzieLet4_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_6MQNone_1_argbuf_r) && (! lizzieLet4_6MQNone_bufchan_buf[0])))
        lizzieLet4_6MQNone_bufchan_buf <= lizzieLet4_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet4_6MQVal,Pointer_CTmain_mask_Bool) > (lizzieLet4_6MQVal_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQVal_bufchan_d;
  logic lizzieLet4_6MQVal_bufchan_r;
  assign lizzieLet4_6MQVal_r = ((! lizzieLet4_6MQVal_bufchan_d[0]) || lizzieLet4_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_6MQVal_r)
        lizzieLet4_6MQVal_bufchan_d <= lizzieLet4_6MQVal_d;
  Pointer_CTmain_mask_Bool_t lizzieLet4_6MQVal_bufchan_buf;
  assign lizzieLet4_6MQVal_bufchan_r = (! lizzieLet4_6MQVal_bufchan_buf[0]);
  assign lizzieLet4_6MQVal_1_argbuf_d = (lizzieLet4_6MQVal_bufchan_buf[0] ? lizzieLet4_6MQVal_bufchan_buf :
                                         lizzieLet4_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_6MQVal_1_argbuf_r && lizzieLet4_6MQVal_bufchan_buf[0]))
        lizzieLet4_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_6MQVal_1_argbuf_r) && (! lizzieLet4_6MQVal_bufchan_buf[0])))
        lizzieLet4_6MQVal_bufchan_buf <= lizzieLet4_6MQVal_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (m1acL_goMux_mux,Pointer_QTree_Bool) > (m1acL_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m1acL_goMux_mux_bufchan_d;
  logic m1acL_goMux_mux_bufchan_r;
  assign m1acL_goMux_mux_r = ((! m1acL_goMux_mux_bufchan_d[0]) || m1acL_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acL_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1acL_goMux_mux_r)
        m1acL_goMux_mux_bufchan_d <= m1acL_goMux_mux_d;
  Pointer_QTree_Bool_t m1acL_goMux_mux_bufchan_buf;
  assign m1acL_goMux_mux_bufchan_r = (! m1acL_goMux_mux_bufchan_buf[0]);
  assign m1acL_1_argbuf_d = (m1acL_goMux_mux_bufchan_buf[0] ? m1acL_goMux_mux_bufchan_buf :
                             m1acL_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acL_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1acL_1_argbuf_r && m1acL_goMux_mux_bufchan_buf[0]))
        m1acL_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1acL_1_argbuf_r) && (! m1acL_goMux_mux_bufchan_buf[0])))
        m1acL_goMux_mux_bufchan_buf <= m1acL_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (m2acM_2_2,Pointer_QTree_Bool) > (m2acM_2_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2acM_2_2_bufchan_d;
  logic m2acM_2_2_bufchan_r;
  assign m2acM_2_2_r = ((! m2acM_2_2_bufchan_d[0]) || m2acM_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_2_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2acM_2_2_r) m2acM_2_2_bufchan_d <= m2acM_2_2_d;
  Pointer_QTree_Bool_t m2acM_2_2_bufchan_buf;
  assign m2acM_2_2_bufchan_r = (! m2acM_2_2_bufchan_buf[0]);
  assign m2acM_2_2_argbuf_d = (m2acM_2_2_bufchan_buf[0] ? m2acM_2_2_bufchan_buf :
                               m2acM_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_2_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acM_2_2_argbuf_r && m2acM_2_2_bufchan_buf[0]))
        m2acM_2_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acM_2_2_argbuf_r) && (! m2acM_2_2_bufchan_buf[0])))
        m2acM_2_2_bufchan_buf <= m2acM_2_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2acM_2_destruct,Pointer_QTree_Bool) > [(m2acM_2_1,Pointer_QTree_Bool),
                                                                        (m2acM_2_2,Pointer_QTree_Bool)] */
  logic [1:0] m2acM_2_destruct_emitted;
  logic [1:0] m2acM_2_destruct_done;
  assign m2acM_2_1_d = {m2acM_2_destruct_d[16:1],
                        (m2acM_2_destruct_d[0] && (! m2acM_2_destruct_emitted[0]))};
  assign m2acM_2_2_d = {m2acM_2_destruct_d[16:1],
                        (m2acM_2_destruct_d[0] && (! m2acM_2_destruct_emitted[1]))};
  assign m2acM_2_destruct_done = (m2acM_2_destruct_emitted | ({m2acM_2_2_d[0],
                                                               m2acM_2_1_d[0]} & {m2acM_2_2_r,
                                                                                  m2acM_2_1_r}));
  assign m2acM_2_destruct_r = (& m2acM_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_2_destruct_emitted <= 2'd0;
    else
      m2acM_2_destruct_emitted <= (m2acM_2_destruct_r ? 2'd0 :
                                   m2acM_2_destruct_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2acM_3_2,Pointer_QTree_Bool) > (m2acM_3_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2acM_3_2_bufchan_d;
  logic m2acM_3_2_bufchan_r;
  assign m2acM_3_2_r = ((! m2acM_3_2_bufchan_d[0]) || m2acM_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_3_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2acM_3_2_r) m2acM_3_2_bufchan_d <= m2acM_3_2_d;
  Pointer_QTree_Bool_t m2acM_3_2_bufchan_buf;
  assign m2acM_3_2_bufchan_r = (! m2acM_3_2_bufchan_buf[0]);
  assign m2acM_3_2_argbuf_d = (m2acM_3_2_bufchan_buf[0] ? m2acM_3_2_bufchan_buf :
                               m2acM_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_3_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acM_3_2_argbuf_r && m2acM_3_2_bufchan_buf[0]))
        m2acM_3_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acM_3_2_argbuf_r) && (! m2acM_3_2_bufchan_buf[0])))
        m2acM_3_2_bufchan_buf <= m2acM_3_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2acM_3_destruct,Pointer_QTree_Bool) > [(m2acM_3_1,Pointer_QTree_Bool),
                                                                        (m2acM_3_2,Pointer_QTree_Bool)] */
  logic [1:0] m2acM_3_destruct_emitted;
  logic [1:0] m2acM_3_destruct_done;
  assign m2acM_3_1_d = {m2acM_3_destruct_d[16:1],
                        (m2acM_3_destruct_d[0] && (! m2acM_3_destruct_emitted[0]))};
  assign m2acM_3_2_d = {m2acM_3_destruct_d[16:1],
                        (m2acM_3_destruct_d[0] && (! m2acM_3_destruct_emitted[1]))};
  assign m2acM_3_destruct_done = (m2acM_3_destruct_emitted | ({m2acM_3_2_d[0],
                                                               m2acM_3_1_d[0]} & {m2acM_3_2_r,
                                                                                  m2acM_3_1_r}));
  assign m2acM_3_destruct_r = (& m2acM_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_3_destruct_emitted <= 2'd0;
    else
      m2acM_3_destruct_emitted <= (m2acM_3_destruct_r ? 2'd0 :
                                   m2acM_3_destruct_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2acM_4_destruct,Pointer_QTree_Bool) > (m2acM_4_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2acM_4_destruct_bufchan_d;
  logic m2acM_4_destruct_bufchan_r;
  assign m2acM_4_destruct_r = ((! m2acM_4_destruct_bufchan_d[0]) || m2acM_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2acM_4_destruct_r)
        m2acM_4_destruct_bufchan_d <= m2acM_4_destruct_d;
  Pointer_QTree_Bool_t m2acM_4_destruct_bufchan_buf;
  assign m2acM_4_destruct_bufchan_r = (! m2acM_4_destruct_bufchan_buf[0]);
  assign m2acM_4_1_argbuf_d = (m2acM_4_destruct_bufchan_buf[0] ? m2acM_4_destruct_bufchan_buf :
                               m2acM_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acM_4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acM_4_1_argbuf_r && m2acM_4_destruct_bufchan_buf[0]))
        m2acM_4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acM_4_1_argbuf_r) && (! m2acM_4_destruct_bufchan_buf[0])))
        m2acM_4_destruct_bufchan_buf <= m2acM_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (macD_goMux_mux,Pointer_QTree_Bool) > (macD_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t macD_goMux_mux_bufchan_d;
  logic macD_goMux_mux_bufchan_r;
  assign macD_goMux_mux_r = ((! macD_goMux_mux_bufchan_d[0]) || macD_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macD_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (macD_goMux_mux_r) macD_goMux_mux_bufchan_d <= macD_goMux_mux_d;
  Pointer_QTree_Bool_t macD_goMux_mux_bufchan_buf;
  assign macD_goMux_mux_bufchan_r = (! macD_goMux_mux_bufchan_buf[0]);
  assign macD_1_argbuf_d = (macD_goMux_mux_bufchan_buf[0] ? macD_goMux_mux_bufchan_buf :
                            macD_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macD_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((macD_1_argbuf_r && macD_goMux_mux_bufchan_buf[0]))
        macD_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! macD_1_argbuf_r) && (! macD_goMux_mux_bufchan_buf[0])))
        macD_goMux_mux_bufchan_buf <= macD_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (maci_1,Pointer_QTree_Bool) > (maci_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t maci_1_bufchan_d;
  logic maci_1_bufchan_r;
  assign maci_1_r = ((! maci_1_bufchan_d[0]) || maci_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) maci_1_bufchan_d <= {16'd0, 1'd0};
    else if (maci_1_r) maci_1_bufchan_d <= maci_1_d;
  Pointer_QTree_Bool_t maci_1_bufchan_buf;
  assign maci_1_bufchan_r = (! maci_1_bufchan_buf[0]);
  assign maci_1_argbuf_d = (maci_1_bufchan_buf[0] ? maci_1_bufchan_buf :
                            maci_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) maci_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((maci_1_argbuf_r && maci_1_bufchan_buf[0]))
        maci_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! maci_1_argbuf_r) && (! maci_1_bufchan_buf[0])))
        maci_1_bufchan_buf <= maci_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (maci_goMux_mux,Pointer_QTree_Bool) > [(maci_1,Pointer_QTree_Bool),
                                                                      (maci_2,Pointer_QTree_Bool)] */
  logic [1:0] maci_goMux_mux_emitted;
  logic [1:0] maci_goMux_mux_done;
  assign maci_1_d = {maci_goMux_mux_d[16:1],
                     (maci_goMux_mux_d[0] && (! maci_goMux_mux_emitted[0]))};
  assign maci_2_d = {maci_goMux_mux_d[16:1],
                     (maci_goMux_mux_d[0] && (! maci_goMux_mux_emitted[1]))};
  assign maci_goMux_mux_done = (maci_goMux_mux_emitted | ({maci_2_d[0],
                                                           maci_1_d[0]} & {maci_2_r, maci_1_r}));
  assign maci_goMux_mux_r = (& maci_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) maci_goMux_mux_emitted <= 2'd0;
    else
      maci_goMux_mux_emitted <= (maci_goMux_mux_r ? 2'd0 :
                                 maci_goMux_mux_done);
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) > [(main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8,Go),
                                                                                                                                                                                    (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1,Pointer_QTree_Bool),
                                                                                                                                                                                    (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1,Pointer_MaskQTree)] */
  logic [2:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted;
  logic [2:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[0]));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_d = {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[16:1],
                                                                                 (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[1]))};
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_d = {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[32:17],
                                                                                   (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[2]))};
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted | ({main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_d[0],
                                                                                                                                                           main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_d[0],
                                                                                                                                                           main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_d[0]} & {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_r,
                                                                                                                                                                                                                                     main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_r,
                                                                                                                                                                                                                                     main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_r}));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r = (& main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted <= 3'd0;
    else
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted <= (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r ? 3'd0 :
                                                                                 main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done);
  
  /* fork (Ty Go) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8,Go) > [(go_8_1,Go),
                                                                                        (go_8_2,Go)] */
  logic [1:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted;
  logic [1:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_done;
  assign go_8_1_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted[0]));
  assign go_8_2_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted[1]));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_done = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted | ({go_8_2_d[0],
                                                                                                                                                               go_8_1_d[0]} & {go_8_2_r,
                                                                                                                                                                               go_8_1_r}));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_r = (& main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted <= 2'd0;
    else
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_emitted <= (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_r ? 2'd0 :
                                                                                   main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_8_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1,Pointer_QTree_Bool) > (maci_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_r;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_r = ((! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d[0]) || main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d <= {16'd0,
                                                                                       1'd0};
    else
      if (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_r)
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_d;
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_r = (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf[0]);
  assign maci_1_1_argbuf_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf[0] ? main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf :
                              main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
    else
      if ((maci_1_1_argbuf_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf[0]))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
      else if (((! maci_1_1_argbuf_r) && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf[0])))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_buf <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemaci_1_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1,Pointer_MaskQTree) > (mskacj_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_r;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_r = ((! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d[0]) || main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d <= {16'd0,
                                                                                         1'd0};
    else
      if (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_r)
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_d;
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_r = (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf[0]);
  assign mskacj_1_1_argbuf_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf[0] ? main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf :
                                main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
    else
      if ((mskacj_1_1_argbuf_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf[0]))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf <= {16'd0,
                                                                                             1'd0};
      else if (((! mskacj_1_1_argbuf_r) && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf[0])))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_buf <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemskacj_1_bufchan_d;
  
  /* sink (Ty Pointer_QTree_Bool) : (main_mask_Bool_resbuf,Pointer_QTree_Bool) > */
  assign {main_mask_Bool_resbuf_r,
          main_mask_Bool_resbuf_dout} = {main_mask_Bool_resbuf_rout,
                                         main_mask_Bool_resbuf_d};
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) > [(map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9,Go),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1,MyDTBool_Bool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1,MyBool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1,Pointer_QTree_Bool)] */
  logic [4:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted ;
  logic [4:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [0]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [1]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [2]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_d  = {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [1:1],
                                                                                                                          (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [3]))};
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_d  = {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [17:2],
                                                                                                                         (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [4]))};
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  | ({\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_d [0]} & {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_r ,
                                                                                                                                                                                                                                                                                                                                                             \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_r ,
                                                                                                                                                                                                                                                                                                                                                             \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_r ,
                                                                                                                                                                                                                                                                                                                                                             \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_r ,
                                                                                                                                                                                                                                                                                                                                                             \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_r }));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  = (& \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  <= 5'd0;
    else
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  <= (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  ? 5'd0 :
                                                                                                                         \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done );
  
  /* buf (Ty MyDTBool_Bool_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1,MyDTBool_Bool_Bool) > (gacB_1_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_d ;
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf [0]);
  assign gacB_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf  :
                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf  <= 1'd0;
    else
      if ((gacB_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf  <= 1'd0;
      else if (((! gacB_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacB_1_bufchan_d ;
  
  /* fork (Ty Go) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9,Go) > [(go_9_1,Go),
                                                                                                                              (go_9_2,Go)] */
  logic [1:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted ;
  logic [1:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_done ;
  assign go_9_1_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted [0]));
  assign go_9_2_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted [1]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_done  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted  | ({go_9_2_d[0],
                                                                                                                                                                                                                                               go_9_1_d[0]} & {go_9_2_r,
                                                                                                                                                                                                                                                               go_9_1_r}));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_r  = (& \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted  <= 2'd0;
    else
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_emitted  <= (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_r  ? 2'd0 :
                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_9_done );
  
  /* buf (Ty MyDTBool_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1,MyDTBool_Bool) > (isZacA_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_d ;
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf [0]);
  assign isZacA_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf  :
                                \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacA_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf  <= 1'd0;
      else if (((! isZacA_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacA_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1,Pointer_QTree_Bool) > (macD_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d  <= {16'd0,
                                                                                                                               1'd0};
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_d ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf [0]);
  assign macD_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf  :
                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf  <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((macD_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf  <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! macD_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolmacD_1_bufchan_d ;
  
  /* buf (Ty MyBool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1,MyBool) > (v'acC_1_1_argbuf,MyBool) */
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d  <= {1'd0,
                                                                                                                                1'd0};
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_d ;
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf [0]);
  assign \v'acC_1_1_argbuf_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf  :
                                 \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf  <= {1'd0,
                                                                                                                                  1'd0};
    else
      if ((\v'acC_1_1_argbuf_r  && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf  <= {1'd0,
                                                                                                                                    1'd0};
      else if (((! \v'acC_1_1_argbuf_r ) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'acC_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (map''_map''_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) > (lizzieLet11_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d ;
  logic \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r ;
  assign \map''_map''_Bool_Bool_Bool_resbuf_r  = ((! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d [0]) || \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\map''_map''_Bool_Bool_Bool_resbuf_r )
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d  <= \map''_map''_Bool_Bool_Bool_resbuf_d ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf ;
  assign \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r  = (! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0]);
  assign lizzieLet11_1_argbuf_d = (\map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0] ? \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  :
                                   \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0]))
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0])))
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (mskacj_goMux_mux,Pointer_MaskQTree) > (mskacj_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t mskacj_goMux_mux_bufchan_d;
  logic mskacj_goMux_mux_bufchan_r;
  assign mskacj_goMux_mux_r = ((! mskacj_goMux_mux_bufchan_d[0]) || mskacj_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mskacj_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (mskacj_goMux_mux_r)
        mskacj_goMux_mux_bufchan_d <= mskacj_goMux_mux_d;
  Pointer_MaskQTree_t mskacj_goMux_mux_bufchan_buf;
  assign mskacj_goMux_mux_bufchan_r = (! mskacj_goMux_mux_bufchan_buf[0]);
  assign mskacj_1_argbuf_d = (mskacj_goMux_mux_bufchan_buf[0] ? mskacj_goMux_mux_bufchan_buf :
                              mskacj_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mskacj_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mskacj_1_argbuf_r && mskacj_goMux_mux_bufchan_buf[0]))
        mskacj_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mskacj_1_argbuf_r) && (! mskacj_goMux_mux_bufchan_buf[0])))
        mskacj_goMux_mux_bufchan_buf <= mskacj_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1acF_3_destruct,Pointer_QTree_Bool) > (q1acF_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1acF_3_destruct_bufchan_d;
  logic q1acF_3_destruct_bufchan_r;
  assign q1acF_3_destruct_r = ((! q1acF_3_destruct_bufchan_d[0]) || q1acF_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acF_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acF_3_destruct_r)
        q1acF_3_destruct_bufchan_d <= q1acF_3_destruct_d;
  Pointer_QTree_Bool_t q1acF_3_destruct_bufchan_buf;
  assign q1acF_3_destruct_bufchan_r = (! q1acF_3_destruct_bufchan_buf[0]);
  assign q1acF_3_1_argbuf_d = (q1acF_3_destruct_bufchan_buf[0] ? q1acF_3_destruct_bufchan_buf :
                               q1acF_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acF_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acF_3_1_argbuf_r && q1acF_3_destruct_bufchan_buf[0]))
        q1acF_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acF_3_1_argbuf_r) && (! q1acF_3_destruct_bufchan_buf[0])))
        q1acF_3_destruct_bufchan_buf <= q1acF_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1acO_3_destruct,Pointer_QTree_Bool) > (q1acO_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1acO_3_destruct_bufchan_d;
  logic q1acO_3_destruct_bufchan_r;
  assign q1acO_3_destruct_r = ((! q1acO_3_destruct_bufchan_d[0]) || q1acO_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acO_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acO_3_destruct_r)
        q1acO_3_destruct_bufchan_d <= q1acO_3_destruct_d;
  Pointer_QTree_Bool_t q1acO_3_destruct_bufchan_buf;
  assign q1acO_3_destruct_bufchan_r = (! q1acO_3_destruct_bufchan_buf[0]);
  assign q1acO_3_1_argbuf_d = (q1acO_3_destruct_bufchan_buf[0] ? q1acO_3_destruct_bufchan_buf :
                               q1acO_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acO_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acO_3_1_argbuf_r && q1acO_3_destruct_bufchan_buf[0]))
        q1acO_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acO_3_1_argbuf_r) && (! q1acO_3_destruct_bufchan_buf[0])))
        q1acO_3_destruct_bufchan_buf <= q1acO_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1ack_3_destruct,Pointer_MaskQTree) > (q1ack_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1ack_3_destruct_bufchan_d;
  logic q1ack_3_destruct_bufchan_r;
  assign q1ack_3_destruct_r = ((! q1ack_3_destruct_bufchan_d[0]) || q1ack_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ack_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ack_3_destruct_r)
        q1ack_3_destruct_bufchan_d <= q1ack_3_destruct_d;
  Pointer_MaskQTree_t q1ack_3_destruct_bufchan_buf;
  assign q1ack_3_destruct_bufchan_r = (! q1ack_3_destruct_bufchan_buf[0]);
  assign q1ack_3_1_argbuf_d = (q1ack_3_destruct_bufchan_buf[0] ? q1ack_3_destruct_bufchan_buf :
                               q1ack_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ack_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ack_3_1_argbuf_r && q1ack_3_destruct_bufchan_buf[0]))
        q1ack_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ack_3_1_argbuf_r) && (! q1ack_3_destruct_bufchan_buf[0])))
        q1ack_3_destruct_bufchan_buf <= q1ack_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2acG_2_destruct,Pointer_QTree_Bool) > (q2acG_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2acG_2_destruct_bufchan_d;
  logic q2acG_2_destruct_bufchan_r;
  assign q2acG_2_destruct_r = ((! q2acG_2_destruct_bufchan_d[0]) || q2acG_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acG_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acG_2_destruct_r)
        q2acG_2_destruct_bufchan_d <= q2acG_2_destruct_d;
  Pointer_QTree_Bool_t q2acG_2_destruct_bufchan_buf;
  assign q2acG_2_destruct_bufchan_r = (! q2acG_2_destruct_bufchan_buf[0]);
  assign q2acG_2_1_argbuf_d = (q2acG_2_destruct_bufchan_buf[0] ? q2acG_2_destruct_bufchan_buf :
                               q2acG_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acG_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acG_2_1_argbuf_r && q2acG_2_destruct_bufchan_buf[0]))
        q2acG_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acG_2_1_argbuf_r) && (! q2acG_2_destruct_bufchan_buf[0])))
        q2acG_2_destruct_bufchan_buf <= q2acG_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2acP_2_destruct,Pointer_QTree_Bool) > (q2acP_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2acP_2_destruct_bufchan_d;
  logic q2acP_2_destruct_bufchan_r;
  assign q2acP_2_destruct_r = ((! q2acP_2_destruct_bufchan_d[0]) || q2acP_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acP_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acP_2_destruct_r)
        q2acP_2_destruct_bufchan_d <= q2acP_2_destruct_d;
  Pointer_QTree_Bool_t q2acP_2_destruct_bufchan_buf;
  assign q2acP_2_destruct_bufchan_r = (! q2acP_2_destruct_bufchan_buf[0]);
  assign q2acP_2_1_argbuf_d = (q2acP_2_destruct_bufchan_buf[0] ? q2acP_2_destruct_bufchan_buf :
                               q2acP_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acP_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acP_2_1_argbuf_r && q2acP_2_destruct_bufchan_buf[0]))
        q2acP_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acP_2_1_argbuf_r) && (! q2acP_2_destruct_bufchan_buf[0])))
        q2acP_2_destruct_bufchan_buf <= q2acP_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2acl_2_destruct,Pointer_MaskQTree) > (q2acl_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2acl_2_destruct_bufchan_d;
  logic q2acl_2_destruct_bufchan_r;
  assign q2acl_2_destruct_r = ((! q2acl_2_destruct_bufchan_d[0]) || q2acl_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acl_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acl_2_destruct_r)
        q2acl_2_destruct_bufchan_d <= q2acl_2_destruct_d;
  Pointer_MaskQTree_t q2acl_2_destruct_bufchan_buf;
  assign q2acl_2_destruct_bufchan_r = (! q2acl_2_destruct_bufchan_buf[0]);
  assign q2acl_2_1_argbuf_d = (q2acl_2_destruct_bufchan_buf[0] ? q2acl_2_destruct_bufchan_buf :
                               q2acl_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acl_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acl_2_1_argbuf_r && q2acl_2_destruct_bufchan_buf[0]))
        q2acl_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acl_2_1_argbuf_r) && (! q2acl_2_destruct_bufchan_buf[0])))
        q2acl_2_destruct_bufchan_buf <= q2acl_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3acH_1_destruct,Pointer_QTree_Bool) > (q3acH_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3acH_1_destruct_bufchan_d;
  logic q3acH_1_destruct_bufchan_r;
  assign q3acH_1_destruct_r = ((! q3acH_1_destruct_bufchan_d[0]) || q3acH_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acH_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acH_1_destruct_r)
        q3acH_1_destruct_bufchan_d <= q3acH_1_destruct_d;
  Pointer_QTree_Bool_t q3acH_1_destruct_bufchan_buf;
  assign q3acH_1_destruct_bufchan_r = (! q3acH_1_destruct_bufchan_buf[0]);
  assign q3acH_1_1_argbuf_d = (q3acH_1_destruct_bufchan_buf[0] ? q3acH_1_destruct_bufchan_buf :
                               q3acH_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acH_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acH_1_1_argbuf_r && q3acH_1_destruct_bufchan_buf[0]))
        q3acH_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acH_1_1_argbuf_r) && (! q3acH_1_destruct_bufchan_buf[0])))
        q3acH_1_destruct_bufchan_buf <= q3acH_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3acQ_1_destruct,Pointer_QTree_Bool) > (q3acQ_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3acQ_1_destruct_bufchan_d;
  logic q3acQ_1_destruct_bufchan_r;
  assign q3acQ_1_destruct_r = ((! q3acQ_1_destruct_bufchan_d[0]) || q3acQ_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acQ_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acQ_1_destruct_r)
        q3acQ_1_destruct_bufchan_d <= q3acQ_1_destruct_d;
  Pointer_QTree_Bool_t q3acQ_1_destruct_bufchan_buf;
  assign q3acQ_1_destruct_bufchan_r = (! q3acQ_1_destruct_bufchan_buf[0]);
  assign q3acQ_1_1_argbuf_d = (q3acQ_1_destruct_bufchan_buf[0] ? q3acQ_1_destruct_bufchan_buf :
                               q3acQ_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acQ_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acQ_1_1_argbuf_r && q3acQ_1_destruct_bufchan_buf[0]))
        q3acQ_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acQ_1_1_argbuf_r) && (! q3acQ_1_destruct_bufchan_buf[0])))
        q3acQ_1_destruct_bufchan_buf <= q3acQ_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3acm_1_destruct,Pointer_MaskQTree) > (q3acm_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3acm_1_destruct_bufchan_d;
  logic q3acm_1_destruct_bufchan_r;
  assign q3acm_1_destruct_r = ((! q3acm_1_destruct_bufchan_d[0]) || q3acm_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acm_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acm_1_destruct_r)
        q3acm_1_destruct_bufchan_d <= q3acm_1_destruct_d;
  Pointer_MaskQTree_t q3acm_1_destruct_bufchan_buf;
  assign q3acm_1_destruct_bufchan_r = (! q3acm_1_destruct_bufchan_buf[0]);
  assign q3acm_1_1_argbuf_d = (q3acm_1_destruct_bufchan_buf[0] ? q3acm_1_destruct_bufchan_buf :
                               q3acm_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acm_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acm_1_1_argbuf_r && q3acm_1_destruct_bufchan_buf[0]))
        q3acm_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acm_1_1_argbuf_r) && (! q3acm_1_destruct_bufchan_buf[0])))
        q3acm_1_destruct_bufchan_buf <= q3acm_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4acI_destruct,Pointer_QTree_Bool) > (q4acI_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4acI_destruct_bufchan_d;
  logic q4acI_destruct_bufchan_r;
  assign q4acI_destruct_r = ((! q4acI_destruct_bufchan_d[0]) || q4acI_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acI_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acI_destruct_r) q4acI_destruct_bufchan_d <= q4acI_destruct_d;
  Pointer_QTree_Bool_t q4acI_destruct_bufchan_buf;
  assign q4acI_destruct_bufchan_r = (! q4acI_destruct_bufchan_buf[0]);
  assign q4acI_1_argbuf_d = (q4acI_destruct_bufchan_buf[0] ? q4acI_destruct_bufchan_buf :
                             q4acI_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acI_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acI_1_argbuf_r && q4acI_destruct_bufchan_buf[0]))
        q4acI_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acI_1_argbuf_r) && (! q4acI_destruct_bufchan_buf[0])))
        q4acI_destruct_bufchan_buf <= q4acI_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4acR_destruct,Pointer_QTree_Bool) > (q4acR_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4acR_destruct_bufchan_d;
  logic q4acR_destruct_bufchan_r;
  assign q4acR_destruct_r = ((! q4acR_destruct_bufchan_d[0]) || q4acR_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acR_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acR_destruct_r) q4acR_destruct_bufchan_d <= q4acR_destruct_d;
  Pointer_QTree_Bool_t q4acR_destruct_bufchan_buf;
  assign q4acR_destruct_bufchan_r = (! q4acR_destruct_bufchan_buf[0]);
  assign q4acR_1_argbuf_d = (q4acR_destruct_bufchan_buf[0] ? q4acR_destruct_bufchan_buf :
                             q4acR_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acR_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acR_1_argbuf_r && q4acR_destruct_bufchan_buf[0]))
        q4acR_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acR_1_argbuf_r) && (! q4acR_destruct_bufchan_buf[0])))
        q4acR_destruct_bufchan_buf <= q4acR_destruct_bufchan_d;
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf,CTkron_kron_Bool_Bool_Bool) > (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r = ((! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d <= {83'd0,
                                                                            1'd0};
    else
      if (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r)
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d <= readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r = (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d = (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf :
                                                                          readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= {83'd0,
                                                                              1'd0};
    else
      if ((readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r && readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= {83'd0,
                                                                                1'd0};
      else if (((! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r) && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CTkron_kron_Bool_Bool_Bool) : (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb,CTkron_kron_Bool_Bool_Bool) > [(lizzieLet20_1,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet20_2,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet20_3,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet20_4,CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet20_1_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet20_2_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet20_3_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet20_4_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done = (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet20_4_d[0],
                                                                                                                                                     lizzieLet20_3_d[0],
                                                                                                                                                     lizzieLet20_2_d[0],
                                                                                                                                                     lizzieLet20_1_d[0]} & {lizzieLet20_4_r,
                                                                                                                                                                            lizzieLet20_3_r,
                                                                                                                                                                            lizzieLet20_2_r,
                                                                                                                                                                            lizzieLet20_1_r}));
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r = (& readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                                              readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_mask_Bool) : (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf,CTmain_mask_Bool) > (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb,CTmain_mask_Bool) */
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r = ((! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d <= {115'd0,
                                                                    1'd0};
    else
      if (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r)
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d = (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf :
                                                                  readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                      1'd0};
    else
      if ((readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r && readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                        1'd0};
      else if (((! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CTmain_mask_Bool) : (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb,CTmain_mask_Bool) > [(lizzieLet25_1,CTmain_mask_Bool),
                                                                                                       (lizzieLet25_2,CTmain_mask_Bool),
                                                                                                       (lizzieLet25_3,CTmain_mask_Bool),
                                                                                                       (lizzieLet25_4,CTmain_mask_Bool)] */
  logic [3:0] readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet25_1_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet25_2_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet25_3_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet25_4_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done = (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet25_4_d[0],
                                                                                                                                     lizzieLet25_3_d[0],
                                                                                                                                     lizzieLet25_2_d[0],
                                                                                                                                     lizzieLet25_1_d[0]} & {lizzieLet25_4_r,
                                                                                                                                                            lizzieLet25_3_r,
                                                                                                                                                            lizzieLet25_2_r,
                                                                                                                                                            lizzieLet25_1_r}));
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                                      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf,CTmap''_map''_Bool_Bool_Bool) > (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d  <= {68'd0,
                                                                                  1'd0};
    else
      if (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r )
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  :
                                                                                \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {68'd0,
                                                                                    1'd0};
    else
      if ((\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {68'd0,
                                                                                      1'd0};
      else if (((! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmap''_map''_Bool_Bool_Bool) : (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb,CTmap''_map''_Bool_Bool_Bool) > [(lizzieLet30_1,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet30_2,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet30_3,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet30_4,CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet30_1_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet30_2_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet30_3_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet30_4_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet30_4_d[0],
                                                                                                                                                                 lizzieLet30_3_d[0],
                                                                                                                                                                 lizzieLet30_2_d[0],
                                                                                                                                                                 lizzieLet30_1_d[0]} & {lizzieLet30_4_r,
                                                                                                                                                                                        lizzieLet30_3_r,
                                                                                                                                                                                        lizzieLet30_2_r,
                                                                                                                                                                                        lizzieLet30_1_r}));
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                                    \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreemskacj_1_argbuf,MaskQTree) > (readPointer_MaskQTreemskacj_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreemskacj_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreemskacj_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreemskacj_1_argbuf_r = ((! readPointer_MaskQTreemskacj_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreemskacj_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacj_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreemskacj_1_argbuf_r)
        readPointer_MaskQTreemskacj_1_argbuf_bufchan_d <= readPointer_MaskQTreemskacj_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreemskacj_1_argbuf_bufchan_r = (! readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreemskacj_1_argbuf_rwb_d = (readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf :
                                                       readPointer_MaskQTreemskacj_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreemskacj_1_argbuf_rwb_r && readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreemskacj_1_argbuf_rwb_r) && (! readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreemskacj_1_argbuf_bufchan_buf <= readPointer_MaskQTreemskacj_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreemskacj_1_argbuf_rwb,MaskQTree) > [(lizzieLet4_1,MaskQTree),
                                                                              (lizzieLet4_2,MaskQTree),
                                                                              (lizzieLet4_3,MaskQTree),
                                                                              (lizzieLet4_4,MaskQTree),
                                                                              (lizzieLet4_5,MaskQTree),
                                                                              (lizzieLet4_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreemskacj_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet4_5_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet4_6_d = {readPointer_MaskQTreemskacj_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreemskacj_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreemskacj_1_argbuf_rwb_done = (readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted | ({lizzieLet4_6_d[0],
                                                                                                               lizzieLet4_5_d[0],
                                                                                                               lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_6_r,
                                                                                                                                     lizzieLet4_5_r,
                                                                                                                                     lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_MaskQTreemskacj_1_argbuf_rwb_r = (& readPointer_MaskQTreemskacj_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreemskacj_1_argbuf_rwb_emitted <= (readPointer_MaskQTreemskacj_1_argbuf_rwb_r ? 6'd0 :
                                                           readPointer_MaskQTreemskacj_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm1acL_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm1acL_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm1acL_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm1acL_1_argbuf_r = ((! readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm1acL_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm1acL_1_argbuf_r)
        readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d <= readPointer_QTree_Boolm1acL_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm1acL_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm1acL_1_argbuf_rwb_d = (readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm1acL_1_argbuf_rwb_r && readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm1acL_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm1acL_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm1acL_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolm1acL_1_argbuf_rwb,QTree_Bool) > [(lizzieLet0_1,QTree_Bool),
                                                                                (lizzieLet0_2,QTree_Bool),
                                                                                (lizzieLet0_3,QTree_Bool),
                                                                                (lizzieLet0_4,QTree_Bool),
                                                                                (lizzieLet0_5,QTree_Bool),
                                                                                (lizzieLet0_6,QTree_Bool),
                                                                                (lizzieLet0_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Boolm1acL_1_argbuf_rwb_done;
  assign lizzieLet0_1_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet0_2_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet0_3_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet0_4_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet0_5_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet0_6_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet0_7_d = {readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1acL_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Boolm1acL_1_argbuf_rwb_done = (readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted | ({lizzieLet0_7_d[0],
                                                                                                               lizzieLet0_6_d[0],
                                                                                                               lizzieLet0_5_d[0],
                                                                                                               lizzieLet0_4_d[0],
                                                                                                               lizzieLet0_3_d[0],
                                                                                                               lizzieLet0_2_d[0],
                                                                                                               lizzieLet0_1_d[0]} & {lizzieLet0_7_r,
                                                                                                                                     lizzieLet0_6_r,
                                                                                                                                     lizzieLet0_5_r,
                                                                                                                                     lizzieLet0_4_r,
                                                                                                                                     lizzieLet0_3_r,
                                                                                                                                     lizzieLet0_2_r,
                                                                                                                                     lizzieLet0_1_r}));
  assign readPointer_QTree_Boolm1acL_1_argbuf_rwb_r = (& readPointer_QTree_Boolm1acL_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Boolm1acL_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolm1acL_1_argbuf_rwb_r ? 7'd0 :
                                                           readPointer_QTree_Boolm1acL_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_BoolmacD_1_argbuf,QTree_Bool) > (readPointer_QTree_BoolmacD_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_BoolmacD_1_argbuf_bufchan_d;
  logic readPointer_QTree_BoolmacD_1_argbuf_bufchan_r;
  assign readPointer_QTree_BoolmacD_1_argbuf_r = ((! readPointer_QTree_BoolmacD_1_argbuf_bufchan_d[0]) || readPointer_QTree_BoolmacD_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacD_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_BoolmacD_1_argbuf_r)
        readPointer_QTree_BoolmacD_1_argbuf_bufchan_d <= readPointer_QTree_BoolmacD_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf;
  assign readPointer_QTree_BoolmacD_1_argbuf_bufchan_r = (! readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_BoolmacD_1_argbuf_rwb_d = (readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf[0] ? readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_BoolmacD_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_BoolmacD_1_argbuf_rwb_r && readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_BoolmacD_1_argbuf_rwb_r) && (! readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_BoolmacD_1_argbuf_bufchan_buf <= readPointer_QTree_BoolmacD_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_BoolmacD_1_argbuf_rwb,QTree_Bool) > [(lizzieLet11_1_1,QTree_Bool),
                                                                               (lizzieLet11_1_2,QTree_Bool),
                                                                               (lizzieLet11_1_3,QTree_Bool),
                                                                               (lizzieLet11_1_4,QTree_Bool),
                                                                               (lizzieLet11_1_5,QTree_Bool),
                                                                               (lizzieLet11_1_6,QTree_Bool),
                                                                               (lizzieLet11_1_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_BoolmacD_1_argbuf_rwb_done;
  assign lizzieLet11_1_1_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet11_1_2_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet11_1_3_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet11_1_4_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet11_1_5_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet11_1_6_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet11_1_7_d = {readPointer_QTree_BoolmacD_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_BoolmacD_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_BoolmacD_1_argbuf_rwb_done = (readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted | ({lizzieLet11_1_7_d[0],
                                                                                                             lizzieLet11_1_6_d[0],
                                                                                                             lizzieLet11_1_5_d[0],
                                                                                                             lizzieLet11_1_4_d[0],
                                                                                                             lizzieLet11_1_3_d[0],
                                                                                                             lizzieLet11_1_2_d[0],
                                                                                                             lizzieLet11_1_1_d[0]} & {lizzieLet11_1_7_r,
                                                                                                                                      lizzieLet11_1_6_r,
                                                                                                                                      lizzieLet11_1_5_r,
                                                                                                                                      lizzieLet11_1_4_r,
                                                                                                                                      lizzieLet11_1_3_r,
                                                                                                                                      lizzieLet11_1_2_r,
                                                                                                                                      lizzieLet11_1_1_r}));
  assign readPointer_QTree_BoolmacD_1_argbuf_rwb_r = (& readPointer_QTree_BoolmacD_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_BoolmacD_1_argbuf_rwb_emitted <= (readPointer_QTree_BoolmacD_1_argbuf_rwb_r ? 7'd0 :
                                                          readPointer_QTree_BoolmacD_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolmaci_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolmaci_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolmaci_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolmaci_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolmaci_1_argbuf_r = ((! readPointer_QTree_Boolmaci_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolmaci_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolmaci_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolmaci_1_argbuf_r)
        readPointer_QTree_Boolmaci_1_argbuf_bufchan_d <= readPointer_QTree_Boolmaci_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolmaci_1_argbuf_bufchan_r = (! readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolmaci_1_argbuf_rwb_d = (readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Boolmaci_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolmaci_1_argbuf_rwb_r && readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolmaci_1_argbuf_rwb_r) && (! readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolmaci_1_argbuf_bufchan_buf <= readPointer_QTree_Boolmaci_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (sc_0_10_destruct,Pointer_CTmain_mask_Bool) > (sc_0_10_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  Pointer_CTmain_mask_Bool_t sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (sc_0_14_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sc_0_14_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (sc_0_6_destruct,Pointer_CTkron_kron_Bool_Bool_Bool) > (sc_0_6_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (scfarg_0_1_goMux_mux,Pointer_CTmain_mask_Bool) > (scfarg_0_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (scfarg_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) > (scfarg_0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (scfarg_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) > (scfarg_0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1acp_3_destruct,Pointer_QTree_Bool) > (t1acp_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1acp_3_destruct_bufchan_d;
  logic t1acp_3_destruct_bufchan_r;
  assign t1acp_3_destruct_r = ((! t1acp_3_destruct_bufchan_d[0]) || t1acp_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1acp_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1acp_3_destruct_r)
        t1acp_3_destruct_bufchan_d <= t1acp_3_destruct_d;
  Pointer_QTree_Bool_t t1acp_3_destruct_bufchan_buf;
  assign t1acp_3_destruct_bufchan_r = (! t1acp_3_destruct_bufchan_buf[0]);
  assign t1acp_3_1_argbuf_d = (t1acp_3_destruct_bufchan_buf[0] ? t1acp_3_destruct_bufchan_buf :
                               t1acp_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1acp_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1acp_3_1_argbuf_r && t1acp_3_destruct_bufchan_buf[0]))
        t1acp_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1acp_3_1_argbuf_r) && (! t1acp_3_destruct_bufchan_buf[0])))
        t1acp_3_destruct_bufchan_buf <= t1acp_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2acq_2_destruct,Pointer_QTree_Bool) > (t2acq_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2acq_2_destruct_bufchan_d;
  logic t2acq_2_destruct_bufchan_r;
  assign t2acq_2_destruct_r = ((! t2acq_2_destruct_bufchan_d[0]) || t2acq_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2acq_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2acq_2_destruct_r)
        t2acq_2_destruct_bufchan_d <= t2acq_2_destruct_d;
  Pointer_QTree_Bool_t t2acq_2_destruct_bufchan_buf;
  assign t2acq_2_destruct_bufchan_r = (! t2acq_2_destruct_bufchan_buf[0]);
  assign t2acq_2_1_argbuf_d = (t2acq_2_destruct_bufchan_buf[0] ? t2acq_2_destruct_bufchan_buf :
                               t2acq_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2acq_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2acq_2_1_argbuf_r && t2acq_2_destruct_bufchan_buf[0]))
        t2acq_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2acq_2_1_argbuf_r) && (! t2acq_2_destruct_bufchan_buf[0])))
        t2acq_2_destruct_bufchan_buf <= t2acq_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3acr_1_destruct,Pointer_QTree_Bool) > (t3acr_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3acr_1_destruct_bufchan_d;
  logic t3acr_1_destruct_bufchan_r;
  assign t3acr_1_destruct_r = ((! t3acr_1_destruct_bufchan_d[0]) || t3acr_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3acr_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3acr_1_destruct_r)
        t3acr_1_destruct_bufchan_d <= t3acr_1_destruct_d;
  Pointer_QTree_Bool_t t3acr_1_destruct_bufchan_buf;
  assign t3acr_1_destruct_bufchan_r = (! t3acr_1_destruct_bufchan_buf[0]);
  assign t3acr_1_1_argbuf_d = (t3acr_1_destruct_bufchan_buf[0] ? t3acr_1_destruct_bufchan_buf :
                               t3acr_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3acr_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3acr_1_1_argbuf_r && t3acr_1_destruct_bufchan_buf[0]))
        t3acr_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3acr_1_1_argbuf_r) && (! t3acr_1_destruct_bufchan_buf[0])))
        t3acr_1_destruct_bufchan_buf <= t3acr_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4acs_destruct,Pointer_QTree_Bool) > (t4acs_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4acs_destruct_bufchan_d;
  logic t4acs_destruct_bufchan_r;
  assign t4acs_destruct_r = ((! t4acs_destruct_bufchan_d[0]) || t4acs_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4acs_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4acs_destruct_r) t4acs_destruct_bufchan_d <= t4acs_destruct_d;
  Pointer_QTree_Bool_t t4acs_destruct_bufchan_buf;
  assign t4acs_destruct_bufchan_r = (! t4acs_destruct_bufchan_buf[0]);
  assign t4acs_1_argbuf_d = (t4acs_destruct_bufchan_buf[0] ? t4acs_destruct_bufchan_buf :
                             t4acs_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4acs_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4acs_1_argbuf_r && t4acs_destruct_bufchan_buf[0]))
        t4acs_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4acs_1_argbuf_r) && (! t4acs_destruct_bufchan_buf[0])))
        t4acs_destruct_bufchan_buf <= t4acs_destruct_bufchan_d;
  
  /* buf (Ty MyBool) : (v'acC_2_2,MyBool) > (v'acC_2_2_argbuf,MyBool) */
  MyBool_t \v'acC_2_2_bufchan_d ;
  logic \v'acC_2_2_bufchan_r ;
  assign \v'acC_2_2_r  = ((! \v'acC_2_2_bufchan_d [0]) || \v'acC_2_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_2_2_bufchan_d  <= {1'd0, 1'd0};
    else if (\v'acC_2_2_r ) \v'acC_2_2_bufchan_d  <= \v'acC_2_2_d ;
  MyBool_t \v'acC_2_2_bufchan_buf ;
  assign \v'acC_2_2_bufchan_r  = (! \v'acC_2_2_bufchan_buf [0]);
  assign \v'acC_2_2_argbuf_d  = (\v'acC_2_2_bufchan_buf [0] ? \v'acC_2_2_bufchan_buf  :
                                 \v'acC_2_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_2_2_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'acC_2_2_argbuf_r  && \v'acC_2_2_bufchan_buf [0]))
        \v'acC_2_2_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'acC_2_2_argbuf_r ) && (! \v'acC_2_2_bufchan_buf [0])))
        \v'acC_2_2_bufchan_buf  <= \v'acC_2_2_bufchan_d ;
  
  /* fork (Ty MyBool) : (v'acC_2_destruct,MyBool) > [(v'acC_2_1,MyBool),
                                                (v'acC_2_2,MyBool)] */
  logic [1:0] \v'acC_2_destruct_emitted ;
  logic [1:0] \v'acC_2_destruct_done ;
  assign \v'acC_2_1_d  = {\v'acC_2_destruct_d [1:1],
                          (\v'acC_2_destruct_d [0] && (! \v'acC_2_destruct_emitted [0]))};
  assign \v'acC_2_2_d  = {\v'acC_2_destruct_d [1:1],
                          (\v'acC_2_destruct_d [0] && (! \v'acC_2_destruct_emitted [1]))};
  assign \v'acC_2_destruct_done  = (\v'acC_2_destruct_emitted  | ({\v'acC_2_2_d [0],
                                                                   \v'acC_2_1_d [0]} & {\v'acC_2_2_r ,
                                                                                        \v'acC_2_1_r }));
  assign \v'acC_2_destruct_r  = (& \v'acC_2_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_2_destruct_emitted  <= 2'd0;
    else
      \v'acC_2_destruct_emitted  <= (\v'acC_2_destruct_r  ? 2'd0 :
                                     \v'acC_2_destruct_done );
  
  /* buf (Ty MyBool) : (v'acC_3_2,MyBool) > (v'acC_3_2_argbuf,MyBool) */
  MyBool_t \v'acC_3_2_bufchan_d ;
  logic \v'acC_3_2_bufchan_r ;
  assign \v'acC_3_2_r  = ((! \v'acC_3_2_bufchan_d [0]) || \v'acC_3_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_3_2_bufchan_d  <= {1'd0, 1'd0};
    else if (\v'acC_3_2_r ) \v'acC_3_2_bufchan_d  <= \v'acC_3_2_d ;
  MyBool_t \v'acC_3_2_bufchan_buf ;
  assign \v'acC_3_2_bufchan_r  = (! \v'acC_3_2_bufchan_buf [0]);
  assign \v'acC_3_2_argbuf_d  = (\v'acC_3_2_bufchan_buf [0] ? \v'acC_3_2_bufchan_buf  :
                                 \v'acC_3_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_3_2_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'acC_3_2_argbuf_r  && \v'acC_3_2_bufchan_buf [0]))
        \v'acC_3_2_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'acC_3_2_argbuf_r ) && (! \v'acC_3_2_bufchan_buf [0])))
        \v'acC_3_2_bufchan_buf  <= \v'acC_3_2_bufchan_d ;
  
  /* fork (Ty MyBool) : (v'acC_3_destruct,MyBool) > [(v'acC_3_1,MyBool),
                                                (v'acC_3_2,MyBool)] */
  logic [1:0] \v'acC_3_destruct_emitted ;
  logic [1:0] \v'acC_3_destruct_done ;
  assign \v'acC_3_1_d  = {\v'acC_3_destruct_d [1:1],
                          (\v'acC_3_destruct_d [0] && (! \v'acC_3_destruct_emitted [0]))};
  assign \v'acC_3_2_d  = {\v'acC_3_destruct_d [1:1],
                          (\v'acC_3_destruct_d [0] && (! \v'acC_3_destruct_emitted [1]))};
  assign \v'acC_3_destruct_done  = (\v'acC_3_destruct_emitted  | ({\v'acC_3_2_d [0],
                                                                   \v'acC_3_1_d [0]} & {\v'acC_3_2_r ,
                                                                                        \v'acC_3_1_r }));
  assign \v'acC_3_destruct_r  = (& \v'acC_3_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_3_destruct_emitted  <= 2'd0;
    else
      \v'acC_3_destruct_emitted  <= (\v'acC_3_destruct_r  ? 2'd0 :
                                     \v'acC_3_destruct_done );
  
  /* buf (Ty MyBool) : (v'acC_4_destruct,MyBool) > (v'acC_4_1_argbuf,MyBool) */
  MyBool_t \v'acC_4_destruct_bufchan_d ;
  logic \v'acC_4_destruct_bufchan_r ;
  assign \v'acC_4_destruct_r  = ((! \v'acC_4_destruct_bufchan_d [0]) || \v'acC_4_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acC_4_destruct_bufchan_d  <= {1'd0, 1'd0};
    else
      if (\v'acC_4_destruct_r )
        \v'acC_4_destruct_bufchan_d  <= \v'acC_4_destruct_d ;
  MyBool_t \v'acC_4_destruct_bufchan_buf ;
  assign \v'acC_4_destruct_bufchan_r  = (! \v'acC_4_destruct_bufchan_buf [0]);
  assign \v'acC_4_1_argbuf_d  = (\v'acC_4_destruct_bufchan_buf [0] ? \v'acC_4_destruct_bufchan_buf  :
                                 \v'acC_4_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \v'acC_4_destruct_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'acC_4_1_argbuf_r  && \v'acC_4_destruct_bufchan_buf [0]))
        \v'acC_4_destruct_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'acC_4_1_argbuf_r ) && (! \v'acC_4_destruct_bufchan_buf [0])))
        \v'acC_4_destruct_bufchan_buf  <= \v'acC_4_destruct_bufchan_d ;
  
  /* buf (Ty MyBool) : (vacE_destruct,MyBool) > (vacE_1_argbuf,MyBool) */
  MyBool_t vacE_destruct_bufchan_d;
  logic vacE_destruct_bufchan_r;
  assign vacE_destruct_r = ((! vacE_destruct_bufchan_d[0]) || vacE_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacE_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (vacE_destruct_r) vacE_destruct_bufchan_d <= vacE_destruct_d;
  MyBool_t vacE_destruct_bufchan_buf;
  assign vacE_destruct_bufchan_r = (! vacE_destruct_bufchan_buf[0]);
  assign vacE_1_argbuf_d = (vacE_destruct_bufchan_buf[0] ? vacE_destruct_bufchan_buf :
                            vacE_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacE_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((vacE_1_argbuf_r && vacE_destruct_bufchan_buf[0]))
        vacE_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! vacE_1_argbuf_r) && (! vacE_destruct_bufchan_buf[0])))
        vacE_destruct_bufchan_buf <= vacE_destruct_bufchan_d;
  
  /* buf (Ty MyBool) : (vacN_destruct,MyBool) > (vacN_1_argbuf,MyBool) */
  MyBool_t vacN_destruct_bufchan_d;
  logic vacN_destruct_bufchan_r;
  assign vacN_destruct_r = ((! vacN_destruct_bufchan_d[0]) || vacN_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacN_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (vacN_destruct_r) vacN_destruct_bufchan_d <= vacN_destruct_d;
  MyBool_t vacN_destruct_bufchan_buf;
  assign vacN_destruct_bufchan_r = (! vacN_destruct_bufchan_buf[0]);
  assign vacN_1_argbuf_d = (vacN_destruct_bufchan_buf[0] ? vacN_destruct_bufchan_buf :
                            vacN_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacN_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((vacN_1_argbuf_r && vacN_destruct_bufchan_buf[0]))
        vacN_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! vacN_1_argbuf_r) && (! vacN_destruct_bufchan_buf[0])))
        vacN_destruct_bufchan_buf <= vacN_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet13_1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf :
                                     writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca2_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca1_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca0_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf :
                                                                     writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca3_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                           1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
    else
      if ((sca3_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                               1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet18_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet18_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet18_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet26_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet26_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet26_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca2_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet27_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet27_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet27_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca1_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet28_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet28_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet28_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca0_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet9_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet9_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet9_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca3_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca3_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet15_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet9_1_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet9_1_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet19_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca2_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet31_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca1_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet32_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet33_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_r = ((! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_1_argbuf_r)
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet12_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet12_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet12_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet12_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet13_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_argbuf_r = ((! writeQTree_BoollizzieLet13_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_argbuf_r)
        writeQTree_BoollizzieLet13_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet13_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet13_1_argbuf_rwb_d = (writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet13_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet13_1_argbuf_rwb_r && writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet13_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet13_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet13_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet13_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_r = ((! writeQTree_BoollizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_r)
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_d = (writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet14_1_argbuf_rwb_r && writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet14_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet16_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet16_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet16_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet16_1_argbuf_r = ((! writeQTree_BoollizzieLet16_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet16_1_argbuf_r)
        writeQTree_BoollizzieLet16_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet16_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet16_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet16_1_argbuf_rwb_d = (writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet16_1_argbuf_rwb_r && writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet16_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet16_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet16_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet16_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet16_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet16_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet1_1_argbuf_r = ((! writeQTree_BoollizzieLet1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet1_1_argbuf_r)
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet1_1_argbuf_rwb_r && writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet10_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet24_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet24_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet24_1_argbuf_r = ((! writeQTree_BoollizzieLet24_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet24_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet24_1_argbuf_r)
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet24_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet24_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_d = (writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet24_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet24_1_argbuf_rwb_r && writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet24_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet24_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet24_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet24_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet24_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet24_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet24_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet29_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet29_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet29_1_argbuf_r = ((! writeQTree_BoollizzieLet29_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet29_1_argbuf_r)
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet29_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet29_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_d = (writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet29_1_argbuf_rwb_r && writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet29_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet29_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet29_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet29_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet29_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_r = ((! writeQTree_BoollizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_r)
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_d = (writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet34_1_argbuf_rwb_r && writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet34_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_r = ((! writeQTree_BoollizzieLet3_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_r)
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_d = (writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet3_1_argbuf_rwb_r && writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet3_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet12_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_r = ((! writeQTree_BoollizzieLet5_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_r)
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_d = (writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet5_1_argbuf_rwb_r && writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet5_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_r = ((! writeQTree_BoollizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_r)
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_d = (writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet7_1_argbuf_rwb_r && writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet7_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet8_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet8_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet8_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet8_1_argbuf_r = ((! writeQTree_BoollizzieLet8_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet8_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet8_1_argbuf_r)
        writeQTree_BoollizzieLet8_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet8_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet8_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet8_1_argbuf_rwb_d = (writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet8_1_argbuf_rwb_r && writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet8_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet8_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet8_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet8_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet8_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet8_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty MyBool) : (xabY_1,MyBool) > (xabY_1_argbuf,MyBool) */
  MyBool_t xabY_1_bufchan_d;
  logic xabY_1_bufchan_r;
  assign xabY_1_r = ((! xabY_1_bufchan_d[0]) || xabY_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xabY_1_bufchan_d <= {1'd0, 1'd0};
    else if (xabY_1_r) xabY_1_bufchan_d <= xabY_1_d;
  MyBool_t xabY_1_bufchan_buf;
  assign xabY_1_bufchan_r = (! xabY_1_bufchan_buf[0]);
  assign xabY_1_argbuf_d = (xabY_1_bufchan_buf[0] ? xabY_1_bufchan_buf :
                            xabY_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xabY_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((xabY_1_argbuf_r && xabY_1_bufchan_buf[0]))
        xabY_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! xabY_1_argbuf_r) && (! xabY_1_bufchan_buf[0])))
        xabY_1_bufchan_buf <= xabY_1_bufchan_d;
endmodule