`timescale 1ns/1ns
import mMaskKron_package::*;

module mMaskKron(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1adl_0_d,
  output logic m1adl_0_r,
  input Pointer_QTree_Int_t m2adm_1_d,
  output logic m2adm_1_r,
  input Pointer_QTree_Int_t m3adn_2_d,
  output logic m3adn_2_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Int_t \es_7_1I#_dout ,
  input logic \es_7_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1adl_0, 16, 65536, Pointer_MaskQTree), (m2adm_1, 16, 65536, Pointer_QTree_Int), (m3adn_2, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (es_7_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTmain_mask_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
CTmap__027__027_map__027__027_Int_Int_Int 16 3 (0,[0]) (1,[16p,0,0,32,16p,16p,16p]) (2,[16p,16p,0,0,32,16p,16p]) (3,[16p,16p,16p,0,0,32,16p]) (4,[16p,16p,16p,16p])
CTkron_kron_Int_Int_Int 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,0,0,16p,16p]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz_Int 16 0 (0,[0,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int 16 0 (0,[0,0,0,16p,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int 16 0 (0,[0,16p,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap__027__027_map__027__027_Int_Int_Int 16 0 (0,[0,0,0,32,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,0,0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_MaskQTree 16 0 (0,[0,16p,16p])
TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int 16 0 (0,[0,0,0,32,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go_5_d;
  logic go_5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  Go_t go__11_d;
  logic go__11_r;
  Go_t go__12_d;
  logic go__12_r;
  Go_t go__13_d;
  logic go__13_r;
  \Word16#_t  initHP_CT$wnnz_Int_d;
  logic initHP_CT$wnnz_Int_r;
  \Word16#_t  incrHP_CT$wnnz_Int_d;
  logic incrHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_d;
  logic incrHP_mergeCT$wnnz_Int_r;
  Go_t incrHP_CT$wnnz_Int1_d;
  logic incrHP_CT$wnnz_Int1_r;
  Go_t incrHP_CT$wnnz_Int2_d;
  logic incrHP_CT$wnnz_Int2_r;
  \Word16#_t  addHP_CT$wnnz_Int_d;
  logic addHP_CT$wnnz_Int_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_d;
  logic mergeHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_buf_d;
  logic incrHP_mergeCT$wnnz_Int_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_buf_d;
  logic mergeHP_CT$wnnz_Int_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_Int_d;
  logic forkHP1_CT$wnnz_Int_r;
  \Word16#_t  forkHP1_CT$wnnz_In2_d;
  logic forkHP1_CT$wnnz_In2_r;
  \Word16#_t  forkHP1_CT$wnnz_In3_d;
  logic forkHP1_CT$wnnz_In3_r;
  C2_t memMergeChoice_CT$wnnz_Int_d;
  logic memMergeChoice_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_d;
  logic memMergeIn_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_d;
  logic memOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memReadOut_CT$wnnz_Int_d;
  logic memReadOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memWriteOut_CT$wnnz_Int_d;
  logic memWriteOut_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_dbuf_d;
  logic memMergeIn_CT$wnnz_Int_dbuf_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_rbuf_d;
  logic memMergeIn_CT$wnnz_Int_rbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_dbuf_d;
  logic memOut_CT$wnnz_Int_dbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_rbuf_d;
  logic memOut_CT$wnnz_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_Int_d;
  logic destructReadIn_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t dconReadIn_CT$wnnz_Int_d;
  logic dconReadIn_CT$wnnz_Int_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_Int_d;
  logic writeMerge_choice_CT$wnnz_Int_r;
  CT$wnnz_Int_t writeMerge_data_CT$wnnz_Int_d;
  logic writeMerge_data_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_r;
  MemIn_CT$wnnz_Int_t dconWriteIn_CT$wnnz_Int_d;
  logic dconWriteIn_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t dconPtr_CT$wnnz_Int_d;
  logic dconPtr_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_CT$wnnz_Int_t demuxWriteResult_CT$wnnz_Int_d;
  logic demuxWriteResult_CT$wnnz_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C4_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1acN_1_argbuf_d;
  logic readPointer_QTree_Intm1acN_1_argbuf_r;
  QTree_Int_t readPointer_QTree_IntmacF_1_argbuf_d;
  logic readPointer_QTree_IntmacF_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intmack_1_argbuf_d;
  logic readPointer_QTree_Intmack_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intwsxl_1_1_argbuf_d;
  logic readPointer_QTree_Intwsxl_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C14_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_d;
  logic writeQTree_IntlizzieLet14_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_d;
  logic writeQTree_IntlizzieLet44_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  initHP_CTmain_mask_Int_d;
  logic initHP_CTmain_mask_Int_r;
  \Word16#_t  incrHP_CTmain_mask_Int_d;
  logic incrHP_CTmain_mask_Int_r;
  Go_t incrHP_mergeCTmain_mask_Int_d;
  logic incrHP_mergeCTmain_mask_Int_r;
  Go_t incrHP_CTmain_mask_Int1_d;
  logic incrHP_CTmain_mask_Int1_r;
  Go_t incrHP_CTmain_mask_Int2_d;
  logic incrHP_CTmain_mask_Int2_r;
  \Word16#_t  addHP_CTmain_mask_Int_d;
  logic addHP_CTmain_mask_Int_r;
  \Word16#_t  mergeHP_CTmain_mask_Int_d;
  logic mergeHP_CTmain_mask_Int_r;
  Go_t incrHP_mergeCTmain_mask_Int_buf_d;
  logic incrHP_mergeCTmain_mask_Int_buf_r;
  \Word16#_t  mergeHP_CTmain_mask_Int_buf_d;
  logic mergeHP_CTmain_mask_Int_buf_r;
  \Word16#_t  forkHP1_CTmain_mask_Int_d;
  logic forkHP1_CTmain_mask_Int_r;
  \Word16#_t  forkHP1_CTmain_mask_In2_d;
  logic forkHP1_CTmain_mask_In2_r;
  \Word16#_t  forkHP1_CTmain_mask_In3_d;
  logic forkHP1_CTmain_mask_In3_r;
  C2_t memMergeChoice_CTmain_mask_Int_d;
  logic memMergeChoice_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_d;
  logic memMergeIn_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_d;
  logic memOut_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memReadOut_CTmain_mask_Int_d;
  logic memReadOut_CTmain_mask_Int_r;
  MemOut_CTmain_mask_Int_t memWriteOut_CTmain_mask_Int_d;
  logic memWriteOut_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_dbuf_d;
  logic memMergeIn_CTmain_mask_Int_dbuf_r;
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_rbuf_d;
  logic memMergeIn_CTmain_mask_Int_rbuf_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_dbuf_d;
  logic memOut_CTmain_mask_Int_dbuf_r;
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_rbuf_d;
  logic memOut_CTmain_mask_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTmain_mask_Int_d;
  logic destructReadIn_CTmain_mask_Int_r;
  MemIn_CTmain_mask_Int_t dconReadIn_CTmain_mask_Int_d;
  logic dconReadIn_CTmain_mask_Int_r;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTmain_mask_Int_d;
  logic writeMerge_choice_CTmain_mask_Int_r;
  CTmain_mask_Int_t writeMerge_data_CTmain_mask_Int_d;
  logic writeMerge_data_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet15_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet24_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet36_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet37_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_d;
  logic writeCTmain_mask_IntlizzieLet38_1_argbuf_r;
  MemIn_CTmain_mask_Int_t dconWriteIn_CTmain_mask_Int_d;
  logic dconWriteIn_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t dconPtr_CTmain_mask_Int_d;
  logic dconPtr_CTmain_mask_Int_r;
  Pointer_CTmain_mask_Int_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Pointer_CTmain_mask_Int_t demuxWriteResult_CTmain_mask_Int_d;
  logic demuxWriteResult_CTmain_mask_Int_r;
  \Word16#_t  \initHP_CTmap''_map''_Int_Int_Int_d ;
  logic \initHP_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \incrHP_CTmap''_map''_Int_Int_Int_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_CTmap''_map''_Int_Int_Int1_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int1_r ;
  Go_t \incrHP_CTmap''_map''_Int_Int_Int2_d ;
  logic \incrHP_CTmap''_map''_Int_Int_Int2_r ;
  \Word16#_t  \addHP_CTmap''_map''_Int_Int_Int_d ;
  logic \addHP_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_buf_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_buf_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_Int_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_In2_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_In2_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Int_Int_In3_d ;
  logic \forkHP1_CTmap''_map''_Int_Int_In3_r ;
  C2_t \memMergeChoice_CTmap''_map''_Int_Int_Int_d ;
  logic \memMergeChoice_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memReadOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memReadOut_CTmap''_map''_Int_Int_Int_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memWriteOut_CTmap''_map''_Int_Int_Int_d ;
  logic \memWriteOut_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_dbuf_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_dbuf_r ;
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_rbuf_d ;
  logic \memOut_CTmap''_map''_Int_Int_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmap''_map''_Int_Int_Int_d ;
  logic \destructReadIn_CTmap''_map''_Int_Int_Int_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \dconReadIn_CTmap''_map''_Int_Int_Int_d ;
  logic \dconReadIn_CTmap''_map''_Int_Int_Int_r ;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmap''_map''_Int_Int_Int_d ;
  logic \writeMerge_choice_CTmap''_map''_Int_Int_Int_r ;
  \CTmap''_map''_Int_Int_Int_t  \writeMerge_data_CTmap''_map''_Int_Int_Int_d ;
  logic \writeMerge_data_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_r ;
  \MemIn_CTmap''_map''_Int_Int_Int_t  \dconWriteIn_CTmap''_map''_Int_Int_Int_d ;
  logic \dconWriteIn_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \dconPtr_CTmap''_map''_Int_Int_Int_d ;
  logic \dconPtr_CTmap''_map''_Int_Int_Int_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \demuxWriteResult_CTmap''_map''_Int_Int_Int_d ;
  logic \demuxWriteResult_CTmap''_map''_Int_Int_Int_r ;
  \Word16#_t  initHP_CTkron_kron_Int_Int_Int_d;
  logic initHP_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  incrHP_CTkron_kron_Int_Int_Int_d;
  logic incrHP_CTkron_kron_Int_Int_Int_r;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_r;
  Go_t incrHP_CTkron_kron_Int_Int_Int1_d;
  logic incrHP_CTkron_kron_Int_Int_Int1_r;
  Go_t incrHP_CTkron_kron_Int_Int_Int2_d;
  logic incrHP_CTkron_kron_Int_Int_Int2_r;
  \Word16#_t  addHP_CTkron_kron_Int_Int_Int_d;
  logic addHP_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_r;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_buf_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_buf_r;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_buf_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_buf_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_Int_d;
  logic forkHP1_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_In2_d;
  logic forkHP1_CTkron_kron_Int_Int_In2_r;
  \Word16#_t  forkHP1_CTkron_kron_Int_Int_In3_d;
  logic forkHP1_CTkron_kron_Int_Int_In3_r;
  C2_t memMergeChoice_CTkron_kron_Int_Int_Int_d;
  logic memMergeChoice_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_d;
  logic memOut_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memReadOut_CTkron_kron_Int_Int_Int_d;
  logic memReadOut_CTkron_kron_Int_Int_Int_r;
  MemOut_CTkron_kron_Int_Int_Int_t memWriteOut_CTkron_kron_Int_Int_Int_d;
  logic memWriteOut_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r;
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d;
  logic memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_dbuf_d;
  logic memOut_CTkron_kron_Int_Int_Int_dbuf_r;
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_rbuf_d;
  logic memOut_CTkron_kron_Int_Int_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTkron_kron_Int_Int_Int_d;
  logic destructReadIn_CTkron_kron_Int_Int_Int_r;
  MemIn_CTkron_kron_Int_Int_Int_t dconReadIn_CTkron_kron_Int_Int_Int_d;
  logic dconReadIn_CTkron_kron_Int_Int_Int_r;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CTkron_kron_Int_Int_Int_d;
  logic writeMerge_choice_CTkron_kron_Int_Int_Int_r;
  CTkron_kron_Int_Int_Int_t writeMerge_data_CTkron_kron_Int_Int_Int_d;
  logic writeMerge_data_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r;
  MemIn_CTkron_kron_Int_Int_Int_t dconWriteIn_CTkron_kron_Int_Int_Int_d;
  logic dconWriteIn_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t dconPtr_CTkron_kron_Int_Int_Int_d;
  logic dconPtr_CTkron_kron_Int_Int_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Pointer_CTkron_kron_Int_Int_Int_t demuxWriteResult_CTkron_kron_Int_Int_Int_d;
  logic demuxWriteResult_CTkron_kron_Int_Int_Int_r;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreemskacl_1_argbuf_d;
  logic readPointer_MaskQTreemskacl_1_argbuf_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_r ;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Int_t wsxl_1_argbuf_d;
  logic wsxl_1_argbuf_r;
  Int_t \es_7_1I#_d ;
  logic \es_7_1I#_r ;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t es_0_2_1_d;
  logic es_0_2_1_r;
  MyBool_t es_0_2_2_d;
  logic es_0_2_2_r;
  MyBool_t es_0_2_3_d;
  logic es_0_2_3_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r;
  MyDTInt_Int_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t xac0_1_d;
  logic xac0_1_r;
  Int_t xac0_2_d;
  logic xac0_2_r;
  Int_t arg0_1Dcon_main1_d;
  logic arg0_1Dcon_main1_r;
  Int_t arg0_1Dcon_main1_1_d;
  logic arg0_1Dcon_main1_1_r;
  Int_t arg0_1Dcon_main1_2_d;
  logic arg0_1Dcon_main1_2_r;
  Int_t arg0_1Dcon_main1_3_d;
  logic arg0_1Dcon_main1_3_r;
  Int_t arg0_1Dcon_main1_4_d;
  logic arg0_1Dcon_main1_4_r;
  \Int#_t  xase_destruct_d;
  logic xase_destruct_r;
  Int_t \arg0_1Dcon_main1_1I#_d ;
  logic \arg0_1Dcon_main1_1I#_r ;
  Go_t \arg0_1Dcon_main1_3I#_d ;
  logic \arg0_1Dcon_main1_3I#_r ;
  Go_t \arg0_1Dcon_main1_3I#_1_d ;
  logic \arg0_1Dcon_main1_3I#_1_r ;
  Go_t \arg0_1Dcon_main1_3I#_2_d ;
  logic \arg0_1Dcon_main1_3I#_2_r ;
  Go_t \arg0_1Dcon_main1_3I#_3_d ;
  logic \arg0_1Dcon_main1_3I#_3_r ;
  Go_t \arg0_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_main1_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_main1_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1X1j_1_Eq_d;
  logic lizzieLet1_1wild1X1j_1_Eq_r;
  Go_t \arg0_1Dcon_main1_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_main1_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_main1_d;
  logic arg0_2Dcon_main1_r;
  Int_t \arg0_2_1Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_2_1Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_4_r ;
  \Int#_t  xa1m0_destruct_d;
  logic xa1m0_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_1I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_r ;
  \Int#_t  ya1m1_destruct_d;
  logic ya1m1_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d ;
  logic \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r ;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r;
  Pointer_QTree_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r;
  Go_t call_$wnnz_Int_initBufi_d;
  logic call_$wnnz_Int_initBufi_r;
  C5_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t call_$wnnz_Int_unlockFork1_d;
  logic call_$wnnz_Int_unlockFork1_r;
  Go_t call_$wnnz_Int_unlockFork2_d;
  logic call_$wnnz_Int_unlockFork2_r;
  Go_t call_$wnnz_Int_unlockFork3_d;
  logic call_$wnnz_Int_unlockFork3_r;
  Go_t call_$wnnz_Int_initBuf_d;
  logic call_$wnnz_Int_initBuf_r;
  Go_t call_$wnnz_Int_goMux1_d;
  logic call_$wnnz_Int_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_Int_goMux2_d;
  logic call_$wnnz_Int_goMux2_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_Int_goMux3_d;
  logic call_$wnnz_Int_goMux3_r;
  Go_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_r;
  MyDTInt_Bool_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_r;
  MyDTInt_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_r;
  Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r;
  Go_t call_kron_kron_Int_Int_Int_initBufi_d;
  logic call_kron_kron_Int_Int_Int_initBufi_r;
  C5_t go_9_goMux_choice_d;
  logic go_9_goMux_choice_r;
  Go_t go_9_goMux_data_d;
  logic go_9_goMux_data_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork1_d;
  logic call_kron_kron_Int_Int_Int_unlockFork1_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork2_d;
  logic call_kron_kron_Int_Int_Int_unlockFork2_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork3_d;
  logic call_kron_kron_Int_Int_Int_unlockFork3_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork4_d;
  logic call_kron_kron_Int_Int_Int_unlockFork4_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork5_d;
  logic call_kron_kron_Int_Int_Int_unlockFork5_r;
  Go_t call_kron_kron_Int_Int_Int_unlockFork6_d;
  logic call_kron_kron_Int_Int_Int_unlockFork6_r;
  Go_t call_kron_kron_Int_Int_Int_initBuf_d;
  logic call_kron_kron_Int_Int_Int_initBuf_r;
  Go_t call_kron_kron_Int_Int_Int_goMux1_d;
  logic call_kron_kron_Int_Int_Int_goMux1_r;
  MyDTInt_Bool_t call_kron_kron_Int_Int_Int_goMux2_d;
  logic call_kron_kron_Int_Int_Int_goMux2_r;
  MyDTInt_Int_Int_t call_kron_kron_Int_Int_Int_goMux3_d;
  logic call_kron_kron_Int_Int_Int_goMux3_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_Int_goMux4_d;
  logic call_kron_kron_Int_Int_Int_goMux4_r;
  Pointer_QTree_Int_t call_kron_kron_Int_Int_Int_goMux5_d;
  logic call_kron_kron_Int_Int_Int_goMux5_r;
  Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_Int_goMux6_d;
  logic call_kron_kron_Int_Int_Int_goMux6_r;
  Go_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_r;
  Pointer_QTree_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_r;
  Pointer_MaskQTree_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_r;
  Pointer_CTmain_mask_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r;
  Go_t call_main_mask_Int_initBufi_d;
  logic call_main_mask_Int_initBufi_r;
  C5_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t call_main_mask_Int_unlockFork1_d;
  logic call_main_mask_Int_unlockFork1_r;
  Go_t call_main_mask_Int_unlockFork2_d;
  logic call_main_mask_Int_unlockFork2_r;
  Go_t call_main_mask_Int_unlockFork3_d;
  logic call_main_mask_Int_unlockFork3_r;
  Go_t call_main_mask_Int_unlockFork4_d;
  logic call_main_mask_Int_unlockFork4_r;
  Go_t call_main_mask_Int_initBuf_d;
  logic call_main_mask_Int_initBuf_r;
  Go_t call_main_mask_Int_goMux1_d;
  logic call_main_mask_Int_goMux1_r;
  Pointer_QTree_Int_t call_main_mask_Int_goMux2_d;
  logic call_main_mask_Int_goMux2_r;
  Pointer_MaskQTree_t call_main_mask_Int_goMux3_d;
  logic call_main_mask_Int_goMux3_r;
  Pointer_CTmain_mask_Int_t call_main_mask_Int_goMux4_d;
  logic call_main_mask_Int_goMux4_r;
  Go_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_r ;
  MyDTInt_Bool_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_r ;
  MyDTInt_Int_Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_r ;
  Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_r ;
  Pointer_QTree_Int_t \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r ;
  Go_t \call_map''_map''_Int_Int_Int_initBufi_d ;
  logic \call_map''_map''_Int_Int_Int_initBufi_r ;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork1_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork1_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork2_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork2_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork3_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork3_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork4_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork4_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork5_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork5_r ;
  Go_t \call_map''_map''_Int_Int_Int_unlockFork6_d ;
  logic \call_map''_map''_Int_Int_Int_unlockFork6_r ;
  Go_t \call_map''_map''_Int_Int_Int_initBuf_d ;
  logic \call_map''_map''_Int_Int_Int_initBuf_r ;
  Go_t \call_map''_map''_Int_Int_Int_goMux1_d ;
  logic \call_map''_map''_Int_Int_Int_goMux1_r ;
  MyDTInt_Bool_t \call_map''_map''_Int_Int_Int_goMux2_d ;
  logic \call_map''_map''_Int_Int_Int_goMux2_r ;
  MyDTInt_Int_Int_t \call_map''_map''_Int_Int_Int_goMux3_d ;
  logic \call_map''_map''_Int_Int_Int_goMux3_r ;
  Int_t \call_map''_map''_Int_Int_Int_goMux4_d ;
  logic \call_map''_map''_Int_Int_Int_goMux4_r ;
  Pointer_QTree_Int_t \call_map''_map''_Int_Int_Int_goMux5_d ;
  logic \call_map''_map''_Int_Int_Int_goMux5_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_Int_goMux6_d ;
  logic \call_map''_map''_Int_Int_Int_goMux6_r ;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Go_t es_0_2_1MyFalse_d;
  logic es_0_2_1MyFalse_r;
  Go_t es_0_2_1MyTrue_d;
  logic es_0_2_1MyTrue_r;
  Go_t es_0_2_1MyFalse_1_argbuf_d;
  logic es_0_2_1MyFalse_1_argbuf_r;
  Go_t es_0_2_1MyTrue_1_d;
  logic es_0_2_1MyTrue_1_r;
  Go_t es_0_2_1MyTrue_2_d;
  logic es_0_2_1MyTrue_2_r;
  QTree_Int_t es_0_2_1MyTrue_1QNone_Int_d;
  logic es_0_2_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Go_t es_0_2_1MyTrue_2_argbuf_d;
  logic es_0_2_1MyTrue_2_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyFalse_d;
  logic es_0_2_2MyFalse_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyTrue_d;
  logic es_0_2_2MyTrue_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyFalse_1_argbuf_d;
  logic es_0_2_2MyFalse_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyTrue_1_argbuf_d;
  logic es_0_2_2MyTrue_1_argbuf_r;
  Int_t es_0_2_3MyFalse_d;
  logic es_0_2_3MyFalse_r;
  Int_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  QTree_Int_t es_0_2_3MyFalse_1QVal_Int_d;
  logic es_0_2_3MyFalse_1QVal_Int_r;
  QTree_Int_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  \Int#_t  es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_d;
  logic es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_r;
  MyDTInt_Int_Int_t gacD_2_2_argbuf_d;
  logic gacD_2_2_argbuf_r;
  MyDTInt_Int_Int_t gacD_2_1_d;
  logic gacD_2_1_r;
  MyDTInt_Int_Int_t gacD_2_2_d;
  logic gacD_2_2_r;
  MyDTInt_Int_Int_t gacD_3_2_argbuf_d;
  logic gacD_3_2_argbuf_r;
  MyDTInt_Int_Int_t gacD_3_1_d;
  logic gacD_3_1_r;
  MyDTInt_Int_Int_t gacD_3_2_d;
  logic gacD_3_2_r;
  MyDTInt_Int_Int_t gacD_4_1_argbuf_d;
  logic gacD_4_1_argbuf_r;
  MyDTInt_Int_Int_t gacM_2_2_argbuf_d;
  logic gacM_2_2_argbuf_r;
  MyDTInt_Int_Int_t gacM_2_1_d;
  logic gacM_2_1_r;
  MyDTInt_Int_Int_t gacM_2_2_d;
  logic gacM_2_2_r;
  MyDTInt_Int_Int_t gacM_3_2_argbuf_d;
  logic gacM_3_2_argbuf_r;
  MyDTInt_Int_Int_t gacM_3_1_d;
  logic gacM_3_1_r;
  MyDTInt_Int_Int_t gacM_3_2_d;
  logic gacM_3_2_r;
  MyDTInt_Int_Int_t gacM_4_1_argbuf_d;
  logic gacM_4_1_argbuf_r;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$ctimes_d ;
  logic \go_1Dcon_$fNumInt_$ctimes_r ;
  C5_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C5_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  C5_t go_10_goMux_choice_3_d;
  logic go_10_goMux_choice_3_r;
  Pointer_QTree_Int_t mack_goMux_mux_d;
  logic mack_goMux_mux_r;
  Pointer_MaskQTree_t mskacl_goMux_mux_d;
  logic mskacl_goMux_mux_r;
  Pointer_CTmain_mask_Int_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  C5_t go_11_goMux_choice_3_d;
  logic go_11_goMux_choice_3_r;
  C5_t go_11_goMux_choice_4_d;
  logic go_11_goMux_choice_4_r;
  C5_t go_11_goMux_choice_5_d;
  logic go_11_goMux_choice_5_r;
  MyDTInt_Bool_t isZacC_goMux_mux_d;
  logic isZacC_goMux_mux_r;
  MyDTInt_Int_Int_t gacD_goMux_mux_d;
  logic gacD_goMux_mux_r;
  Int_t \v'acE_goMux_mux_d ;
  logic \v'acE_goMux_mux_r ;
  Pointer_QTree_Int_t macF_goMux_mux_d;
  logic macF_goMux_mux_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_3_goMux_mux_d;
  logic sc_0_3_goMux_mux_r;
  CTkron_kron_Int_Int_Int_t go_12_1Lkron_kron_Int_Int_Intsbos_d;
  logic go_12_1Lkron_kron_Int_Int_Intsbos_r;
  CTkron_kron_Int_Int_Int_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t go_12_2_argbuf_d;
  logic go_12_2_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_t call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d;
  logic call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r;
  CTmain_mask_Int_t go_13_1Lmain_mask_Intsbos_d;
  logic go_13_1Lmain_mask_Intsbos_r;
  CTmain_mask_Int_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Go_t go_13_2_argbuf_d;
  logic go_13_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_t call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d;
  logic call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r;
  \CTmap''_map''_Int_Int_Int_t  \go_14_1Lmap''_map''_Int_Int_Intsbos_d ;
  logic \go_14_1Lmap''_map''_Int_Int_Intsbos_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Go_t go_14_2_argbuf_d;
  logic go_14_2_argbuf_r;
  \TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_t  \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d ;
  logic \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r ;
  C4_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C4_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C4_t go_16_goMux_choice_1_d;
  logic go_16_goMux_choice_1_r;
  C4_t go_16_goMux_choice_2_d;
  logic go_16_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C6_t go_17_goMux_choice_1_d;
  logic go_17_goMux_choice_1_r;
  C6_t go_17_goMux_choice_2_d;
  logic go_17_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  C5_t go_18_goMux_choice_1_d;
  logic go_18_goMux_choice_1_r;
  C5_t go_18_goMux_choice_2_d;
  logic go_18_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_3_goMux_mux_d;
  logic srtarg_0_3_goMux_mux_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_d;
  logic scfarg_0_3_goMux_mux_r;
  MyDTInt_Int_Int_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  MyDTInt_Bool_t go_2Dcon_main1_d;
  logic go_2Dcon_main1_r;
  MyDTInt_Bool_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r;
  Go_t go_4_argbuf_d;
  logic go_4_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r;
  Go_t go_5_argbuf_d;
  logic go_5_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_d;
  logic go_6_1L$wnnz_Intsbos_r;
  CT$wnnz_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r;
  C5_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C5_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  Pointer_QTree_Int_t wsxl_1_goMux_mux_d;
  logic wsxl_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_9_goMux_choice_1_d;
  logic go_9_goMux_choice_1_r;
  C5_t go_9_goMux_choice_2_d;
  logic go_9_goMux_choice_2_r;
  C5_t go_9_goMux_choice_3_d;
  logic go_9_goMux_choice_3_r;
  C5_t go_9_goMux_choice_4_d;
  logic go_9_goMux_choice_4_r;
  C5_t go_9_goMux_choice_5_d;
  logic go_9_goMux_choice_5_r;
  MyDTInt_Bool_t isZacL_goMux_mux_d;
  logic isZacL_goMux_mux_r;
  MyDTInt_Int_Int_t gacM_goMux_mux_d;
  logic gacM_goMux_mux_r;
  Pointer_QTree_Int_t m1acN_goMux_mux_d;
  logic m1acN_goMux_mux_r;
  Pointer_QTree_Int_t m2acO_goMux_mux_d;
  logic m2acO_goMux_mux_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  MyDTInt_Bool_t isZacC_2_2_argbuf_d;
  logic isZacC_2_2_argbuf_r;
  MyDTInt_Bool_t isZacC_2_1_d;
  logic isZacC_2_1_r;
  MyDTInt_Bool_t isZacC_2_2_d;
  logic isZacC_2_2_r;
  MyDTInt_Bool_t isZacC_3_2_argbuf_d;
  logic isZacC_3_2_argbuf_r;
  MyDTInt_Bool_t isZacC_3_1_d;
  logic isZacC_3_1_r;
  MyDTInt_Bool_t isZacC_3_2_d;
  logic isZacC_3_2_r;
  MyDTInt_Bool_t isZacC_4_1_argbuf_d;
  logic isZacC_4_1_argbuf_r;
  MyDTInt_Bool_t isZacL_2_2_argbuf_d;
  logic isZacL_2_2_argbuf_r;
  MyDTInt_Bool_t isZacL_2_1_d;
  logic isZacL_2_1_r;
  MyDTInt_Bool_t isZacL_2_2_d;
  logic isZacL_2_2_r;
  MyDTInt_Bool_t isZacL_3_2_argbuf_d;
  logic isZacL_3_2_argbuf_r;
  MyDTInt_Bool_t isZacL_3_1_d;
  logic isZacL_3_1_r;
  MyDTInt_Bool_t isZacL_3_2_d;
  logic isZacL_3_2_r;
  MyDTInt_Bool_t isZacL_4_1_argbuf_d;
  logic isZacL_4_1_argbuf_r;
  Go_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_r;
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_r;
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_r;
  MyDTInt_Int_Int_t gacM_1_1_argbuf_d;
  logic gacM_1_1_argbuf_r;
  Go_t go_12_1_d;
  logic go_12_1_r;
  Go_t go_12_2_d;
  logic go_12_2_r;
  MyDTInt_Bool_t isZacL_1_1_argbuf_d;
  logic isZacL_1_1_argbuf_r;
  Pointer_QTree_Int_t m1acN_1_1_argbuf_d;
  logic m1acN_1_1_argbuf_r;
  Pointer_QTree_Int_t m2acO_1_1_argbuf_d;
  logic m2acO_1_1_argbuf_r;
  Pointer_QTree_Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Pointer_MaskQTree_t q1acm_destruct_d;
  logic q1acm_destruct_r;
  Pointer_MaskQTree_t q2acn_destruct_d;
  logic q2acn_destruct_r;
  Pointer_MaskQTree_t q3aco_destruct_d;
  logic q3aco_destruct_r;
  Pointer_MaskQTree_t q4acp_destruct_d;
  logic q4acp_destruct_r;
  MaskQTree_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  MaskQTree_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  MaskQTree_t lizzieLet10_1_1MQNode_d;
  logic lizzieLet10_1_1MQNode_r;
  Go_t lizzieLet10_1_3MQNone_d;
  logic lizzieLet10_1_3MQNone_r;
  Go_t lizzieLet10_1_3MQVal_d;
  logic lizzieLet10_1_3MQVal_r;
  Go_t lizzieLet10_1_3MQNode_d;
  logic lizzieLet10_1_3MQNode_r;
  Go_t lizzieLet10_1_3MQNone_1_d;
  logic lizzieLet10_1_3MQNone_1_r;
  Go_t lizzieLet10_1_3MQNone_2_d;
  logic lizzieLet10_1_3MQNone_2_r;
  QTree_Int_t lizzieLet10_1_3MQNone_1QNone_Int_d;
  logic lizzieLet10_1_3MQNone_1QNone_Int_r;
  QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet10_1_3MQNone_2_argbuf_d;
  logic lizzieLet10_1_3MQNone_2_argbuf_r;
  C6_t go_17_goMux_choice_d;
  logic go_17_goMux_choice_r;
  Go_t go_17_goMux_data_d;
  logic go_17_goMux_data_r;
  Go_t lizzieLet10_1_3MQVal_1_argbuf_d;
  logic lizzieLet10_1_3MQVal_1_argbuf_r;
  QTree_Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  QTree_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  QTree_Int_t lizzieLet10_1_4MQNode_d;
  logic lizzieLet10_1_4MQNode_r;
  QTree_Int_t lizzieLet10_1_4MQNode_1_d;
  logic lizzieLet10_1_4MQNode_1_r;
  QTree_Int_t lizzieLet10_1_4MQNode_2_d;
  logic lizzieLet10_1_4MQNode_2_r;
  QTree_Int_t lizzieLet10_1_4MQNode_3_d;
  logic lizzieLet10_1_4MQNode_3_r;
  QTree_Int_t lizzieLet10_1_4MQNode_4_d;
  logic lizzieLet10_1_4MQNode_4_r;
  QTree_Int_t lizzieLet10_1_4MQNode_5_d;
  logic lizzieLet10_1_4MQNode_5_r;
  QTree_Int_t lizzieLet10_1_4MQNode_6_d;
  logic lizzieLet10_1_4MQNode_6_r;
  QTree_Int_t lizzieLet10_1_4MQNode_7_d;
  logic lizzieLet10_1_4MQNode_7_r;
  QTree_Int_t lizzieLet10_1_4MQNode_8_d;
  logic lizzieLet10_1_4MQNode_8_r;
  Pointer_QTree_Int_t t1acr_destruct_d;
  logic t1acr_destruct_r;
  Pointer_QTree_Int_t t2acs_destruct_d;
  logic t2acs_destruct_r;
  Pointer_QTree_Int_t t3act_destruct_d;
  logic t3act_destruct_r;
  Pointer_QTree_Int_t t4acu_destruct_d;
  logic t4acu_destruct_r;
  QTree_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  QTree_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  QTree_Int_t lizzieLet10_1_4MQNode_1QNode_Int_d;
  logic lizzieLet10_1_4MQNode_1QNode_Int_r;
  QTree_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_r;
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_r;
  Go_t lizzieLet10_1_4MQNode_3QNode_Int_d;
  logic lizzieLet10_1_4MQNode_3QNode_Int_r;
  Go_t lizzieLet10_1_4MQNode_3QError_Int_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_r;
  Go_t lizzieLet10_1_4MQNode_3QError_Int_1_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_1_r;
  Go_t lizzieLet10_1_4MQNode_3QError_Int_2_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_2_r;
  QTree_Int_t lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_d;
  logic lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_1_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_1_r;
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_2_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_2_r;
  QTree_Int_t lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_1_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_1_r;
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_2_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_2_r;
  QTree_Int_t lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet14_2_1_argbuf_d;
  logic lizzieLet14_2_1_argbuf_r;
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNone_Int_d;
  logic lizzieLet10_1_4MQNode_4QNone_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QVal_Int_d;
  logic lizzieLet10_1_4MQNode_4QVal_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNode_Int_d;
  logic lizzieLet10_1_4MQNode_4QNode_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QError_Int_d;
  logic lizzieLet10_1_4MQNode_4QError_Int_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_d;
  logic lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d;
  logic lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r;
  CTmain_mask_Int_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_d;
  logic lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_d;
  logic lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_r;
  Pointer_MaskQTree_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_MaskQTree_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_5QNode_Int_d;
  logic lizzieLet10_1_4MQNode_5QNode_Int_r;
  Pointer_MaskQTree_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Pointer_MaskQTree_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Pointer_MaskQTree_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_6QNode_Int_d;
  logic lizzieLet10_1_4MQNode_6QNode_Int_r;
  Pointer_MaskQTree_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_MaskQTree_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Pointer_MaskQTree_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_7QNode_Int_d;
  logic lizzieLet10_1_4MQNode_7QNode_Int_r;
  Pointer_MaskQTree_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  Pointer_MaskQTree_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  Pointer_MaskQTree_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_8QNode_Int_d;
  logic lizzieLet10_1_4MQNode_8QNode_Int_r;
  Pointer_MaskQTree_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_d;
  logic lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet10_1_5MQVal_d;
  logic lizzieLet10_1_5MQVal_r;
  Pointer_QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet10_1_5MQVal_1_argbuf_d;
  logic lizzieLet10_1_5MQVal_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQNone_d;
  logic lizzieLet10_1_6MQNone_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQVal_d;
  logic lizzieLet10_1_6MQVal_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQNode_d;
  logic lizzieLet10_1_6MQNode_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQNone_1_argbuf_d;
  logic lizzieLet10_1_6MQNone_1_argbuf_r;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQVal_1_argbuf_d;
  logic lizzieLet10_1_6MQVal_1_argbuf_r;
  Pointer_QTree_Int_t q1acH_destruct_d;
  logic q1acH_destruct_r;
  Pointer_QTree_Int_t q2acI_destruct_d;
  logic q2acI_destruct_r;
  Pointer_QTree_Int_t q3acJ_destruct_d;
  logic q3acJ_destruct_r;
  Pointer_QTree_Int_t q4acK_destruct_d;
  logic q4acK_destruct_r;
  Int_t vacG_destruct_d;
  logic vacG_destruct_r;
  QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  QTree_Int_t lizzieLet17_1QVal_Int_d;
  logic lizzieLet17_1QVal_Int_r;
  QTree_Int_t lizzieLet17_1QNode_Int_d;
  logic lizzieLet17_1QNode_Int_r;
  QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MyDTInt_Int_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_3QVal_Int_d;
  logic lizzieLet17_3QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_d;
  logic lizzieLet17_3QNode_Int_r;
  MyDTInt_Int_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_1_d;
  logic lizzieLet17_3QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_2_d;
  logic lizzieLet17_3QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_2_argbuf_d;
  logic lizzieLet17_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet17_3QVal_Int_1_argbuf_d;
  logic lizzieLet17_3QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  Go_t lizzieLet17_4QNone_Int_d;
  logic lizzieLet17_4QNone_Int_r;
  Go_t lizzieLet17_4QVal_Int_d;
  logic lizzieLet17_4QVal_Int_r;
  Go_t lizzieLet17_4QNode_Int_d;
  logic lizzieLet17_4QNode_Int_r;
  Go_t lizzieLet17_4QError_Int_d;
  logic lizzieLet17_4QError_Int_r;
  Go_t lizzieLet17_4QError_Int_1_d;
  logic lizzieLet17_4QError_Int_1_r;
  Go_t lizzieLet17_4QError_Int_2_d;
  logic lizzieLet17_4QError_Int_2_r;
  QTree_Int_t lizzieLet17_4QError_Int_1QError_Int_d;
  logic lizzieLet17_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t lizzieLet17_4QError_Int_2_argbuf_d;
  logic lizzieLet17_4QError_Int_2_argbuf_r;
  Go_t lizzieLet17_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet17_4QNone_Int_1_d;
  logic lizzieLet17_4QNone_Int_1_r;
  Go_t lizzieLet17_4QNone_Int_2_d;
  logic lizzieLet17_4QNone_Int_2_r;
  QTree_Int_t lizzieLet17_4QNone_Int_1QNone_Int_d;
  logic lizzieLet17_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet17_4QNone_Int_2_argbuf_d;
  logic lizzieLet17_4QNone_Int_2_argbuf_r;
  C5_t go_18_goMux_choice_d;
  logic go_18_goMux_choice_r;
  Go_t go_18_goMux_data_d;
  logic go_18_goMux_data_r;
  Go_t lizzieLet17_4QVal_Int_1_d;
  logic lizzieLet17_4QVal_Int_1_r;
  Go_t lizzieLet17_4QVal_Int_2_d;
  logic lizzieLet17_4QVal_Int_2_r;
  Go_t lizzieLet17_4QVal_Int_1_argbuf_d;
  logic lizzieLet17_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_d;
  logic lizzieLet17_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_r;
  MyDTInt_Bool_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QNone_Int_d;
  logic lizzieLet17_6QNone_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QVal_Int_d;
  logic lizzieLet17_6QVal_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QNode_Int_d;
  logic lizzieLet17_6QNode_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QError_Int_d;
  logic lizzieLet17_6QError_Int_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QError_Int_1_argbuf_d;
  logic lizzieLet17_6QError_Int_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QNone_Int_1_argbuf_d;
  logic lizzieLet17_6QNone_Int_1_argbuf_r;
  Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Int_t lizzieLet17_7QVal_Int_d;
  logic lizzieLet17_7QVal_Int_r;
  Int_t lizzieLet17_7QNode_Int_d;
  logic lizzieLet17_7QNode_Int_r;
  Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Int_t lizzieLet17_7QNode_Int_1_d;
  logic lizzieLet17_7QNode_Int_1_r;
  Int_t lizzieLet17_7QNode_Int_2_d;
  logic lizzieLet17_7QNode_Int_2_r;
  Int_t lizzieLet17_7QNode_Int_2_argbuf_d;
  logic lizzieLet17_7QNode_Int_2_argbuf_r;
  Int_t lizzieLet17_7QVal_Int_1_argbuf_d;
  logic lizzieLet17_7QVal_Int_1_argbuf_r;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  \Int#_t  wwsxo_4_destruct_d;
  logic wwsxo_4_destruct_r;
  \Int#_t  ww1XyC_2_destruct_d;
  logic ww1XyC_2_destruct_r;
  \Int#_t  ww2XyF_1_destruct_d;
  logic ww2XyF_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  \Int#_t  wwsxo_3_destruct_d;
  logic wwsxo_3_destruct_r;
  \Int#_t  ww1XyC_1_destruct_d;
  logic ww1XyC_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Int_t q4acY_3_destruct_d;
  logic q4acY_3_destruct_r;
  \Int#_t  wwsxo_2_destruct_d;
  logic wwsxo_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4acY_2_destruct_d;
  logic q4acY_2_destruct_r;
  Pointer_QTree_Int_t q3acX_2_destruct_d;
  logic q3acX_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4acY_1_destruct_d;
  logic q4acY_1_destruct_r;
  Pointer_QTree_Int_t q3acX_1_destruct_d;
  logic q3acX_1_destruct_r;
  Pointer_QTree_Int_t q2acW_1_destruct_d;
  logic q2acW_1_destruct_r;
  CT$wnnz_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  CT$wnnz_Int_t lizzieLet26_1Lcall_$wnnz_Int3_d;
  logic lizzieLet26_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet26_1Lcall_$wnnz_Int2_d;
  logic lizzieLet26_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet26_1Lcall_$wnnz_Int1_d;
  logic lizzieLet26_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet26_1Lcall_$wnnz_Int0_d;
  logic lizzieLet26_1Lcall_$wnnz_Int0_r;
  Go_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Go_t lizzieLet26_3Lcall_$wnnz_Int3_d;
  logic lizzieLet26_3Lcall_$wnnz_Int3_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int2_d;
  logic lizzieLet26_3Lcall_$wnnz_Int2_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int1_d;
  logic lizzieLet26_3Lcall_$wnnz_Int1_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int0_d;
  logic lizzieLet26_3Lcall_$wnnz_Int0_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_d;
  logic lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_d;
  logic lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_d;
  logic lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_r;
  Go_t lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_d;
  logic lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_r;
  \Int#_t  lizzieLet26_4L$wnnz_Intsbos_d;
  logic lizzieLet26_4L$wnnz_Intsbos_r;
  \Int#_t  lizzieLet26_4Lcall_$wnnz_Int3_d;
  logic lizzieLet26_4Lcall_$wnnz_Int3_r;
  \Int#_t  lizzieLet26_4Lcall_$wnnz_Int2_d;
  logic lizzieLet26_4Lcall_$wnnz_Int2_r;
  \Int#_t  lizzieLet26_4Lcall_$wnnz_Int1_d;
  logic lizzieLet26_4Lcall_$wnnz_Int1_r;
  \Int#_t  lizzieLet26_4Lcall_$wnnz_Int0_d;
  logic lizzieLet26_4Lcall_$wnnz_Int0_r;
  \Int#_t  lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_Int_goConst_d;
  logic call_$wnnz_Int_goConst_r;
  \Int#_t  \$wnnz_Int_resbuf_d ;
  logic \$wnnz_Int_resbuf_r ;
  CT$wnnz_Int_t lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_d;
  logic lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  Pointer_QTree_Int_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Int_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Int_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t es_2_destruct_d;
  logic es_2_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  MyDTInt_Bool_t isZacL_4_destruct_d;
  logic isZacL_4_destruct_r;
  MyDTInt_Int_Int_t gacM_4_destruct_d;
  logic gacM_4_destruct_r;
  Pointer_QTree_Int_t q1acQ_3_destruct_d;
  logic q1acQ_3_destruct_r;
  Pointer_QTree_Int_t m2acO_4_destruct_d;
  logic m2acO_4_destruct_r;
  Pointer_QTree_Int_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  MyDTInt_Bool_t isZacL_3_destruct_d;
  logic isZacL_3_destruct_r;
  MyDTInt_Int_Int_t gacM_3_destruct_d;
  logic gacM_3_destruct_r;
  Pointer_QTree_Int_t q1acQ_2_destruct_d;
  logic q1acQ_2_destruct_r;
  Pointer_QTree_Int_t m2acO_3_destruct_d;
  logic m2acO_3_destruct_r;
  Pointer_QTree_Int_t q2acR_2_destruct_d;
  logic q2acR_2_destruct_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  MyDTInt_Bool_t isZacL_2_destruct_d;
  logic isZacL_2_destruct_r;
  MyDTInt_Int_Int_t gacM_2_destruct_d;
  logic gacM_2_destruct_r;
  Pointer_QTree_Int_t q1acQ_1_destruct_d;
  logic q1acQ_1_destruct_r;
  Pointer_QTree_Int_t m2acO_2_destruct_d;
  logic m2acO_2_destruct_r;
  Pointer_QTree_Int_t q2acR_1_destruct_d;
  logic q2acR_1_destruct_r;
  Pointer_QTree_Int_t q3acS_1_destruct_d;
  logic q3acS_1_destruct_r;
  CTkron_kron_Int_Int_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_r;
  Go_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d;
  logic lizzieLet30_4Lkron_kron_Int_Int_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_r;
  Pointer_QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_r;
  Pointer_QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_r;
  Pointer_QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_r;
  QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_r;
  QTree_Int_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r;
  CTkron_kron_Int_Int_Int_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_kron_kron_Int_Int_Int_goConst_d;
  logic call_kron_kron_Int_Int_Int_goConst_r;
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_d;
  logic kron_kron_Int_Int_Int_resbuf_r;
  Pointer_QTree_Int_t es_1_2_destruct_d;
  logic es_1_2_destruct_r;
  Pointer_QTree_Int_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Int_t es_3_6_destruct_d;
  logic es_3_6_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_15_destruct_d;
  logic sc_0_15_destruct_r;
  Pointer_QTree_Int_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Int_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t t1acr_3_destruct_d;
  logic t1acr_3_destruct_r;
  Pointer_MaskQTree_t q1acm_3_destruct_d;
  logic q1acm_3_destruct_r;
  Pointer_QTree_Int_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t t1acr_2_destruct_d;
  logic t1acr_2_destruct_r;
  Pointer_MaskQTree_t q1acm_2_destruct_d;
  logic q1acm_2_destruct_r;
  Pointer_QTree_Int_t t2acs_2_destruct_d;
  logic t2acs_2_destruct_r;
  Pointer_MaskQTree_t q2acn_2_destruct_d;
  logic q2acn_2_destruct_r;
  Pointer_CTmain_mask_Int_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t t1acr_1_destruct_d;
  logic t1acr_1_destruct_r;
  Pointer_MaskQTree_t q1acm_1_destruct_d;
  logic q1acm_1_destruct_r;
  Pointer_QTree_Int_t t2acs_1_destruct_d;
  logic t2acs_1_destruct_r;
  Pointer_MaskQTree_t q2acn_1_destruct_d;
  logic q2acn_1_destruct_r;
  Pointer_QTree_Int_t t3act_1_destruct_d;
  logic t3act_1_destruct_r;
  Pointer_MaskQTree_t q3aco_1_destruct_d;
  logic q3aco_1_destruct_r;
  CTmain_mask_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  CTmain_mask_Int_t lizzieLet35_1Lcall_main_mask_Int3_d;
  logic lizzieLet35_1Lcall_main_mask_Int3_r;
  CTmain_mask_Int_t lizzieLet35_1Lcall_main_mask_Int2_d;
  logic lizzieLet35_1Lcall_main_mask_Int2_r;
  CTmain_mask_Int_t lizzieLet35_1Lcall_main_mask_Int1_d;
  logic lizzieLet35_1Lcall_main_mask_Int1_r;
  CTmain_mask_Int_t lizzieLet35_1Lcall_main_mask_Int0_d;
  logic lizzieLet35_1Lcall_main_mask_Int0_r;
  Go_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Go_t lizzieLet35_3Lcall_main_mask_Int3_d;
  logic lizzieLet35_3Lcall_main_mask_Int3_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int2_d;
  logic lizzieLet35_3Lcall_main_mask_Int2_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int1_d;
  logic lizzieLet35_3Lcall_main_mask_Int1_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int0_d;
  logic lizzieLet35_3Lcall_main_mask_Int0_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_d;
  logic lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_d;
  logic lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_d;
  logic lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_r;
  Go_t lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_d;
  logic lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet35_4Lmain_mask_Intsbos_d;
  logic lizzieLet35_4Lmain_mask_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet35_4Lcall_main_mask_Int3_d;
  logic lizzieLet35_4Lcall_main_mask_Int3_r;
  Pointer_QTree_Int_t lizzieLet35_4Lcall_main_mask_Int2_d;
  logic lizzieLet35_4Lcall_main_mask_Int2_r;
  Pointer_QTree_Int_t lizzieLet35_4Lcall_main_mask_Int1_d;
  logic lizzieLet35_4Lcall_main_mask_Int1_r;
  Pointer_QTree_Int_t lizzieLet35_4Lcall_main_mask_Int0_d;
  logic lizzieLet35_4Lcall_main_mask_Int0_r;
  QTree_Int_t lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_d;
  logic lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_r;
  QTree_Int_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_d;
  logic lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_r;
  CTmain_mask_Int_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_d;
  logic lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_r;
  CTmain_mask_Int_t lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_d;
  logic lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_r;
  CTmain_mask_Int_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_main_mask_Int_goConst_d;
  logic call_main_mask_Int_goConst_r;
  Pointer_QTree_Int_t main_mask_Int_resbuf_d;
  logic main_mask_Int_resbuf_r;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  Pointer_QTree_Int_t es_2_4_destruct_d;
  logic es_2_4_destruct_r;
  Pointer_QTree_Int_t es_3_8_destruct_d;
  logic es_3_8_destruct_r;
  Pointer_QTree_Int_t es_4_4_destruct_d;
  logic es_4_4_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_d;
  logic sc_0_19_destruct_r;
  Pointer_QTree_Int_t es_3_7_destruct_d;
  logic es_3_7_destruct_r;
  Pointer_QTree_Int_t es_4_3_destruct_d;
  logic es_4_3_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_18_destruct_d;
  logic sc_0_18_destruct_r;
  MyDTInt_Bool_t isZacC_4_destruct_d;
  logic isZacC_4_destruct_r;
  MyDTInt_Int_Int_t gacD_4_destruct_d;
  logic gacD_4_destruct_r;
  Int_t \v'acE_4_destruct_d ;
  logic \v'acE_4_destruct_r ;
  Pointer_QTree_Int_t q1acH_3_destruct_d;
  logic q1acH_3_destruct_r;
  Pointer_QTree_Int_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_17_destruct_d;
  logic sc_0_17_destruct_r;
  MyDTInt_Bool_t isZacC_3_destruct_d;
  logic isZacC_3_destruct_r;
  MyDTInt_Int_Int_t gacD_3_destruct_d;
  logic gacD_3_destruct_r;
  Int_t \v'acE_3_destruct_d ;
  logic \v'acE_3_destruct_r ;
  Pointer_QTree_Int_t q1acH_2_destruct_d;
  logic q1acH_2_destruct_r;
  Pointer_QTree_Int_t q2acI_2_destruct_d;
  logic q2acI_2_destruct_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_16_destruct_d;
  logic sc_0_16_destruct_r;
  MyDTInt_Bool_t isZacC_2_destruct_d;
  logic isZacC_2_destruct_r;
  MyDTInt_Int_Int_t gacD_2_destruct_d;
  logic gacD_2_destruct_r;
  Int_t \v'acE_2_destruct_d ;
  logic \v'acE_2_destruct_r ;
  Pointer_QTree_Int_t q1acH_1_destruct_d;
  logic q1acH_1_destruct_r;
  Pointer_QTree_Int_t q2acI_1_destruct_d;
  logic q2acI_1_destruct_r;
  Pointer_QTree_Int_t q3acJ_1_destruct_d;
  logic q3acJ_1_destruct_r;
  \CTmap''_map''_Int_Int_Int_t  _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_r ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_r ;
  Go_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d ;
  logic \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_r ;
  QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_r ;
  QTree_Int_t lizzieLet44_1_argbuf_d;
  logic lizzieLet44_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_map''_map''_Int_Int_Int_goConst_d ;
  logic \call_map''_map''_Int_Int_Int_goConst_r ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_d ;
  logic \map''_map''_Int_Int_Int_resbuf_r ;
  Pointer_QTree_Int_t q1acV_destruct_d;
  logic q1acV_destruct_r;
  Pointer_QTree_Int_t q2acW_destruct_d;
  logic q2acW_destruct_r;
  Pointer_QTree_Int_t q3acX_destruct_d;
  logic q3acX_destruct_r;
  Pointer_QTree_Int_t q4acY_destruct_d;
  logic q4acY_destruct_r;
  QTree_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  QTree_Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_d;
  logic lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t q1acQ_destruct_d;
  logic q1acQ_destruct_r;
  Pointer_QTree_Int_t q2acR_destruct_d;
  logic q2acR_destruct_r;
  Pointer_QTree_Int_t q3acS_destruct_d;
  logic q3acS_destruct_r;
  Pointer_QTree_Int_t q4acT_destruct_d;
  logic q4acT_destruct_r;
  Int_t vacP_destruct_d;
  logic vacP_destruct_r;
  QTree_Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  QTree_Int_t lizzieLet6_1QVal_Int_d;
  logic lizzieLet6_1QVal_Int_r;
  QTree_Int_t lizzieLet6_1QNode_Int_d;
  logic lizzieLet6_1QNode_Int_r;
  QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  MyDTInt_Int_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_d;
  logic lizzieLet6_3QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_d;
  logic lizzieLet6_3QNode_Int_r;
  MyDTInt_Int_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_1_d;
  logic lizzieLet6_3QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_d;
  logic lizzieLet6_3QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_argbuf_d;
  logic lizzieLet6_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_1_argbuf_d;
  logic lizzieLet6_3QVal_Int_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_d;
  logic lizzieLet6_4QNone_Int_r;
  Go_t lizzieLet6_4QVal_Int_d;
  logic lizzieLet6_4QVal_Int_r;
  Go_t lizzieLet6_4QNode_Int_d;
  logic lizzieLet6_4QNode_Int_r;
  Go_t lizzieLet6_4QError_Int_d;
  logic lizzieLet6_4QError_Int_r;
  Go_t lizzieLet6_4QError_Int_1_d;
  logic lizzieLet6_4QError_Int_1_r;
  Go_t lizzieLet6_4QError_Int_2_d;
  logic lizzieLet6_4QError_Int_2_r;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_d;
  logic lizzieLet6_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t lizzieLet6_4QError_Int_2_argbuf_d;
  logic lizzieLet6_4QError_Int_2_argbuf_r;
  Go_t lizzieLet6_4QNode_Int_1_argbuf_d;
  logic lizzieLet6_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_1_d;
  logic lizzieLet6_4QNone_Int_1_r;
  Go_t lizzieLet6_4QNone_Int_2_d;
  logic lizzieLet6_4QNone_Int_2_r;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_2_argbuf_d;
  logic lizzieLet6_4QNone_Int_2_argbuf_r;
  C4_t go_16_goMux_choice_d;
  logic go_16_goMux_choice_r;
  Go_t go_16_goMux_data_d;
  logic go_16_goMux_data_r;
  Go_t lizzieLet6_4QVal_Int_1_d;
  logic lizzieLet6_4QVal_Int_1_r;
  Go_t lizzieLet6_4QVal_Int_2_d;
  logic lizzieLet6_4QVal_Int_2_r;
  Go_t lizzieLet6_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r ;
  Go_t lizzieLet6_4QVal_Int_2_argbuf_d;
  logic lizzieLet6_4QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_r;
  MyDTInt_Bool_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_d;
  logic lizzieLet6_6QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_d;
  logic lizzieLet6_6QNode_Int_r;
  Pointer_QTree_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_1_d;
  logic lizzieLet6_6QNode_Int_1_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_d;
  logic lizzieLet6_6QNode_Int_2_r;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_argbuf_d;
  logic lizzieLet6_6QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_1_argbuf_d;
  logic lizzieLet6_6QVal_Int_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_d;
  logic lizzieLet6_7QNone_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_d;
  logic lizzieLet6_7QVal_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_d;
  logic lizzieLet6_7QNode_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_d;
  logic lizzieLet6_7QError_Int_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_1_argbuf_d;
  logic lizzieLet6_7QError_Int_1_argbuf_r;
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_d;
  logic lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_1_argbuf_d;
  logic lizzieLet6_7QNone_Int_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_1_argbuf_d;
  logic lizzieLet6_7QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t m1acN_1_argbuf_d;
  logic m1acN_1_argbuf_r;
  Pointer_QTree_Int_t m2acO_2_2_argbuf_d;
  logic m2acO_2_2_argbuf_r;
  Pointer_QTree_Int_t m2acO_2_1_d;
  logic m2acO_2_1_r;
  Pointer_QTree_Int_t m2acO_2_2_d;
  logic m2acO_2_2_r;
  Pointer_QTree_Int_t m2acO_3_2_argbuf_d;
  logic m2acO_3_2_argbuf_r;
  Pointer_QTree_Int_t m2acO_3_1_d;
  logic m2acO_3_1_r;
  Pointer_QTree_Int_t m2acO_3_2_d;
  logic m2acO_3_2_r;
  Pointer_QTree_Int_t m2acO_4_1_argbuf_d;
  logic m2acO_4_1_argbuf_r;
  Pointer_QTree_Int_t macF_1_argbuf_d;
  logic macF_1_argbuf_r;
  Pointer_QTree_Int_t mack_1_argbuf_d;
  logic mack_1_argbuf_r;
  Pointer_QTree_Int_t mack_1_d;
  logic mack_1_r;
  Pointer_QTree_Int_t mack_2_d;
  logic mack_2_r;
  Go_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_r;
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_r;
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_r;
  Go_t go_13_1_d;
  logic go_13_1_r;
  Go_t go_13_2_d;
  logic go_13_2_r;
  Pointer_QTree_Int_t mack_1_1_argbuf_d;
  logic mack_1_1_argbuf_r;
  Pointer_MaskQTree_t mskacl_1_1_argbuf_d;
  logic mskacl_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  Go_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_r ;
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_r ;
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_r ;
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_r ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_r ;
  MyDTInt_Int_Int_t gacD_1_1_argbuf_d;
  logic gacD_1_1_argbuf_r;
  Go_t go_14_1_d;
  logic go_14_1_r;
  Go_t go_14_2_d;
  logic go_14_2_r;
  MyDTInt_Bool_t isZacC_1_1_argbuf_d;
  logic isZacC_1_1_argbuf_r;
  Pointer_QTree_Int_t macF_1_1_argbuf_d;
  logic macF_1_1_argbuf_r;
  Int_t \v'acE_1_1_argbuf_d ;
  logic \v'acE_1_1_argbuf_r ;
  Pointer_QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_MaskQTree_t mskacl_1_argbuf_d;
  logic mskacl_1_argbuf_r;
  Pointer_QTree_Int_t q1acH_3_1_argbuf_d;
  logic q1acH_3_1_argbuf_r;
  Pointer_QTree_Int_t q1acQ_3_1_argbuf_d;
  logic q1acQ_3_1_argbuf_r;
  Pointer_QTree_Int_t q1acV_1_argbuf_d;
  logic q1acV_1_argbuf_r;
  Pointer_MaskQTree_t q1acm_3_1_argbuf_d;
  logic q1acm_3_1_argbuf_r;
  Pointer_QTree_Int_t q2acI_2_1_argbuf_d;
  logic q2acI_2_1_argbuf_r;
  Pointer_QTree_Int_t q2acR_2_1_argbuf_d;
  logic q2acR_2_1_argbuf_r;
  Pointer_QTree_Int_t q2acW_1_1_argbuf_d;
  logic q2acW_1_1_argbuf_r;
  Pointer_MaskQTree_t q2acn_2_1_argbuf_d;
  logic q2acn_2_1_argbuf_r;
  Pointer_QTree_Int_t q3acJ_1_1_argbuf_d;
  logic q3acJ_1_1_argbuf_r;
  Pointer_QTree_Int_t q3acS_1_1_argbuf_d;
  logic q3acS_1_1_argbuf_r;
  Pointer_QTree_Int_t q3acX_2_1_argbuf_d;
  logic q3acX_2_1_argbuf_r;
  Pointer_MaskQTree_t q3aco_1_1_argbuf_d;
  logic q3aco_1_1_argbuf_r;
  Pointer_QTree_Int_t q4acK_1_argbuf_d;
  logic q4acK_1_argbuf_r;
  Pointer_QTree_Int_t q4acT_1_argbuf_d;
  logic q4acT_1_argbuf_r;
  Pointer_QTree_Int_t q4acY_3_1_argbuf_d;
  logic q4acY_3_1_argbuf_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_Int_t lizzieLet26_1_d;
  logic lizzieLet26_1_r;
  CT$wnnz_Int_t lizzieLet26_2_d;
  logic lizzieLet26_2_r;
  CT$wnnz_Int_t lizzieLet26_3_d;
  logic lizzieLet26_3_r;
  CT$wnnz_Int_t lizzieLet26_4_d;
  logic lizzieLet26_4_r;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_1_d;
  logic lizzieLet30_1_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_2_d;
  logic lizzieLet30_2_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_3_d;
  logic lizzieLet30_3_r;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4_d;
  logic lizzieLet30_4_r;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r;
  CTmain_mask_Int_t lizzieLet35_1_d;
  logic lizzieLet35_1_r;
  CTmain_mask_Int_t lizzieLet35_2_d;
  logic lizzieLet35_2_r;
  CTmain_mask_Int_t lizzieLet35_3_d;
  logic lizzieLet35_3_r;
  CTmain_mask_Int_t lizzieLet35_4_d;
  logic lizzieLet35_4_r;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r ;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet40_1_d;
  logic lizzieLet40_1_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet40_2_d;
  logic lizzieLet40_2_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet40_3_d;
  logic lizzieLet40_3_r;
  \CTmap''_map''_Int_Int_Int_t  lizzieLet40_4_d;
  logic lizzieLet40_4_r;
  MaskQTree_t readPointer_MaskQTreemskacl_1_argbuf_rwb_d;
  logic readPointer_MaskQTreemskacl_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet10_1_1_d;
  logic lizzieLet10_1_1_r;
  MaskQTree_t lizzieLet10_1_2_d;
  logic lizzieLet10_1_2_r;
  MaskQTree_t lizzieLet10_1_3_d;
  logic lizzieLet10_1_3_r;
  MaskQTree_t lizzieLet10_1_4_d;
  logic lizzieLet10_1_4_r;
  MaskQTree_t lizzieLet10_1_5_d;
  logic lizzieLet10_1_5_r;
  MaskQTree_t lizzieLet10_1_6_d;
  logic lizzieLet10_1_6_r;
  QTree_Int_t readPointer_QTree_Intm1acN_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1acN_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Int_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Int_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Int_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Int_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Int_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t lizzieLet6_7_d;
  logic lizzieLet6_7_r;
  QTree_Int_t readPointer_QTree_IntmacF_1_argbuf_rwb_d;
  logic readPointer_QTree_IntmacF_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet17_1_d;
  logic lizzieLet17_1_r;
  QTree_Int_t lizzieLet17_2_d;
  logic lizzieLet17_2_r;
  QTree_Int_t lizzieLet17_3_d;
  logic lizzieLet17_3_r;
  QTree_Int_t lizzieLet17_4_d;
  logic lizzieLet17_4_r;
  QTree_Int_t lizzieLet17_5_d;
  logic lizzieLet17_5_r;
  QTree_Int_t lizzieLet17_6_d;
  logic lizzieLet17_6_r;
  QTree_Int_t lizzieLet17_7_d;
  logic lizzieLet17_7_r;
  QTree_Int_t readPointer_QTree_Intmack_1_argbuf_rwb_d;
  logic readPointer_QTree_Intmack_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intwsxl_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_1_argbuf_d;
  logic sc_0_11_1_argbuf_r;
  Pointer_CTmain_mask_Int_t sc_0_15_1_argbuf_d;
  logic sc_0_15_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_1_argbuf_d;
  logic sc_0_19_1_argbuf_r;
  Pointer_CT$wnnz_Int_t sc_0_7_1_argbuf_d;
  logic sc_0_7_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_1_argbuf_d;
  logic scfarg_0_3_1_argbuf_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1acr_3_1_argbuf_d;
  logic t1acr_3_1_argbuf_r;
  Pointer_QTree_Int_t t2acs_2_1_argbuf_d;
  logic t2acs_2_1_argbuf_r;
  Pointer_QTree_Int_t t3act_1_1_argbuf_d;
  logic t3act_1_1_argbuf_r;
  Pointer_QTree_Int_t t4acu_1_argbuf_d;
  logic t4acu_1_argbuf_r;
  Int_t \v'acE_2_2_argbuf_d ;
  logic \v'acE_2_2_argbuf_r ;
  Int_t \v'acE_2_1_d ;
  logic \v'acE_2_1_r ;
  Int_t \v'acE_2_2_d ;
  logic \v'acE_2_2_r ;
  Int_t \v'acE_3_2_argbuf_d ;
  logic \v'acE_3_2_argbuf_r ;
  Int_t \v'acE_3_1_d ;
  logic \v'acE_3_1_r ;
  Int_t \v'acE_3_2_d ;
  logic \v'acE_3_2_r ;
  Int_t \v'acE_4_1_argbuf_d ;
  logic \v'acE_4_1_argbuf_r ;
  Int_t vacG_1_argbuf_d;
  logic vacG_1_argbuf_r;
  Int_t vacP_1_argbuf_d;
  logic vacP_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Int_Int_Int_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_d;
  logic writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Int_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca3_3_1_argbuf_d;
  logic sca3_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca2_3_1_argbuf_d;
  logic sca2_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca1_3_1_argbuf_d;
  logic sca1_3_1_argbuf_r;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sca0_3_1_argbuf_d;
  logic sca0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet14_2_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet16_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet44_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_3_1_argbuf_d;
  logic contRet_0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Int_t wsxl_1_1_argbuf_d;
  logic wsxl_1_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CT$wnnz_Int_t wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_d;
  logic wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  CT$wnnz_Int_t wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  logic wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r;
  \Int#_t  es_6_1ww2XyF_1_1_Add32_d;
  logic es_6_1ww2XyF_1_1_Add32_r;
  \Int#_t  wwsxo_4_1ww1XyC_2_1_Add32_d;
  logic wwsxo_4_1ww1XyC_2_1_Add32_r;
  Int_t xac0_1_argbuf_d;
  logic xac0_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go_5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go),
                                (go__11,Go),
                                (go__12,Go),
                                (go__13,Go)] */
  logic [12:0] sourceGo_emitted;
  logic [12:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign go__11_d = (sourceGo_d[0] && (! sourceGo_emitted[10]));
  assign go__12_d = (sourceGo_d[0] && (! sourceGo_emitted[11]));
  assign go__13_d = (sourceGo_d[0] && (! sourceGo_emitted[12]));
  assign sourceGo_done = (sourceGo_emitted | ({go__13_d[0],
                                               go__12_d[0],
                                               go__11_d[0],
                                               go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go_5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__13_r,
                                                             go__12_r,
                                                             go__11_r,
                                                             go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go_5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 13'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 13'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go__6,Go) > (initHP_CT$wnnz_Int,Word16#) */
  assign initHP_CT$wnnz_Int_d = {16'd0, go__6_d[0]};
  assign go__6_r = initHP_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz_Int1,Go) > (incrHP_CT$wnnz_Int,Word16#) */
  assign incrHP_CT$wnnz_Int_d = {16'd1, incrHP_CT$wnnz_Int1_d[0]};
  assign incrHP_CT$wnnz_Int1_r = incrHP_CT$wnnz_Int_r;
  
  /* merge (Ty Go) : [(go__7,Go),
                 (incrHP_CT$wnnz_Int2,Go)] > (incrHP_mergeCT$wnnz_Int,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_Int_selected;
  logic [1:0] incrHP_mergeCT$wnnz_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_Int_select))
        incrHP_mergeCT$wnnz_Int_selected = incrHP_mergeCT$wnnz_Int_select;
      else
        if (go__7_d[0]) incrHP_mergeCT$wnnz_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz_Int2_d[0])
          incrHP_mergeCT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_select <= (incrHP_mergeCT$wnnz_Int_r ? 2'd0 :
                                         incrHP_mergeCT$wnnz_Int_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_Int_selected[0])
      incrHP_mergeCT$wnnz_Int_d = go__7_d;
    else if (incrHP_mergeCT$wnnz_Int_selected[1])
      incrHP_mergeCT$wnnz_Int_d = incrHP_CT$wnnz_Int2_d;
    else incrHP_mergeCT$wnnz_Int_d = 1'd0;
  assign {incrHP_CT$wnnz_Int2_r,
          go__7_r} = (incrHP_mergeCT$wnnz_Int_r ? incrHP_mergeCT$wnnz_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_Int_buf,Go) > [(incrHP_CT$wnnz_Int1,Go),
                                                   (incrHP_CT$wnnz_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_done;
  assign incrHP_CT$wnnz_Int1_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[0]));
  assign incrHP_CT$wnnz_Int2_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_Int_buf_done = (incrHP_mergeCT$wnnz_Int_buf_emitted | ({incrHP_CT$wnnz_Int2_d[0],
                                                                                     incrHP_CT$wnnz_Int1_d[0]} & {incrHP_CT$wnnz_Int2_r,
                                                                                                                  incrHP_CT$wnnz_Int1_r}));
  assign incrHP_mergeCT$wnnz_Int_buf_r = (& incrHP_mergeCT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_buf_emitted <= (incrHP_mergeCT$wnnz_Int_buf_r ? 2'd0 :
                                              incrHP_mergeCT$wnnz_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz_Int,Word16#) (forkHP1_CT$wnnz_Int,Word16#) > (addHP_CT$wnnz_Int,Word16#) */
  assign addHP_CT$wnnz_Int_d = {(incrHP_CT$wnnz_Int_d[16:1] + forkHP1_CT$wnnz_Int_d[16:1]),
                                (incrHP_CT$wnnz_Int_d[0] && forkHP1_CT$wnnz_Int_d[0])};
  assign {incrHP_CT$wnnz_Int_r,
          forkHP1_CT$wnnz_Int_r} = {2 {(addHP_CT$wnnz_Int_r && addHP_CT$wnnz_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz_Int,Word16#),
                      (addHP_CT$wnnz_Int,Word16#)] > (mergeHP_CT$wnnz_Int,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_Int_selected;
  logic [1:0] mergeHP_CT$wnnz_Int_select;
  always_comb
    begin
      mergeHP_CT$wnnz_Int_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_Int_select))
        mergeHP_CT$wnnz_Int_selected = mergeHP_CT$wnnz_Int_select;
      else
        if (initHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_select <= 2'd0;
    else
      mergeHP_CT$wnnz_Int_select <= (mergeHP_CT$wnnz_Int_r ? 2'd0 :
                                     mergeHP_CT$wnnz_Int_selected);
  always_comb
    if (mergeHP_CT$wnnz_Int_selected[0])
      mergeHP_CT$wnnz_Int_d = initHP_CT$wnnz_Int_d;
    else if (mergeHP_CT$wnnz_Int_selected[1])
      mergeHP_CT$wnnz_Int_d = addHP_CT$wnnz_Int_d;
    else mergeHP_CT$wnnz_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_Int_r,
          initHP_CT$wnnz_Int_r} = (mergeHP_CT$wnnz_Int_r ? mergeHP_CT$wnnz_Int_selected :
                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz_Int,Go) > (incrHP_mergeCT$wnnz_Int_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_d;
  logic incrHP_mergeCT$wnnz_Int_bufchan_r;
  assign incrHP_mergeCT$wnnz_Int_r = ((! incrHP_mergeCT$wnnz_Int_bufchan_d[0]) || incrHP_mergeCT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_Int_r)
        incrHP_mergeCT$wnnz_Int_bufchan_d <= incrHP_mergeCT$wnnz_Int_d;
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_buf;
  assign incrHP_mergeCT$wnnz_Int_bufchan_r = (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_Int_buf_d = (incrHP_mergeCT$wnnz_Int_bufchan_buf[0] ? incrHP_mergeCT$wnnz_Int_bufchan_buf :
                                          incrHP_mergeCT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_Int_buf_r && incrHP_mergeCT$wnnz_Int_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_Int_buf_r) && (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= incrHP_mergeCT$wnnz_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz_Int,Word16#) > (mergeHP_CT$wnnz_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_d;
  logic mergeHP_CT$wnnz_Int_bufchan_r;
  assign mergeHP_CT$wnnz_Int_r = ((! mergeHP_CT$wnnz_Int_bufchan_d[0]) || mergeHP_CT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_Int_r)
        mergeHP_CT$wnnz_Int_bufchan_d <= mergeHP_CT$wnnz_Int_d;
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_buf;
  assign mergeHP_CT$wnnz_Int_bufchan_r = (! mergeHP_CT$wnnz_Int_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_Int_buf_d = (mergeHP_CT$wnnz_Int_bufchan_buf[0] ? mergeHP_CT$wnnz_Int_bufchan_buf :
                                      mergeHP_CT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_Int_buf_r && mergeHP_CT$wnnz_Int_bufchan_buf[0]))
        mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_Int_buf_r) && (! mergeHP_CT$wnnz_Int_bufchan_buf[0])))
        mergeHP_CT$wnnz_Int_bufchan_buf <= mergeHP_CT$wnnz_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_Int_buf,Word16#) > [(forkHP1_CT$wnnz_Int,Word16#),
                                                         (forkHP1_CT$wnnz_In2,Word16#),
                                                         (forkHP1_CT$wnnz_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_Int_buf_done;
  assign forkHP1_CT$wnnz_Int_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[0]))};
  assign forkHP1_CT$wnnz_In2_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[1]))};
  assign forkHP1_CT$wnnz_In3_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_Int_buf_done = (mergeHP_CT$wnnz_Int_buf_emitted | ({forkHP1_CT$wnnz_In3_d[0],
                                                                             forkHP1_CT$wnnz_In2_d[0],
                                                                             forkHP1_CT$wnnz_Int_d[0]} & {forkHP1_CT$wnnz_In3_r,
                                                                                                          forkHP1_CT$wnnz_In2_r,
                                                                                                          forkHP1_CT$wnnz_Int_r}));
  assign mergeHP_CT$wnnz_Int_buf_r = (& mergeHP_CT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_Int_buf_emitted <= (mergeHP_CT$wnnz_Int_buf_r ? 3'd0 :
                                          mergeHP_CT$wnnz_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz_Int) : [(dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int),
                                    (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int)] > (memMergeChoice_CT$wnnz_Int,C2) (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  logic [1:0] dconReadIn_CT$wnnz_Int_select_d;
  assign dconReadIn_CT$wnnz_Int_select_d = ((| dconReadIn_CT$wnnz_Int_select_q) ? dconReadIn_CT$wnnz_Int_select_q :
                                            (dconReadIn_CT$wnnz_Int_d[0] ? 2'd1 :
                                             (dconWriteIn_CT$wnnz_Int_d[0] ? 2'd2 :
                                              2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_select_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                          dconReadIn_CT$wnnz_Int_select_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_emit_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                        dconReadIn_CT$wnnz_Int_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_d;
  assign dconReadIn_CT$wnnz_Int_emit_d = (dconReadIn_CT$wnnz_Int_emit_q | ({memMergeChoice_CT$wnnz_Int_d[0],
                                                                            memMergeIn_CT$wnnz_Int_d[0]} & {memMergeChoice_CT$wnnz_Int_r,
                                                                                                            memMergeIn_CT$wnnz_Int_r}));
  logic dconReadIn_CT$wnnz_Int_done;
  assign dconReadIn_CT$wnnz_Int_done = (& dconReadIn_CT$wnnz_Int_emit_d);
  assign {dconWriteIn_CT$wnnz_Int_r,
          dconReadIn_CT$wnnz_Int_r} = (dconReadIn_CT$wnnz_Int_done ? dconReadIn_CT$wnnz_Int_select_d :
                                       2'd0);
  assign memMergeIn_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconReadIn_CT$wnnz_Int_d :
                                     ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconWriteIn_CT$wnnz_Int_d :
                                      {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz_Int,
      Ty MemOut_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) > (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) */
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_din;
  logic [114:0] memOut_CT$wnnz_Int_q;
  logic memOut_CT$wnnz_Int_valid;
  logic memMergeIn_CT$wnnz_Int_dbuf_we;
  logic memOut_CT$wnnz_Int_we;
  assign memMergeIn_CT$wnnz_Int_dbuf_din = memMergeIn_CT$wnnz_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_Int_dbuf_address = memMergeIn_CT$wnnz_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_Int_dbuf_we = (memMergeIn_CT$wnnz_Int_dbuf_d[1:1] && memMergeIn_CT$wnnz_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_Int_we <= 1'd0;
        memOut_CT$wnnz_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_Int_we <= memMergeIn_CT$wnnz_Int_dbuf_we;
        memOut_CT$wnnz_Int_valid <= memMergeIn_CT$wnnz_Int_dbuf_d[0];
        if (memMergeIn_CT$wnnz_Int_dbuf_we)
          begin
            memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address] <= memMergeIn_CT$wnnz_Int_dbuf_din;
            memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_din;
          end
        else
          memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address];
      end
  assign memOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_q,
                                 memOut_CT$wnnz_Int_we,
                                 memOut_CT$wnnz_Int_valid};
  assign memMergeIn_CT$wnnz_Int_dbuf_r = ((! memOut_CT$wnnz_Int_valid) || memOut_CT$wnnz_Int_r);
  logic [31:0] profiling_MemIn_CT$wnnz_Int_read;
  logic [31:0] profiling_MemIn_CT$wnnz_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_Int_write <= 0;
        profiling_MemIn_CT$wnnz_Int_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_Int_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_Int_write <= (profiling_MemIn_CT$wnnz_Int_write + 1);
      else
        if ((memOut_CT$wnnz_Int_valid == 1'd1))
          profiling_MemIn_CT$wnnz_Int_read <= (profiling_MemIn_CT$wnnz_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz_Int) : (memMergeChoice_CT$wnnz_Int,C2) (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) > [(memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int),
                                                                                                                (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int)] */
  logic [1:0] memOut_CT$wnnz_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_Int_d[0] && memOut_CT$wnnz_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_Int_d[1:1])
        1'd0: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                     memOut_CT$wnnz_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                      memOut_CT$wnnz_Int_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_Int_dbuf_r = (| (memOut_CT$wnnz_Int_dbuf_onehotd & {memWriteOut_CT$wnnz_Int_r,
                                                                            memReadOut_CT$wnnz_Int_r}));
  assign memMergeChoice_CT$wnnz_Int_r = memOut_CT$wnnz_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) */
  assign memMergeIn_CT$wnnz_Int_rbuf_r = ((! memMergeIn_CT$wnnz_Int_dbuf_d[0]) || memMergeIn_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wnnz_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_Int_rbuf_r)
        memMergeIn_CT$wnnz_Int_dbuf_d <= memMergeIn_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) */
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_buf;
  assign memMergeIn_CT$wnnz_Int_r = (! memMergeIn_CT$wnnz_Int_buf[0]);
  assign memMergeIn_CT$wnnz_Int_rbuf_d = (memMergeIn_CT$wnnz_Int_buf[0] ? memMergeIn_CT$wnnz_Int_buf :
                                          memMergeIn_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_Int_rbuf_r && memMergeIn_CT$wnnz_Int_buf[0]))
        memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_Int_rbuf_r) && (! memMergeIn_CT$wnnz_Int_buf[0])))
        memMergeIn_CT$wnnz_Int_buf <= memMergeIn_CT$wnnz_Int_d;
  
  /* dbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) */
  assign memOut_CT$wnnz_Int_rbuf_r = ((! memOut_CT$wnnz_Int_dbuf_d[0]) || memOut_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_Int_rbuf_r)
        memOut_CT$wnnz_Int_dbuf_d <= memOut_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) */
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_buf;
  assign memOut_CT$wnnz_Int_r = (! memOut_CT$wnnz_Int_buf[0]);
  assign memOut_CT$wnnz_Int_rbuf_d = (memOut_CT$wnnz_Int_buf[0] ? memOut_CT$wnnz_Int_buf :
                                      memOut_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_Int_rbuf_r && memOut_CT$wnnz_Int_buf[0]))
        memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_Int_rbuf_r) && (! memOut_CT$wnnz_Int_buf[0])))
        memOut_CT$wnnz_Int_buf <= memOut_CT$wnnz_Int_d;
  
  /* destruct (Ty Pointer_CT$wnnz_Int,
          Dcon Pointer_CT$wnnz_Int) : (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) > [(destructReadIn_CT$wnnz_Int,Word16#)] */
  assign destructReadIn_CT$wnnz_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                         scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon ReadIn_CT$wnnz_Int) : [(destructReadIn_CT$wnnz_Int,Word16#)] > (dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconReadIn_CT$wnnz_Int_d = ReadIn_CT$wnnz_Int_dc((& {destructReadIn_CT$wnnz_Int_d[0]}), destructReadIn_CT$wnnz_Int_d);
  assign {destructReadIn_CT$wnnz_Int_r} = {1 {(dconReadIn_CT$wnnz_Int_r && dconReadIn_CT$wnnz_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz_Int,
          Dcon ReadOut_CT$wnnz_Int) : (memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > [(readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int)] */
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_Int_d[116:2],
                                                       memReadOut_CT$wnnz_Int_d[0]};
  assign memReadOut_CT$wnnz_Int_r = readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wnnz_Int) : [(lizzieLet0_1_argbuf,CT$wnnz_Int),
                              (lizzieLet27_1_argbuf,CT$wnnz_Int),
                              (lizzieLet28_1_argbuf,CT$wnnz_Int),
                              (lizzieLet29_1_argbuf,CT$wnnz_Int),
                              (lizzieLet5_1_argbuf,CT$wnnz_Int)] > (writeMerge_choice_CT$wnnz_Int,C5) (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet27_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet28_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet29_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet5_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_Int_d[0],
                                                                      writeMerge_data_CT$wnnz_Int_d[0]} & {writeMerge_choice_CT$wnnz_Int_r,
                                                                                                           writeMerge_data_CT$wnnz_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet5_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                          ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                              {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                            ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz_Int) : (writeMerge_choice_CT$wnnz_Int,C5) (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet27_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet29_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int)] */
  logic [4:0] demuxWriteResult_CT$wnnz_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_Int_d[0] && demuxWriteResult_CT$wnnz_Int_d[0]))
      unique case (writeMerge_choice_CT$wnnz_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[0]};
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[1]};
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[2]};
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[3]};
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_Int_r = (| (demuxWriteResult_CT$wnnz_Int_onehotd & {writeCT$wnnz_IntlizzieLet5_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet29_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet28_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet27_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_Int_r = demuxWriteResult_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon WriteIn_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In2,Word16#),
                                   (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int)] > (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconWriteIn_CT$wnnz_Int_d = WriteIn_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In2_d[0],
                                                                writeMerge_data_CT$wnnz_Int_d[0]}), forkHP1_CT$wnnz_In2_d, writeMerge_data_CT$wnnz_Int_d);
  assign {forkHP1_CT$wnnz_In2_r,
          writeMerge_data_CT$wnnz_Int_r} = {2 {(dconWriteIn_CT$wnnz_Int_r && dconWriteIn_CT$wnnz_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz_Int,
      Dcon Pointer_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In3,Word16#)] > (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) */
  assign dconPtr_CT$wnnz_Int_d = Pointer_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In3_d[0]}), forkHP1_CT$wnnz_In3_d);
  assign {forkHP1_CT$wnnz_In3_r} = {1 {(dconPtr_CT$wnnz_Int_r && dconPtr_CT$wnnz_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz_Int,
       Ty Pointer_CT$wnnz_Int) : (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(_54,Pointer_CT$wnnz_Int),
                                                                                                                           (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int)] */
  logic [1:0] dconPtr_CT$wnnz_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_Int_d[0] && dconPtr_CT$wnnz_Int_d[0]))
      unique case (memWriteOut_CT$wnnz_Int_d[1:1])
        1'd0: dconPtr_CT$wnnz_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_Int_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_Int_onehotd = 2'd0;
  assign _54_d = {dconPtr_CT$wnnz_Int_d[16:1],
                  dconPtr_CT$wnnz_Int_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_Int_d = {dconPtr_CT$wnnz_Int_d[16:1],
                                           dconPtr_CT$wnnz_Int_onehotd[1]};
  assign dconPtr_CT$wnnz_Int_r = (| (dconPtr_CT$wnnz_Int_onehotd & {demuxWriteResult_CT$wnnz_Int_r,
                                                                    _54_r}));
  assign memWriteOut_CT$wnnz_Int_r = dconPtr_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C4,
           Ty Pointer_QTree_Int) : [(m1acN_1_argbuf,Pointer_QTree_Int),
                                    (macF_1_argbuf,Pointer_QTree_Int),
                                    (mack_1_argbuf,Pointer_QTree_Int),
                                    (wsxl_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C4) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [3:0] m1acN_1_argbuf_select_d;
  assign m1acN_1_argbuf_select_d = ((| m1acN_1_argbuf_select_q) ? m1acN_1_argbuf_select_q :
                                    (m1acN_1_argbuf_d[0] ? 4'd1 :
                                     (macF_1_argbuf_d[0] ? 4'd2 :
                                      (mack_1_argbuf_d[0] ? 4'd4 :
                                       (wsxl_1_1_argbuf_d[0] ? 4'd8 :
                                        4'd0)))));
  logic [3:0] m1acN_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acN_1_argbuf_select_q <= 4'd0;
    else
      m1acN_1_argbuf_select_q <= (m1acN_1_argbuf_done ? 4'd0 :
                                  m1acN_1_argbuf_select_d);
  logic [1:0] m1acN_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acN_1_argbuf_emit_q <= 2'd0;
    else
      m1acN_1_argbuf_emit_q <= (m1acN_1_argbuf_done ? 2'd0 :
                                m1acN_1_argbuf_emit_d);
  logic [1:0] m1acN_1_argbuf_emit_d;
  assign m1acN_1_argbuf_emit_d = (m1acN_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1acN_1_argbuf_done;
  assign m1acN_1_argbuf_done = (& m1acN_1_argbuf_emit_d);
  assign {wsxl_1_1_argbuf_r,
          mack_1_argbuf_r,
          macF_1_argbuf_r,
          m1acN_1_argbuf_r} = (m1acN_1_argbuf_done ? m1acN_1_argbuf_select_d :
                               4'd0);
  assign readMerge_data_QTree_Int_d = ((m1acN_1_argbuf_select_d[0] && (! m1acN_1_argbuf_emit_q[0])) ? m1acN_1_argbuf_d :
                                       ((m1acN_1_argbuf_select_d[1] && (! m1acN_1_argbuf_emit_q[0])) ? macF_1_argbuf_d :
                                        ((m1acN_1_argbuf_select_d[2] && (! m1acN_1_argbuf_emit_q[0])) ? mack_1_argbuf_d :
                                         ((m1acN_1_argbuf_select_d[3] && (! m1acN_1_argbuf_emit_q[0])) ? wsxl_1_1_argbuf_d :
                                          {16'd0, 1'd0}))));
  assign readMerge_choice_QTree_Int_d = ((m1acN_1_argbuf_select_d[0] && (! m1acN_1_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                         ((m1acN_1_argbuf_select_d[1] && (! m1acN_1_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                          ((m1acN_1_argbuf_select_d[2] && (! m1acN_1_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                           ((m1acN_1_argbuf_select_d[3] && (! m1acN_1_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                            {2'd0, 1'd0}))));
  
  /* demux (Ty C4,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C4) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1acN_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntmacF_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intmack_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intwsxl_1_1_argbuf,QTree_Int)] */
  logic [3:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 4'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 4'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 4'd4;
        2'd3: destructReadOut_QTree_Int_onehotd = 4'd8;
        default: destructReadOut_QTree_Int_onehotd = 4'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 4'd0;
  assign readPointer_QTree_Intm1acN_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_IntmacF_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intmack_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_Intwsxl_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[3]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intwsxl_1_1_argbuf_r,
                                                                                readPointer_QTree_Intmack_1_argbuf_r,
                                                                                readPointer_QTree_IntmacF_1_argbuf_r,
                                                                                readPointer_QTree_Intm1acN_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C14,
           Ty QTree_Int) : [(lizzieLet11_1_1_argbuf,QTree_Int),
                            (lizzieLet13_1_argbuf,QTree_Int),
                            (lizzieLet14_2_1_argbuf,QTree_Int),
                            (lizzieLet16_1_1_argbuf,QTree_Int),
                            (lizzieLet18_1_argbuf,QTree_Int),
                            (lizzieLet19_1_argbuf,QTree_Int),
                            (lizzieLet20_1_argbuf,QTree_Int),
                            (lizzieLet22_1_argbuf,QTree_Int),
                            (lizzieLet34_1_argbuf,QTree_Int),
                            (lizzieLet39_1_argbuf,QTree_Int),
                            (lizzieLet44_1_argbuf,QTree_Int),
                            (lizzieLet7_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C14) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [13:0] lizzieLet11_1_1_argbuf_select_d;
  assign lizzieLet11_1_1_argbuf_select_d = ((| lizzieLet11_1_1_argbuf_select_q) ? lizzieLet11_1_1_argbuf_select_q :
                                            (lizzieLet11_1_1_argbuf_d[0] ? 14'd1 :
                                             (lizzieLet13_1_argbuf_d[0] ? 14'd2 :
                                              (lizzieLet14_2_1_argbuf_d[0] ? 14'd4 :
                                               (lizzieLet16_1_1_argbuf_d[0] ? 14'd8 :
                                                (lizzieLet18_1_argbuf_d[0] ? 14'd16 :
                                                 (lizzieLet19_1_argbuf_d[0] ? 14'd32 :
                                                  (lizzieLet20_1_argbuf_d[0] ? 14'd64 :
                                                   (lizzieLet22_1_argbuf_d[0] ? 14'd128 :
                                                    (lizzieLet34_1_argbuf_d[0] ? 14'd256 :
                                                     (lizzieLet39_1_argbuf_d[0] ? 14'd512 :
                                                      (lizzieLet44_1_argbuf_d[0] ? 14'd1024 :
                                                       (lizzieLet7_1_argbuf_d[0] ? 14'd2048 :
                                                        (lizzieLet9_1_argbuf_d[0] ? 14'd4096 :
                                                         (dummy_write_QTree_Int_d[0] ? 14'd8192 :
                                                          14'd0)))))))))))))));
  logic [13:0] lizzieLet11_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_select_q <= 14'd0;
    else
      lizzieLet11_1_1_argbuf_select_q <= (lizzieLet11_1_1_argbuf_done ? 14'd0 :
                                          lizzieLet11_1_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_1_argbuf_emit_q <= (lizzieLet11_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet11_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_d;
  assign lizzieLet11_1_1_argbuf_emit_d = (lizzieLet11_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                            writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                               writeMerge_data_QTree_Int_r}));
  logic lizzieLet11_1_1_argbuf_done;
  assign lizzieLet11_1_1_argbuf_done = (& lizzieLet11_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet44_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet14_2_1_argbuf_r,
          lizzieLet13_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r} = (lizzieLet11_1_1_argbuf_done ? lizzieLet11_1_1_argbuf_select_d :
                                       14'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                        ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_argbuf_d :
                                         ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet14_2_1_argbuf_d :
                                          ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet16_1_1_argbuf_d :
                                           ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                            ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                             ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                              ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                               ((lizzieLet11_1_1_argbuf_select_d[8] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                ((lizzieLet11_1_1_argbuf_select_d[9] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                                 ((lizzieLet11_1_1_argbuf_select_d[10] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet44_1_argbuf_d :
                                                  ((lizzieLet11_1_1_argbuf_select_d[11] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                   ((lizzieLet11_1_1_argbuf_select_d[12] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                    ((lizzieLet11_1_1_argbuf_select_d[13] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                     {66'd0, 1'd0}))))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C1_14_dc(1'd1) :
                                          ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C2_14_dc(1'd1) :
                                           ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C3_14_dc(1'd1) :
                                            ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C4_14_dc(1'd1) :
                                             ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C5_14_dc(1'd1) :
                                              ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C6_14_dc(1'd1) :
                                               ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C7_14_dc(1'd1) :
                                                ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C8_14_dc(1'd1) :
                                                 ((lizzieLet11_1_1_argbuf_select_d[8] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C9_14_dc(1'd1) :
                                                  ((lizzieLet11_1_1_argbuf_select_d[9] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C10_14_dc(1'd1) :
                                                   ((lizzieLet11_1_1_argbuf_select_d[10] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C11_14_dc(1'd1) :
                                                    ((lizzieLet11_1_1_argbuf_select_d[11] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C12_14_dc(1'd1) :
                                                     ((lizzieLet11_1_1_argbuf_select_d[12] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C13_14_dc(1'd1) :
                                                      ((lizzieLet11_1_1_argbuf_select_d[13] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C14_14_dc(1'd1) :
                                                       {4'd0, 1'd0}))))))))))))));
  
  /* demux (Ty C14,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C14) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet14_2_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet16_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet19_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet39_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet44_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [13:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[4:1])
        4'd0: demuxWriteResult_QTree_Int_onehotd = 14'd1;
        4'd1: demuxWriteResult_QTree_Int_onehotd = 14'd2;
        4'd2: demuxWriteResult_QTree_Int_onehotd = 14'd4;
        4'd3: demuxWriteResult_QTree_Int_onehotd = 14'd8;
        4'd4: demuxWriteResult_QTree_Int_onehotd = 14'd16;
        4'd5: demuxWriteResult_QTree_Int_onehotd = 14'd32;
        4'd6: demuxWriteResult_QTree_Int_onehotd = 14'd64;
        4'd7: demuxWriteResult_QTree_Int_onehotd = 14'd128;
        4'd8: demuxWriteResult_QTree_Int_onehotd = 14'd256;
        4'd9: demuxWriteResult_QTree_Int_onehotd = 14'd512;
        4'd10: demuxWriteResult_QTree_Int_onehotd = 14'd1024;
        4'd11: demuxWriteResult_QTree_Int_onehotd = 14'd2048;
        4'd12: demuxWriteResult_QTree_Int_onehotd = 14'd4096;
        4'd13: demuxWriteResult_QTree_Int_onehotd = 14'd8192;
        default: demuxWriteResult_QTree_Int_onehotd = 14'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 14'd0;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet13_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet14_2_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet16_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet19_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet39_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet44_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[11]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[12]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[13]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet44_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet39_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet34_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet22_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet20_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet19_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet18_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet16_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet14_2_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet13_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_53,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _53_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _53_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__8,Go) > (initHP_CTmain_mask_Int,Word16#) */
  assign initHP_CTmain_mask_Int_d = {16'd0, go__8_d[0]};
  assign go__8_r = initHP_CTmain_mask_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_mask_Int1,Go) > (incrHP_CTmain_mask_Int,Word16#) */
  assign incrHP_CTmain_mask_Int_d = {16'd1,
                                     incrHP_CTmain_mask_Int1_d[0]};
  assign incrHP_CTmain_mask_Int1_r = incrHP_CTmain_mask_Int_r;
  
  /* merge (Ty Go) : [(go__9,Go),
                 (incrHP_CTmain_mask_Int2,Go)] > (incrHP_mergeCTmain_mask_Int,Go) */
  logic [1:0] incrHP_mergeCTmain_mask_Int_selected;
  logic [1:0] incrHP_mergeCTmain_mask_Int_select;
  always_comb
    begin
      incrHP_mergeCTmain_mask_Int_selected = 2'd0;
      if ((| incrHP_mergeCTmain_mask_Int_select))
        incrHP_mergeCTmain_mask_Int_selected = incrHP_mergeCTmain_mask_Int_select;
      else
        if (go__9_d[0]) incrHP_mergeCTmain_mask_Int_selected[0] = 1'd1;
        else if (incrHP_CTmain_mask_Int2_d[0])
          incrHP_mergeCTmain_mask_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Int_select <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Int_select <= (incrHP_mergeCTmain_mask_Int_r ? 2'd0 :
                                             incrHP_mergeCTmain_mask_Int_selected);
  always_comb
    if (incrHP_mergeCTmain_mask_Int_selected[0])
      incrHP_mergeCTmain_mask_Int_d = go__9_d;
    else if (incrHP_mergeCTmain_mask_Int_selected[1])
      incrHP_mergeCTmain_mask_Int_d = incrHP_CTmain_mask_Int2_d;
    else incrHP_mergeCTmain_mask_Int_d = 1'd0;
  assign {incrHP_CTmain_mask_Int2_r,
          go__9_r} = (incrHP_mergeCTmain_mask_Int_r ? incrHP_mergeCTmain_mask_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_mask_Int_buf,Go) > [(incrHP_CTmain_mask_Int1,Go),
                                                       (incrHP_CTmain_mask_Int2,Go)] */
  logic [1:0] incrHP_mergeCTmain_mask_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTmain_mask_Int_buf_done;
  assign incrHP_CTmain_mask_Int1_d = (incrHP_mergeCTmain_mask_Int_buf_d[0] && (! incrHP_mergeCTmain_mask_Int_buf_emitted[0]));
  assign incrHP_CTmain_mask_Int2_d = (incrHP_mergeCTmain_mask_Int_buf_d[0] && (! incrHP_mergeCTmain_mask_Int_buf_emitted[1]));
  assign incrHP_mergeCTmain_mask_Int_buf_done = (incrHP_mergeCTmain_mask_Int_buf_emitted | ({incrHP_CTmain_mask_Int2_d[0],
                                                                                             incrHP_CTmain_mask_Int1_d[0]} & {incrHP_CTmain_mask_Int2_r,
                                                                                                                              incrHP_CTmain_mask_Int1_r}));
  assign incrHP_mergeCTmain_mask_Int_buf_r = (& incrHP_mergeCTmain_mask_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Int_buf_emitted <= (incrHP_mergeCTmain_mask_Int_buf_r ? 2'd0 :
                                                  incrHP_mergeCTmain_mask_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_mask_Int,Word16#) (forkHP1_CTmain_mask_Int,Word16#) > (addHP_CTmain_mask_Int,Word16#) */
  assign addHP_CTmain_mask_Int_d = {(incrHP_CTmain_mask_Int_d[16:1] + forkHP1_CTmain_mask_Int_d[16:1]),
                                    (incrHP_CTmain_mask_Int_d[0] && forkHP1_CTmain_mask_Int_d[0])};
  assign {incrHP_CTmain_mask_Int_r,
          forkHP1_CTmain_mask_Int_r} = {2 {(addHP_CTmain_mask_Int_r && addHP_CTmain_mask_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_mask_Int,Word16#),
                      (addHP_CTmain_mask_Int,Word16#)] > (mergeHP_CTmain_mask_Int,Word16#) */
  logic [1:0] mergeHP_CTmain_mask_Int_selected;
  logic [1:0] mergeHP_CTmain_mask_Int_select;
  always_comb
    begin
      mergeHP_CTmain_mask_Int_selected = 2'd0;
      if ((| mergeHP_CTmain_mask_Int_select))
        mergeHP_CTmain_mask_Int_selected = mergeHP_CTmain_mask_Int_select;
      else
        if (initHP_CTmain_mask_Int_d[0])
          mergeHP_CTmain_mask_Int_selected[0] = 1'd1;
        else if (addHP_CTmain_mask_Int_d[0])
          mergeHP_CTmain_mask_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Int_select <= 2'd0;
    else
      mergeHP_CTmain_mask_Int_select <= (mergeHP_CTmain_mask_Int_r ? 2'd0 :
                                         mergeHP_CTmain_mask_Int_selected);
  always_comb
    if (mergeHP_CTmain_mask_Int_selected[0])
      mergeHP_CTmain_mask_Int_d = initHP_CTmain_mask_Int_d;
    else if (mergeHP_CTmain_mask_Int_selected[1])
      mergeHP_CTmain_mask_Int_d = addHP_CTmain_mask_Int_d;
    else mergeHP_CTmain_mask_Int_d = {16'd0, 1'd0};
  assign {addHP_CTmain_mask_Int_r,
          initHP_CTmain_mask_Int_r} = (mergeHP_CTmain_mask_Int_r ? mergeHP_CTmain_mask_Int_selected :
                                       2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_mask_Int,Go) > (incrHP_mergeCTmain_mask_Int_buf,Go) */
  Go_t incrHP_mergeCTmain_mask_Int_bufchan_d;
  logic incrHP_mergeCTmain_mask_Int_bufchan_r;
  assign incrHP_mergeCTmain_mask_Int_r = ((! incrHP_mergeCTmain_mask_Int_bufchan_d[0]) || incrHP_mergeCTmain_mask_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTmain_mask_Int_r)
        incrHP_mergeCTmain_mask_Int_bufchan_d <= incrHP_mergeCTmain_mask_Int_d;
  Go_t incrHP_mergeCTmain_mask_Int_bufchan_buf;
  assign incrHP_mergeCTmain_mask_Int_bufchan_r = (! incrHP_mergeCTmain_mask_Int_bufchan_buf[0]);
  assign incrHP_mergeCTmain_mask_Int_buf_d = (incrHP_mergeCTmain_mask_Int_bufchan_buf[0] ? incrHP_mergeCTmain_mask_Int_bufchan_buf :
                                              incrHP_mergeCTmain_mask_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTmain_mask_Int_buf_r && incrHP_mergeCTmain_mask_Int_bufchan_buf[0]))
        incrHP_mergeCTmain_mask_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTmain_mask_Int_buf_r) && (! incrHP_mergeCTmain_mask_Int_bufchan_buf[0])))
        incrHP_mergeCTmain_mask_Int_bufchan_buf <= incrHP_mergeCTmain_mask_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_mask_Int,Word16#) > (mergeHP_CTmain_mask_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTmain_mask_Int_bufchan_d;
  logic mergeHP_CTmain_mask_Int_bufchan_r;
  assign mergeHP_CTmain_mask_Int_r = ((! mergeHP_CTmain_mask_Int_bufchan_d[0]) || mergeHP_CTmain_mask_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTmain_mask_Int_r)
        mergeHP_CTmain_mask_Int_bufchan_d <= mergeHP_CTmain_mask_Int_d;
  \Word16#_t  mergeHP_CTmain_mask_Int_bufchan_buf;
  assign mergeHP_CTmain_mask_Int_bufchan_r = (! mergeHP_CTmain_mask_Int_bufchan_buf[0]);
  assign mergeHP_CTmain_mask_Int_buf_d = (mergeHP_CTmain_mask_Int_bufchan_buf[0] ? mergeHP_CTmain_mask_Int_bufchan_buf :
                                          mergeHP_CTmain_mask_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTmain_mask_Int_buf_r && mergeHP_CTmain_mask_Int_bufchan_buf[0]))
        mergeHP_CTmain_mask_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTmain_mask_Int_buf_r) && (! mergeHP_CTmain_mask_Int_bufchan_buf[0])))
        mergeHP_CTmain_mask_Int_bufchan_buf <= mergeHP_CTmain_mask_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_mask_Int_buf,Word16#) > [(forkHP1_CTmain_mask_Int,Word16#),
                                                             (forkHP1_CTmain_mask_In2,Word16#),
                                                             (forkHP1_CTmain_mask_In3,Word16#)] */
  logic [2:0] mergeHP_CTmain_mask_Int_buf_emitted;
  logic [2:0] mergeHP_CTmain_mask_Int_buf_done;
  assign forkHP1_CTmain_mask_Int_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[0]))};
  assign forkHP1_CTmain_mask_In2_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[1]))};
  assign forkHP1_CTmain_mask_In3_d = {mergeHP_CTmain_mask_Int_buf_d[16:1],
                                      (mergeHP_CTmain_mask_Int_buf_d[0] && (! mergeHP_CTmain_mask_Int_buf_emitted[2]))};
  assign mergeHP_CTmain_mask_Int_buf_done = (mergeHP_CTmain_mask_Int_buf_emitted | ({forkHP1_CTmain_mask_In3_d[0],
                                                                                     forkHP1_CTmain_mask_In2_d[0],
                                                                                     forkHP1_CTmain_mask_Int_d[0]} & {forkHP1_CTmain_mask_In3_r,
                                                                                                                      forkHP1_CTmain_mask_In2_r,
                                                                                                                      forkHP1_CTmain_mask_Int_r}));
  assign mergeHP_CTmain_mask_Int_buf_r = (& mergeHP_CTmain_mask_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTmain_mask_Int_buf_emitted <= (mergeHP_CTmain_mask_Int_buf_r ? 3'd0 :
                                              mergeHP_CTmain_mask_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_mask_Int) : [(dconReadIn_CTmain_mask_Int,MemIn_CTmain_mask_Int),
                                        (dconWriteIn_CTmain_mask_Int,MemIn_CTmain_mask_Int)] > (memMergeChoice_CTmain_mask_Int,C2) (memMergeIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  logic [1:0] dconReadIn_CTmain_mask_Int_select_d;
  assign dconReadIn_CTmain_mask_Int_select_d = ((| dconReadIn_CTmain_mask_Int_select_q) ? dconReadIn_CTmain_mask_Int_select_q :
                                                (dconReadIn_CTmain_mask_Int_d[0] ? 2'd1 :
                                                 (dconWriteIn_CTmain_mask_Int_d[0] ? 2'd2 :
                                                  2'd0)));
  logic [1:0] dconReadIn_CTmain_mask_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Int_select_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Int_select_q <= (dconReadIn_CTmain_mask_Int_done ? 2'd0 :
                                              dconReadIn_CTmain_mask_Int_select_d);
  logic [1:0] dconReadIn_CTmain_mask_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Int_emit_q <= (dconReadIn_CTmain_mask_Int_done ? 2'd0 :
                                            dconReadIn_CTmain_mask_Int_emit_d);
  logic [1:0] dconReadIn_CTmain_mask_Int_emit_d;
  assign dconReadIn_CTmain_mask_Int_emit_d = (dconReadIn_CTmain_mask_Int_emit_q | ({memMergeChoice_CTmain_mask_Int_d[0],
                                                                                    memMergeIn_CTmain_mask_Int_d[0]} & {memMergeChoice_CTmain_mask_Int_r,
                                                                                                                        memMergeIn_CTmain_mask_Int_r}));
  logic dconReadIn_CTmain_mask_Int_done;
  assign dconReadIn_CTmain_mask_Int_done = (& dconReadIn_CTmain_mask_Int_emit_d);
  assign {dconWriteIn_CTmain_mask_Int_r,
          dconReadIn_CTmain_mask_Int_r} = (dconReadIn_CTmain_mask_Int_done ? dconReadIn_CTmain_mask_Int_select_d :
                                           2'd0);
  assign memMergeIn_CTmain_mask_Int_d = ((dconReadIn_CTmain_mask_Int_select_d[0] && (! dconReadIn_CTmain_mask_Int_emit_q[0])) ? dconReadIn_CTmain_mask_Int_d :
                                         ((dconReadIn_CTmain_mask_Int_select_d[1] && (! dconReadIn_CTmain_mask_Int_emit_q[0])) ? dconWriteIn_CTmain_mask_Int_d :
                                          {132'd0, 1'd0}));
  assign memMergeChoice_CTmain_mask_Int_d = ((dconReadIn_CTmain_mask_Int_select_d[0] && (! dconReadIn_CTmain_mask_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                             ((dconReadIn_CTmain_mask_Int_select_d[1] && (! dconReadIn_CTmain_mask_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                              {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_mask_Int,
      Ty MemOut_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int_dbuf,MemIn_CTmain_mask_Int) > (memOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) */
  logic [114:0] memMergeIn_CTmain_mask_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTmain_mask_Int_dbuf_address;
  logic [114:0] memMergeIn_CTmain_mask_Int_dbuf_din;
  logic [114:0] memOut_CTmain_mask_Int_q;
  logic memOut_CTmain_mask_Int_valid;
  logic memMergeIn_CTmain_mask_Int_dbuf_we;
  logic memOut_CTmain_mask_Int_we;
  assign memMergeIn_CTmain_mask_Int_dbuf_din = memMergeIn_CTmain_mask_Int_dbuf_d[132:18];
  assign memMergeIn_CTmain_mask_Int_dbuf_address = memMergeIn_CTmain_mask_Int_dbuf_d[17:2];
  assign memMergeIn_CTmain_mask_Int_dbuf_we = (memMergeIn_CTmain_mask_Int_dbuf_d[1:1] && memMergeIn_CTmain_mask_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTmain_mask_Int_we <= 1'd0;
        memOut_CTmain_mask_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTmain_mask_Int_we <= memMergeIn_CTmain_mask_Int_dbuf_we;
        memOut_CTmain_mask_Int_valid <= memMergeIn_CTmain_mask_Int_dbuf_d[0];
        if (memMergeIn_CTmain_mask_Int_dbuf_we)
          begin
            memMergeIn_CTmain_mask_Int_dbuf_mem[memMergeIn_CTmain_mask_Int_dbuf_address] <= memMergeIn_CTmain_mask_Int_dbuf_din;
            memOut_CTmain_mask_Int_q <= memMergeIn_CTmain_mask_Int_dbuf_din;
          end
        else
          memOut_CTmain_mask_Int_q <= memMergeIn_CTmain_mask_Int_dbuf_mem[memMergeIn_CTmain_mask_Int_dbuf_address];
      end
  assign memOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_q,
                                     memOut_CTmain_mask_Int_we,
                                     memOut_CTmain_mask_Int_valid};
  assign memMergeIn_CTmain_mask_Int_dbuf_r = ((! memOut_CTmain_mask_Int_valid) || memOut_CTmain_mask_Int_r);
  logic [31:0] profiling_MemIn_CTmain_mask_Int_read;
  logic [31:0] profiling_MemIn_CTmain_mask_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTmain_mask_Int_write <= 0;
        profiling_MemIn_CTmain_mask_Int_read <= 0;
      end
    else
      if ((memMergeIn_CTmain_mask_Int_dbuf_we == 1'd1))
        profiling_MemIn_CTmain_mask_Int_write <= (profiling_MemIn_CTmain_mask_Int_write + 1);
      else
        if ((memOut_CTmain_mask_Int_valid == 1'd1))
          profiling_MemIn_CTmain_mask_Int_read <= (profiling_MemIn_CTmain_mask_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_mask_Int) : (memMergeChoice_CTmain_mask_Int,C2) (memOut_CTmain_mask_Int_dbuf,MemOut_CTmain_mask_Int) > [(memReadOut_CTmain_mask_Int,MemOut_CTmain_mask_Int),
                                                                                                                                (memWriteOut_CTmain_mask_Int,MemOut_CTmain_mask_Int)] */
  logic [1:0] memOut_CTmain_mask_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTmain_mask_Int_d[0] && memOut_CTmain_mask_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTmain_mask_Int_d[1:1])
        1'd0: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTmain_mask_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTmain_mask_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_dbuf_d[116:1],
                                         memOut_CTmain_mask_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTmain_mask_Int_d = {memOut_CTmain_mask_Int_dbuf_d[116:1],
                                          memOut_CTmain_mask_Int_dbuf_onehotd[1]};
  assign memOut_CTmain_mask_Int_dbuf_r = (| (memOut_CTmain_mask_Int_dbuf_onehotd & {memWriteOut_CTmain_mask_Int_r,
                                                                                    memReadOut_CTmain_mask_Int_r}));
  assign memMergeChoice_CTmain_mask_Int_r = memOut_CTmain_mask_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int_rbuf,MemIn_CTmain_mask_Int) > (memMergeIn_CTmain_mask_Int_dbuf,MemIn_CTmain_mask_Int) */
  assign memMergeIn_CTmain_mask_Int_rbuf_r = ((! memMergeIn_CTmain_mask_Int_dbuf_d[0]) || memMergeIn_CTmain_mask_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTmain_mask_Int_rbuf_r)
        memMergeIn_CTmain_mask_Int_dbuf_d <= memMergeIn_CTmain_mask_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTmain_mask_Int) : (memMergeIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) > (memMergeIn_CTmain_mask_Int_rbuf,MemIn_CTmain_mask_Int) */
  MemIn_CTmain_mask_Int_t memMergeIn_CTmain_mask_Int_buf;
  assign memMergeIn_CTmain_mask_Int_r = (! memMergeIn_CTmain_mask_Int_buf[0]);
  assign memMergeIn_CTmain_mask_Int_rbuf_d = (memMergeIn_CTmain_mask_Int_buf[0] ? memMergeIn_CTmain_mask_Int_buf :
                                              memMergeIn_CTmain_mask_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTmain_mask_Int_rbuf_r && memMergeIn_CTmain_mask_Int_buf[0]))
        memMergeIn_CTmain_mask_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTmain_mask_Int_rbuf_r) && (! memMergeIn_CTmain_mask_Int_buf[0])))
        memMergeIn_CTmain_mask_Int_buf <= memMergeIn_CTmain_mask_Int_d;
  
  /* dbuf (Ty MemOut_CTmain_mask_Int) : (memOut_CTmain_mask_Int_rbuf,MemOut_CTmain_mask_Int) > (memOut_CTmain_mask_Int_dbuf,MemOut_CTmain_mask_Int) */
  assign memOut_CTmain_mask_Int_rbuf_r = ((! memOut_CTmain_mask_Int_dbuf_d[0]) || memOut_CTmain_mask_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTmain_mask_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTmain_mask_Int_rbuf_r)
        memOut_CTmain_mask_Int_dbuf_d <= memOut_CTmain_mask_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTmain_mask_Int) : (memOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) > (memOut_CTmain_mask_Int_rbuf,MemOut_CTmain_mask_Int) */
  MemOut_CTmain_mask_Int_t memOut_CTmain_mask_Int_buf;
  assign memOut_CTmain_mask_Int_r = (! memOut_CTmain_mask_Int_buf[0]);
  assign memOut_CTmain_mask_Int_rbuf_d = (memOut_CTmain_mask_Int_buf[0] ? memOut_CTmain_mask_Int_buf :
                                          memOut_CTmain_mask_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTmain_mask_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTmain_mask_Int_rbuf_r && memOut_CTmain_mask_Int_buf[0]))
        memOut_CTmain_mask_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTmain_mask_Int_rbuf_r) && (! memOut_CTmain_mask_Int_buf[0])))
        memOut_CTmain_mask_Int_buf <= memOut_CTmain_mask_Int_d;
  
  /* destruct (Ty Pointer_CTmain_mask_Int,
          Dcon Pointer_CTmain_mask_Int) : (scfarg_0_2_1_argbuf,Pointer_CTmain_mask_Int) > [(destructReadIn_CTmain_mask_Int,Word16#)] */
  assign destructReadIn_CTmain_mask_Int_d = {scfarg_0_2_1_argbuf_d[16:1],
                                             scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTmain_mask_Int_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Int,
      Dcon ReadIn_CTmain_mask_Int) : [(destructReadIn_CTmain_mask_Int,Word16#)] > (dconReadIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  assign dconReadIn_CTmain_mask_Int_d = ReadIn_CTmain_mask_Int_dc((& {destructReadIn_CTmain_mask_Int_d[0]}), destructReadIn_CTmain_mask_Int_d);
  assign {destructReadIn_CTmain_mask_Int_r} = {1 {(dconReadIn_CTmain_mask_Int_r && dconReadIn_CTmain_mask_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTmain_mask_Int,
          Dcon ReadOut_CTmain_mask_Int) : (memReadOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) > [(readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf,CTmain_mask_Int)] */
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d = {memReadOut_CTmain_mask_Int_d[116:2],
                                                             memReadOut_CTmain_mask_Int_d[0]};
  assign memReadOut_CTmain_mask_Int_r = readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTmain_mask_Int) : [(lizzieLet15_1_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet24_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet36_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet37_1_argbuf,CTmain_mask_Int),
                                  (lizzieLet38_1_argbuf,CTmain_mask_Int)] > (writeMerge_choice_CTmain_mask_Int,C5) (writeMerge_data_CTmain_mask_Int,CTmain_mask_Int) */
  logic [4:0] lizzieLet15_1_1_argbuf_select_d;
  assign lizzieLet15_1_1_argbuf_select_d = ((| lizzieLet15_1_1_argbuf_select_q) ? lizzieLet15_1_1_argbuf_select_q :
                                            (lizzieLet15_1_1_argbuf_d[0] ? 5'd1 :
                                             (lizzieLet24_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet36_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet37_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet38_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] lizzieLet15_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet15_1_1_argbuf_select_q <= (lizzieLet15_1_1_argbuf_done ? 5'd0 :
                                          lizzieLet15_1_1_argbuf_select_d);
  logic [1:0] lizzieLet15_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet15_1_1_argbuf_emit_q <= (lizzieLet15_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet15_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet15_1_1_argbuf_emit_d;
  assign lizzieLet15_1_1_argbuf_emit_d = (lizzieLet15_1_1_argbuf_emit_q | ({writeMerge_choice_CTmain_mask_Int_d[0],
                                                                            writeMerge_data_CTmain_mask_Int_d[0]} & {writeMerge_choice_CTmain_mask_Int_r,
                                                                                                                     writeMerge_data_CTmain_mask_Int_r}));
  logic lizzieLet15_1_1_argbuf_done;
  assign lizzieLet15_1_1_argbuf_done = (& lizzieLet15_1_1_argbuf_emit_d);
  assign {lizzieLet38_1_argbuf_r,
          lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r} = (lizzieLet15_1_1_argbuf_done ? lizzieLet15_1_1_argbuf_select_d :
                                       5'd0);
  assign writeMerge_data_CTmain_mask_Int_d = ((lizzieLet15_1_1_argbuf_select_d[0] && (! lizzieLet15_1_1_argbuf_emit_q[0])) ? lizzieLet15_1_1_argbuf_d :
                                              ((lizzieLet15_1_1_argbuf_select_d[1] && (! lizzieLet15_1_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                               ((lizzieLet15_1_1_argbuf_select_d[2] && (! lizzieLet15_1_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                ((lizzieLet15_1_1_argbuf_select_d[3] && (! lizzieLet15_1_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                 ((lizzieLet15_1_1_argbuf_select_d[4] && (! lizzieLet15_1_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                                  {115'd0, 1'd0})))));
  assign writeMerge_choice_CTmain_mask_Int_d = ((lizzieLet15_1_1_argbuf_select_d[0] && (! lizzieLet15_1_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                ((lizzieLet15_1_1_argbuf_select_d[1] && (! lizzieLet15_1_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                 ((lizzieLet15_1_1_argbuf_select_d[2] && (! lizzieLet15_1_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                  ((lizzieLet15_1_1_argbuf_select_d[3] && (! lizzieLet15_1_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                   ((lizzieLet15_1_1_argbuf_select_d[4] && (! lizzieLet15_1_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                    {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_mask_Int) : (writeMerge_choice_CTmain_mask_Int,C5) (demuxWriteResult_CTmain_mask_Int,Pointer_CTmain_mask_Int) > [(writeCTmain_mask_IntlizzieLet15_1_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet24_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet36_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet37_1_argbuf,Pointer_CTmain_mask_Int),
                                                                                                                                          (writeCTmain_mask_IntlizzieLet38_1_argbuf,Pointer_CTmain_mask_Int)] */
  logic [4:0] demuxWriteResult_CTmain_mask_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTmain_mask_Int_d[0] && demuxWriteResult_CTmain_mask_Int_d[0]))
      unique case (writeMerge_choice_CTmain_mask_Int_d[3:1])
        3'd0: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTmain_mask_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTmain_mask_Int_onehotd = 5'd0;
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                         demuxWriteResult_CTmain_mask_Int_onehotd[0]};
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[1]};
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[2]};
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[3]};
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_d = {demuxWriteResult_CTmain_mask_Int_d[16:1],
                                                       demuxWriteResult_CTmain_mask_Int_onehotd[4]};
  assign demuxWriteResult_CTmain_mask_Int_r = (| (demuxWriteResult_CTmain_mask_Int_onehotd & {writeCTmain_mask_IntlizzieLet38_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet37_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet36_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet24_1_argbuf_r,
                                                                                              writeCTmain_mask_IntlizzieLet15_1_1_argbuf_r}));
  assign writeMerge_choice_CTmain_mask_Int_r = demuxWriteResult_CTmain_mask_Int_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Int,
      Dcon WriteIn_CTmain_mask_Int) : [(forkHP1_CTmain_mask_In2,Word16#),
                                       (writeMerge_data_CTmain_mask_Int,CTmain_mask_Int)] > (dconWriteIn_CTmain_mask_Int,MemIn_CTmain_mask_Int) */
  assign dconWriteIn_CTmain_mask_Int_d = WriteIn_CTmain_mask_Int_dc((& {forkHP1_CTmain_mask_In2_d[0],
                                                                        writeMerge_data_CTmain_mask_Int_d[0]}), forkHP1_CTmain_mask_In2_d, writeMerge_data_CTmain_mask_Int_d);
  assign {forkHP1_CTmain_mask_In2_r,
          writeMerge_data_CTmain_mask_Int_r} = {2 {(dconWriteIn_CTmain_mask_Int_r && dconWriteIn_CTmain_mask_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTmain_mask_Int,
      Dcon Pointer_CTmain_mask_Int) : [(forkHP1_CTmain_mask_In3,Word16#)] > (dconPtr_CTmain_mask_Int,Pointer_CTmain_mask_Int) */
  assign dconPtr_CTmain_mask_Int_d = Pointer_CTmain_mask_Int_dc((& {forkHP1_CTmain_mask_In3_d[0]}), forkHP1_CTmain_mask_In3_d);
  assign {forkHP1_CTmain_mask_In3_r} = {1 {(dconPtr_CTmain_mask_Int_r && dconPtr_CTmain_mask_Int_d[0])}};
  
  /* demux (Ty MemOut_CTmain_mask_Int,
       Ty Pointer_CTmain_mask_Int) : (memWriteOut_CTmain_mask_Int,MemOut_CTmain_mask_Int) (dconPtr_CTmain_mask_Int,Pointer_CTmain_mask_Int) > [(_52,Pointer_CTmain_mask_Int),
                                                                                                                                               (demuxWriteResult_CTmain_mask_Int,Pointer_CTmain_mask_Int)] */
  logic [1:0] dconPtr_CTmain_mask_Int_onehotd;
  always_comb
    if ((memWriteOut_CTmain_mask_Int_d[0] && dconPtr_CTmain_mask_Int_d[0]))
      unique case (memWriteOut_CTmain_mask_Int_d[1:1])
        1'd0: dconPtr_CTmain_mask_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTmain_mask_Int_onehotd = 2'd2;
        default: dconPtr_CTmain_mask_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTmain_mask_Int_onehotd = 2'd0;
  assign _52_d = {dconPtr_CTmain_mask_Int_d[16:1],
                  dconPtr_CTmain_mask_Int_onehotd[0]};
  assign demuxWriteResult_CTmain_mask_Int_d = {dconPtr_CTmain_mask_Int_d[16:1],
                                               dconPtr_CTmain_mask_Int_onehotd[1]};
  assign dconPtr_CTmain_mask_Int_r = (| (dconPtr_CTmain_mask_Int_onehotd & {demuxWriteResult_CTmain_mask_Int_r,
                                                                            _52_r}));
  assign memWriteOut_CTmain_mask_Int_r = dconPtr_CTmain_mask_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__10,Go) > (initHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \initHP_CTmap''_map''_Int_Int_Int_d  = {16'd0, go__10_d[0]};
  assign go__10_r = \initHP_CTmap''_map''_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmap''_map''_Int_Int_Int1,Go) > (incrHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \incrHP_CTmap''_map''_Int_Int_Int_d  = {16'd1,
                                                 \incrHP_CTmap''_map''_Int_Int_Int1_d [0]};
  assign \incrHP_CTmap''_map''_Int_Int_Int1_r  = \incrHP_CTmap''_map''_Int_Int_Int_r ;
  
  /* merge (Ty Go) : [(go__11,Go),
                 (incrHP_CTmap''_map''_Int_Int_Int2,Go)] > (incrHP_mergeCTmap''_map''_Int_Int_Int,Go) */
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_selected ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTmap''_map''_Int_Int_Int_select ))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  = \incrHP_mergeCTmap''_map''_Int_Int_Int_select ;
      else
        if (go__11_d[0])
          \incrHP_mergeCTmap''_map''_Int_Int_Int_selected [0] = 1'd1;
        else if (\incrHP_CTmap''_map''_Int_Int_Int2_d [0])
          \incrHP_mergeCTmap''_map''_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Int_Int_Int_select  <= (\incrHP_mergeCTmap''_map''_Int_Int_Int_r  ? 2'd0 :
                                                         \incrHP_mergeCTmap''_map''_Int_Int_Int_selected );
  always_comb
    if (\incrHP_mergeCTmap''_map''_Int_Int_Int_selected [0])
      \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = go__11_d;
    else if (\incrHP_mergeCTmap''_map''_Int_Int_Int_selected [1])
      \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = \incrHP_CTmap''_map''_Int_Int_Int2_d ;
    else \incrHP_mergeCTmap''_map''_Int_Int_Int_d  = 1'd0;
  assign {\incrHP_CTmap''_map''_Int_Int_Int2_r ,
          go__11_r} = (\incrHP_mergeCTmap''_map''_Int_Int_Int_r  ? \incrHP_mergeCTmap''_map''_Int_Int_Int_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmap''_map''_Int_Int_Int_buf,Go) > [(incrHP_CTmap''_map''_Int_Int_Int1,Go),
                                                                 (incrHP_CTmap''_map''_Int_Int_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done ;
  assign \incrHP_CTmap''_map''_Int_Int_Int1_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted [0]));
  assign \incrHP_CTmap''_map''_Int_Int_Int2_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted [1]));
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  | ({\incrHP_CTmap''_map''_Int_Int_Int2_d [0],
                                                                                                                     \incrHP_CTmap''_map''_Int_Int_Int1_d [0]} & {\incrHP_CTmap''_map''_Int_Int_Int2_r ,
                                                                                                                                                                  \incrHP_CTmap''_map''_Int_Int_Int1_r }));
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  = (& \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_emitted  <= (\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  ? 2'd0 :
                                                              \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmap''_map''_Int_Int_Int,Word16#) (forkHP1_CTmap''_map''_Int_Int_Int,Word16#) > (addHP_CTmap''_map''_Int_Int_Int,Word16#) */
  assign \addHP_CTmap''_map''_Int_Int_Int_d  = {(\incrHP_CTmap''_map''_Int_Int_Int_d [16:1] + \forkHP1_CTmap''_map''_Int_Int_Int_d [16:1]),
                                                (\incrHP_CTmap''_map''_Int_Int_Int_d [0] && \forkHP1_CTmap''_map''_Int_Int_Int_d [0])};
  assign {\incrHP_CTmap''_map''_Int_Int_Int_r ,
          \forkHP1_CTmap''_map''_Int_Int_Int_r } = {2 {(\addHP_CTmap''_map''_Int_Int_Int_r  && \addHP_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmap''_map''_Int_Int_Int,Word16#),
                      (addHP_CTmap''_map''_Int_Int_Int,Word16#)] > (mergeHP_CTmap''_map''_Int_Int_Int,Word16#) */
  logic [1:0] \mergeHP_CTmap''_map''_Int_Int_Int_selected ;
  logic [1:0] \mergeHP_CTmap''_map''_Int_Int_Int_select ;
  always_comb
    begin
      \mergeHP_CTmap''_map''_Int_Int_Int_selected  = 2'd0;
      if ((| \mergeHP_CTmap''_map''_Int_Int_Int_select ))
        \mergeHP_CTmap''_map''_Int_Int_Int_selected  = \mergeHP_CTmap''_map''_Int_Int_Int_select ;
      else
        if (\initHP_CTmap''_map''_Int_Int_Int_d [0])
          \mergeHP_CTmap''_map''_Int_Int_Int_selected [0] = 1'd1;
        else if (\addHP_CTmap''_map''_Int_Int_Int_d [0])
          \mergeHP_CTmap''_map''_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_select  <= 2'd0;
    else
      \mergeHP_CTmap''_map''_Int_Int_Int_select  <= (\mergeHP_CTmap''_map''_Int_Int_Int_r  ? 2'd0 :
                                                     \mergeHP_CTmap''_map''_Int_Int_Int_selected );
  always_comb
    if (\mergeHP_CTmap''_map''_Int_Int_Int_selected [0])
      \mergeHP_CTmap''_map''_Int_Int_Int_d  = \initHP_CTmap''_map''_Int_Int_Int_d ;
    else if (\mergeHP_CTmap''_map''_Int_Int_Int_selected [1])
      \mergeHP_CTmap''_map''_Int_Int_Int_d  = \addHP_CTmap''_map''_Int_Int_Int_d ;
    else \mergeHP_CTmap''_map''_Int_Int_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTmap''_map''_Int_Int_Int_r ,
          \initHP_CTmap''_map''_Int_Int_Int_r } = (\mergeHP_CTmap''_map''_Int_Int_Int_r  ? \mergeHP_CTmap''_map''_Int_Int_Int_selected  :
                                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmap''_map''_Int_Int_Int,Go) > (incrHP_mergeCTmap''_map''_Int_Int_Int_buf,Go) */
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d ;
  logic \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r ;
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_r  = ((! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d [0]) || \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmap''_map''_Int_Int_Int_r )
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d  <= \incrHP_mergeCTmap''_map''_Int_Int_Int_d ;
  Go_t \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf ;
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_r  = (! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_d  = (\incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0] ? \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  :
                                                          \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r  && \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0]))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmap''_map''_Int_Int_Int_buf_r ) && (! \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf [0])))
        \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_buf  <= \incrHP_mergeCTmap''_map''_Int_Int_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmap''_map''_Int_Int_Int,Word16#) > (mergeHP_CTmap''_map''_Int_Int_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d ;
  logic \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r ;
  assign \mergeHP_CTmap''_map''_Int_Int_Int_r  = ((! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d [0]) || \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmap''_map''_Int_Int_Int_r )
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d  <= \mergeHP_CTmap''_map''_Int_Int_Int_d ;
  \Word16#_t  \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf ;
  assign \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_r  = (! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0]);
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_d  = (\mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0] ? \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  :
                                                      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTmap''_map''_Int_Int_Int_buf_r  && \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0]))
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTmap''_map''_Int_Int_Int_buf_r ) && (! \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf [0])))
        \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_buf  <= \mergeHP_CTmap''_map''_Int_Int_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmap''_map''_Int_Int_Int_buf,Word16#) > [(forkHP1_CTmap''_map''_Int_Int_Int,Word16#),
                                                                       (forkHP1_CTmap''_map''_Int_Int_In2,Word16#),
                                                                       (forkHP1_CTmap''_map''_Int_Int_In3,Word16#)] */
  logic [2:0] \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTmap''_map''_Int_Int_Int_buf_done ;
  assign \forkHP1_CTmap''_map''_Int_Int_Int_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [0]))};
  assign \forkHP1_CTmap''_map''_Int_Int_In2_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [1]))};
  assign \forkHP1_CTmap''_map''_Int_Int_In3_d  = {\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [16:1],
                                                  (\mergeHP_CTmap''_map''_Int_Int_Int_buf_d [0] && (! \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted [2]))};
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_done  = (\mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  | ({\forkHP1_CTmap''_map''_Int_Int_In3_d [0],
                                                                                                             \forkHP1_CTmap''_map''_Int_Int_In2_d [0],
                                                                                                             \forkHP1_CTmap''_map''_Int_Int_Int_d [0]} & {\forkHP1_CTmap''_map''_Int_Int_In3_r ,
                                                                                                                                                          \forkHP1_CTmap''_map''_Int_Int_In2_r ,
                                                                                                                                                          \forkHP1_CTmap''_map''_Int_Int_Int_r }));
  assign \mergeHP_CTmap''_map''_Int_Int_Int_buf_r  = (& \mergeHP_CTmap''_map''_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmap''_map''_Int_Int_Int_buf_emitted  <= (\mergeHP_CTmap''_map''_Int_Int_Int_buf_r  ? 3'd0 :
                                                          \mergeHP_CTmap''_map''_Int_Int_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmap''_map''_Int_Int_Int) : [(dconReadIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int),
                                                  (dconWriteIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int)] > (memMergeChoice_CTmap''_map''_Int_Int_Int,C2) (memMergeIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_select_d ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_select_d  = ((| \dconReadIn_CTmap''_map''_Int_Int_Int_select_q ) ? \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  :
                                                            (\dconReadIn_CTmap''_map''_Int_Int_Int_d [0] ? 2'd1 :
                                                             (\dconWriteIn_CTmap''_map''_Int_Int_Int_d [0] ? 2'd2 :
                                                              2'd0)));
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Int_Int_Int_select_q  <= (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? 2'd0 :
                                                          \dconReadIn_CTmap''_map''_Int_Int_Int_select_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  <= (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? 2'd0 :
                                                        \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d  = (\dconReadIn_CTmap''_map''_Int_Int_Int_emit_q  | ({\memMergeChoice_CTmap''_map''_Int_Int_Int_d [0],
                                                                                                            \memMergeIn_CTmap''_map''_Int_Int_Int_d [0]} & {\memMergeChoice_CTmap''_map''_Int_Int_Int_r ,
                                                                                                                                                            \memMergeIn_CTmap''_map''_Int_Int_Int_r }));
  logic \dconReadIn_CTmap''_map''_Int_Int_Int_done ;
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_done  = (& \dconReadIn_CTmap''_map''_Int_Int_Int_emit_d );
  assign {\dconWriteIn_CTmap''_map''_Int_Int_Int_r ,
          \dconReadIn_CTmap''_map''_Int_Int_Int_r } = (\dconReadIn_CTmap''_map''_Int_Int_Int_done  ? \dconReadIn_CTmap''_map''_Int_Int_Int_select_d  :
                                                       2'd0);
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_d  = ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [0] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [0])) ? \dconReadIn_CTmap''_map''_Int_Int_Int_d  :
                                                     ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [1] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [0])) ? \dconWriteIn_CTmap''_map''_Int_Int_Int_d  :
                                                      {116'd0, 1'd0}));
  assign \memMergeChoice_CTmap''_map''_Int_Int_Int_d  = ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [0] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                         ((\dconReadIn_CTmap''_map''_Int_Int_Int_select_d [1] && (! \dconReadIn_CTmap''_map''_Int_Int_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Ty MemOut_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int_dbuf,MemIn_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) */
  logic [98:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ;
  logic [98:0] \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
  logic [98:0] \memOut_CTmap''_map''_Int_Int_Int_q ;
  logic \memOut_CTmap''_map''_Int_Int_Int_valid ;
  logic \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we ;
  logic \memOut_CTmap''_map''_Int_Int_Int_we ;
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din  = \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [116:18];
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address  = \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [17:2];
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we  = (\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [1:1] && \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmap''_map''_Int_Int_Int_we  <= 1'd0;
        \memOut_CTmap''_map''_Int_Int_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmap''_map''_Int_Int_Int_we  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we ;
        \memOut_CTmap''_map''_Int_Int_Int_valid  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0];
        if (\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we )
          begin
            \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ] <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
            \memOut_CTmap''_map''_Int_Int_Int_q  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_din ;
          end
        else
          \memOut_CTmap''_map''_Int_Int_Int_q  <= \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_mem [\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_address ];
      end
  assign \memOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_q ,
                                                 \memOut_CTmap''_map''_Int_Int_Int_we ,
                                                 \memOut_CTmap''_map''_Int_Int_Int_valid };
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r  = ((! \memOut_CTmap''_map''_Int_Int_Int_valid ) || \memOut_CTmap''_map''_Int_Int_Int_r );
  logic [31:0] \profiling_MemIn_CTmap''_map''_Int_Int_Int_read ;
  logic [31:0] \profiling_MemIn_CTmap''_map''_Int_Int_Int_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTmap''_map''_Int_Int_Int_write  <= 0;
        \profiling_MemIn_CTmap''_map''_Int_Int_Int_read  <= 0;
      end
    else
      if ((\memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_we  == 1'd1))
        \profiling_MemIn_CTmap''_map''_Int_Int_Int_write  <= (\profiling_MemIn_CTmap''_map''_Int_Int_Int_write  + 1);
      else
        if ((\memOut_CTmap''_map''_Int_Int_Int_valid  == 1'd1))
          \profiling_MemIn_CTmap''_map''_Int_Int_Int_read  <= (\profiling_MemIn_CTmap''_map''_Int_Int_Int_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmap''_map''_Int_Int_Int) : (memMergeChoice_CTmap''_map''_Int_Int_Int,C2) (memOut_CTmap''_map''_Int_Int_Int_dbuf,MemOut_CTmap''_map''_Int_Int_Int) > [(memReadOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                        (memWriteOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmap''_map''_Int_Int_Int_d [0] && \memOut_CTmap''_map''_Int_Int_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTmap''_map''_Int_Int_Int_d [1:1])
        1'd0: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_dbuf_d [100:1],
                                                     \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTmap''_map''_Int_Int_Int_d  = {\memOut_CTmap''_map''_Int_Int_Int_dbuf_d [100:1],
                                                      \memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd [1]};
  assign \memOut_CTmap''_map''_Int_Int_Int_dbuf_r  = (| (\memOut_CTmap''_map''_Int_Int_Int_dbuf_onehotd  & {\memWriteOut_CTmap''_map''_Int_Int_Int_r ,
                                                                                                            \memReadOut_CTmap''_map''_Int_Int_Int_r }));
  assign \memMergeChoice_CTmap''_map''_Int_Int_Int_r  = \memOut_CTmap''_map''_Int_Int_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int_rbuf,MemIn_CTmap''_map''_Int_Int_Int) > (memMergeIn_CTmap''_map''_Int_Int_Int_dbuf,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r  = ((! \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d [0]) || \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r )
        \memMergeIn_CTmap''_map''_Int_Int_Int_dbuf_d  <= \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmap''_map''_Int_Int_Int) : (memMergeIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) > (memMergeIn_CTmap''_map''_Int_Int_Int_rbuf,MemIn_CTmap''_map''_Int_Int_Int) */
  \MemIn_CTmap''_map''_Int_Int_Int_t  \memMergeIn_CTmap''_map''_Int_Int_Int_buf ;
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_r  = (! \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0]);
  assign \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_d  = (\memMergeIn_CTmap''_map''_Int_Int_Int_buf [0] ? \memMergeIn_CTmap''_map''_Int_Int_Int_buf  :
                                                          \memMergeIn_CTmap''_map''_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r  && \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0]))
        \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memMergeIn_CTmap''_map''_Int_Int_Int_rbuf_r ) && (! \memMergeIn_CTmap''_map''_Int_Int_Int_buf [0])))
        \memMergeIn_CTmap''_map''_Int_Int_Int_buf  <= \memMergeIn_CTmap''_map''_Int_Int_Int_d ;
  
  /* dbuf (Ty MemOut_CTmap''_map''_Int_Int_Int) : (memOut_CTmap''_map''_Int_Int_Int_rbuf,MemOut_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int_dbuf,MemOut_CTmap''_map''_Int_Int_Int) */
  assign \memOut_CTmap''_map''_Int_Int_Int_rbuf_r  = ((! \memOut_CTmap''_map''_Int_Int_Int_dbuf_d [0]) || \memOut_CTmap''_map''_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Int_Int_Int_dbuf_d  <= {100'd0, 1'd0};
    else
      if (\memOut_CTmap''_map''_Int_Int_Int_rbuf_r )
        \memOut_CTmap''_map''_Int_Int_Int_dbuf_d  <= \memOut_CTmap''_map''_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmap''_map''_Int_Int_Int) : (memOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) > (memOut_CTmap''_map''_Int_Int_Int_rbuf,MemOut_CTmap''_map''_Int_Int_Int) */
  \MemOut_CTmap''_map''_Int_Int_Int_t  \memOut_CTmap''_map''_Int_Int_Int_buf ;
  assign \memOut_CTmap''_map''_Int_Int_Int_r  = (! \memOut_CTmap''_map''_Int_Int_Int_buf [0]);
  assign \memOut_CTmap''_map''_Int_Int_Int_rbuf_d  = (\memOut_CTmap''_map''_Int_Int_Int_buf [0] ? \memOut_CTmap''_map''_Int_Int_Int_buf  :
                                                      \memOut_CTmap''_map''_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Int_Int_Int_buf  <= {100'd0, 1'd0};
    else
      if ((\memOut_CTmap''_map''_Int_Int_Int_rbuf_r  && \memOut_CTmap''_map''_Int_Int_Int_buf [0]))
        \memOut_CTmap''_map''_Int_Int_Int_buf  <= {100'd0, 1'd0};
      else if (((! \memOut_CTmap''_map''_Int_Int_Int_rbuf_r ) && (! \memOut_CTmap''_map''_Int_Int_Int_buf [0])))
        \memOut_CTmap''_map''_Int_Int_Int_buf  <= \memOut_CTmap''_map''_Int_Int_Int_d ;
  
  /* destruct (Ty Pointer_CTmap''_map''_Int_Int_Int,
          Dcon Pointer_CTmap''_map''_Int_Int_Int) : (scfarg_0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > [(destructReadIn_CTmap''_map''_Int_Int_Int,Word16#)] */
  assign \destructReadIn_CTmap''_map''_Int_Int_Int_d  = {scfarg_0_3_1_argbuf_d[16:1],
                                                         scfarg_0_3_1_argbuf_d[0]};
  assign scfarg_0_3_1_argbuf_r = \destructReadIn_CTmap''_map''_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Dcon ReadIn_CTmap''_map''_Int_Int_Int) : [(destructReadIn_CTmap''_map''_Int_Int_Int,Word16#)] > (dconReadIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \dconReadIn_CTmap''_map''_Int_Int_Int_d  = \ReadIn_CTmap''_map''_Int_Int_Int_dc ((& {\destructReadIn_CTmap''_map''_Int_Int_Int_d [0]}), \destructReadIn_CTmap''_map''_Int_Int_Int_d );
  assign {\destructReadIn_CTmap''_map''_Int_Int_Int_r } = {1 {(\dconReadIn_CTmap''_map''_Int_Int_Int_r  && \dconReadIn_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTmap''_map''_Int_Int_Int,
          Dcon ReadOut_CTmap''_map''_Int_Int_Int) : (memReadOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) > [(readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf,CTmap''_map''_Int_Int_Int)] */
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d  = {\memReadOut_CTmap''_map''_Int_Int_Int_d [100:2],
                                                                         \memReadOut_CTmap''_map''_Int_Int_Int_d [0]};
  assign \memReadOut_CTmap''_map''_Int_Int_Int_r  = \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmap''_map''_Int_Int_Int) : [(lizzieLet21_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet25_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet41_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet42_1_argbuf,CTmap''_map''_Int_Int_Int),
                                            (lizzieLet43_1_argbuf,CTmap''_map''_Int_Int_Int)] > (writeMerge_choice_CTmap''_map''_Int_Int_Int,C5) (writeMerge_data_CTmap''_map''_Int_Int_Int,CTmap''_map''_Int_Int_Int) */
  logic [4:0] lizzieLet21_1_argbuf_select_d;
  assign lizzieLet21_1_argbuf_select_d = ((| lizzieLet21_1_argbuf_select_q) ? lizzieLet21_1_argbuf_select_q :
                                          (lizzieLet21_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet25_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet41_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet42_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet43_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet21_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet21_1_argbuf_select_q <= (lizzieLet21_1_argbuf_done ? 5'd0 :
                                        lizzieLet21_1_argbuf_select_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet21_1_argbuf_emit_q <= (lizzieLet21_1_argbuf_done ? 2'd0 :
                                      lizzieLet21_1_argbuf_emit_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_d;
  assign lizzieLet21_1_argbuf_emit_d = (lizzieLet21_1_argbuf_emit_q | ({\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [0],
                                                                        \writeMerge_data_CTmap''_map''_Int_Int_Int_d [0]} & {\writeMerge_choice_CTmap''_map''_Int_Int_Int_r ,
                                                                                                                             \writeMerge_data_CTmap''_map''_Int_Int_Int_r }));
  logic lizzieLet21_1_argbuf_done;
  assign lizzieLet21_1_argbuf_done = (& lizzieLet21_1_argbuf_emit_d);
  assign {lizzieLet43_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet21_1_argbuf_r} = (lizzieLet21_1_argbuf_done ? lizzieLet21_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmap''_map''_Int_Int_Int_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                                          ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                           ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                            ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                             ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                                              {99'd0, 1'd0})))));
  assign \writeMerge_choice_CTmap''_map''_Int_Int_Int_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                            ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                             ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                              ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                               ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeMerge_choice_CTmap''_map''_Int_Int_Int,C5) (demuxWriteResult_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                  (writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [4:0] \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [0] && \demuxWriteResult_CTmap''_map''_Int_Int_Int_d [0]))
      unique case (\writeMerge_choice_CTmap''_map''_Int_Int_Int_d [3:1])
        3'd0: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  = 5'd0;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [0]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [1]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [2]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [3]};
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd [4]};
  assign \demuxWriteResult_CTmap''_map''_Int_Int_Int_r  = (| (\demuxWriteResult_CTmap''_map''_Int_Int_Int_onehotd  & {\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_r ,
                                                                                                                      \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_r }));
  assign \writeMerge_choice_CTmap''_map''_Int_Int_Int_r  = \demuxWriteResult_CTmap''_map''_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Int_Int_Int,
      Dcon WriteIn_CTmap''_map''_Int_Int_Int) : [(forkHP1_CTmap''_map''_Int_Int_In2,Word16#),
                                                 (writeMerge_data_CTmap''_map''_Int_Int_Int,CTmap''_map''_Int_Int_Int)] > (dconWriteIn_CTmap''_map''_Int_Int_Int,MemIn_CTmap''_map''_Int_Int_Int) */
  assign \dconWriteIn_CTmap''_map''_Int_Int_Int_d  = \WriteIn_CTmap''_map''_Int_Int_Int_dc ((& {\forkHP1_CTmap''_map''_Int_Int_In2_d [0],
                                                                                                \writeMerge_data_CTmap''_map''_Int_Int_Int_d [0]}), \forkHP1_CTmap''_map''_Int_Int_In2_d , \writeMerge_data_CTmap''_map''_Int_Int_Int_d );
  assign {\forkHP1_CTmap''_map''_Int_Int_In2_r ,
          \writeMerge_data_CTmap''_map''_Int_Int_Int_r } = {2 {(\dconWriteIn_CTmap''_map''_Int_Int_Int_r  && \dconWriteIn_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTmap''_map''_Int_Int_Int,
      Dcon Pointer_CTmap''_map''_Int_Int_Int) : [(forkHP1_CTmap''_map''_Int_Int_In3,Word16#)] > (dconPtr_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) */
  assign \dconPtr_CTmap''_map''_Int_Int_Int_d  = \Pointer_CTmap''_map''_Int_Int_Int_dc ((& {\forkHP1_CTmap''_map''_Int_Int_In3_d [0]}), \forkHP1_CTmap''_map''_Int_Int_In3_d );
  assign {\forkHP1_CTmap''_map''_Int_Int_In3_r } = {1 {(\dconPtr_CTmap''_map''_Int_Int_Int_r  && \dconPtr_CTmap''_map''_Int_Int_Int_d [0])}};
  
  /* demux (Ty MemOut_CTmap''_map''_Int_Int_Int,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (memWriteOut_CTmap''_map''_Int_Int_Int,MemOut_CTmap''_map''_Int_Int_Int) (dconPtr_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(_51,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                                                                                 (demuxWriteResult_CTmap''_map''_Int_Int_Int,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] \dconPtr_CTmap''_map''_Int_Int_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTmap''_map''_Int_Int_Int_d [0] && \dconPtr_CTmap''_map''_Int_Int_Int_d [0]))
      unique case (\memWriteOut_CTmap''_map''_Int_Int_Int_d [1:1])
        1'd0: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd2;
        default: \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmap''_map''_Int_Int_Int_onehotd  = 2'd0;
  assign _51_d = {\dconPtr_CTmap''_map''_Int_Int_Int_d [16:1],
                  \dconPtr_CTmap''_map''_Int_Int_Int_onehotd [0]};
  assign \demuxWriteResult_CTmap''_map''_Int_Int_Int_d  = {\dconPtr_CTmap''_map''_Int_Int_Int_d [16:1],
                                                           \dconPtr_CTmap''_map''_Int_Int_Int_onehotd [1]};
  assign \dconPtr_CTmap''_map''_Int_Int_Int_r  = (| (\dconPtr_CTmap''_map''_Int_Int_Int_onehotd  & {\demuxWriteResult_CTmap''_map''_Int_Int_Int_r ,
                                                                                                    _51_r}));
  assign \memWriteOut_CTmap''_map''_Int_Int_Int_r  = \dconPtr_CTmap''_map''_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go__12,Go) > (initHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign initHP_CTkron_kron_Int_Int_Int_d = {16'd0, go__12_d[0]};
  assign go__12_r = initHP_CTkron_kron_Int_Int_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTkron_kron_Int_Int_Int1,Go) > (incrHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign incrHP_CTkron_kron_Int_Int_Int_d = {16'd1,
                                             incrHP_CTkron_kron_Int_Int_Int1_d[0]};
  assign incrHP_CTkron_kron_Int_Int_Int1_r = incrHP_CTkron_kron_Int_Int_Int_r;
  
  /* merge (Ty Go) : [(go__13,Go),
                 (incrHP_CTkron_kron_Int_Int_Int2,Go)] > (incrHP_mergeCTkron_kron_Int_Int_Int,Go) */
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_selected;
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_select;
  always_comb
    begin
      incrHP_mergeCTkron_kron_Int_Int_Int_selected = 2'd0;
      if ((| incrHP_mergeCTkron_kron_Int_Int_Int_select))
        incrHP_mergeCTkron_kron_Int_Int_Int_selected = incrHP_mergeCTkron_kron_Int_Int_Int_select;
      else
        if (go__13_d[0])
          incrHP_mergeCTkron_kron_Int_Int_Int_selected[0] = 1'd1;
        else if (incrHP_CTkron_kron_Int_Int_Int2_d[0])
          incrHP_mergeCTkron_kron_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_select <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Int_Int_Int_select <= (incrHP_mergeCTkron_kron_Int_Int_Int_r ? 2'd0 :
                                                     incrHP_mergeCTkron_kron_Int_Int_Int_selected);
  always_comb
    if (incrHP_mergeCTkron_kron_Int_Int_Int_selected[0])
      incrHP_mergeCTkron_kron_Int_Int_Int_d = go__13_d;
    else if (incrHP_mergeCTkron_kron_Int_Int_Int_selected[1])
      incrHP_mergeCTkron_kron_Int_Int_Int_d = incrHP_CTkron_kron_Int_Int_Int2_d;
    else incrHP_mergeCTkron_kron_Int_Int_Int_d = 1'd0;
  assign {incrHP_CTkron_kron_Int_Int_Int2_r,
          go__13_r} = (incrHP_mergeCTkron_kron_Int_Int_Int_r ? incrHP_mergeCTkron_kron_Int_Int_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTkron_kron_Int_Int_Int_buf,Go) > [(incrHP_CTkron_kron_Int_Int_Int1,Go),
                                                               (incrHP_CTkron_kron_Int_Int_Int2,Go)] */
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTkron_kron_Int_Int_Int_buf_done;
  assign incrHP_CTkron_kron_Int_Int_Int1_d = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted[0]));
  assign incrHP_CTkron_kron_Int_Int_Int2_d = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted[1]));
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_done = (incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted | ({incrHP_CTkron_kron_Int_Int_Int2_d[0],
                                                                                                             incrHP_CTkron_kron_Int_Int_Int1_d[0]} & {incrHP_CTkron_kron_Int_Int_Int2_r,
                                                                                                                                                      incrHP_CTkron_kron_Int_Int_Int1_r}));
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_r = (& incrHP_mergeCTkron_kron_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Int_Int_Int_buf_emitted <= (incrHP_mergeCTkron_kron_Int_Int_Int_buf_r ? 2'd0 :
                                                          incrHP_mergeCTkron_kron_Int_Int_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTkron_kron_Int_Int_Int,Word16#) (forkHP1_CTkron_kron_Int_Int_Int,Word16#) > (addHP_CTkron_kron_Int_Int_Int,Word16#) */
  assign addHP_CTkron_kron_Int_Int_Int_d = {(incrHP_CTkron_kron_Int_Int_Int_d[16:1] + forkHP1_CTkron_kron_Int_Int_Int_d[16:1]),
                                            (incrHP_CTkron_kron_Int_Int_Int_d[0] && forkHP1_CTkron_kron_Int_Int_Int_d[0])};
  assign {incrHP_CTkron_kron_Int_Int_Int_r,
          forkHP1_CTkron_kron_Int_Int_Int_r} = {2 {(addHP_CTkron_kron_Int_Int_Int_r && addHP_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTkron_kron_Int_Int_Int,Word16#),
                      (addHP_CTkron_kron_Int_Int_Int,Word16#)] > (mergeHP_CTkron_kron_Int_Int_Int,Word16#) */
  logic [1:0] mergeHP_CTkron_kron_Int_Int_Int_selected;
  logic [1:0] mergeHP_CTkron_kron_Int_Int_Int_select;
  always_comb
    begin
      mergeHP_CTkron_kron_Int_Int_Int_selected = 2'd0;
      if ((| mergeHP_CTkron_kron_Int_Int_Int_select))
        mergeHP_CTkron_kron_Int_Int_Int_selected = mergeHP_CTkron_kron_Int_Int_Int_select;
      else
        if (initHP_CTkron_kron_Int_Int_Int_d[0])
          mergeHP_CTkron_kron_Int_Int_Int_selected[0] = 1'd1;
        else if (addHP_CTkron_kron_Int_Int_Int_d[0])
          mergeHP_CTkron_kron_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_select <= 2'd0;
    else
      mergeHP_CTkron_kron_Int_Int_Int_select <= (mergeHP_CTkron_kron_Int_Int_Int_r ? 2'd0 :
                                                 mergeHP_CTkron_kron_Int_Int_Int_selected);
  always_comb
    if (mergeHP_CTkron_kron_Int_Int_Int_selected[0])
      mergeHP_CTkron_kron_Int_Int_Int_d = initHP_CTkron_kron_Int_Int_Int_d;
    else if (mergeHP_CTkron_kron_Int_Int_Int_selected[1])
      mergeHP_CTkron_kron_Int_Int_Int_d = addHP_CTkron_kron_Int_Int_Int_d;
    else mergeHP_CTkron_kron_Int_Int_Int_d = {16'd0, 1'd0};
  assign {addHP_CTkron_kron_Int_Int_Int_r,
          initHP_CTkron_kron_Int_Int_Int_r} = (mergeHP_CTkron_kron_Int_Int_Int_r ? mergeHP_CTkron_kron_Int_Int_Int_selected :
                                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTkron_kron_Int_Int_Int,Go) > (incrHP_mergeCTkron_kron_Int_Int_Int_buf,Go) */
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d;
  logic incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r;
  assign incrHP_mergeCTkron_kron_Int_Int_Int_r = ((! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d[0]) || incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTkron_kron_Int_Int_Int_r)
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d <= incrHP_mergeCTkron_kron_Int_Int_Int_d;
  Go_t incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf;
  assign incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_r = (! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0]);
  assign incrHP_mergeCTkron_kron_Int_Int_Int_buf_d = (incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0] ? incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf :
                                                      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTkron_kron_Int_Int_Int_buf_r && incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0]))
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTkron_kron_Int_Int_Int_buf_r) && (! incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf[0])))
        incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_buf <= incrHP_mergeCTkron_kron_Int_Int_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTkron_kron_Int_Int_Int,Word16#) > (mergeHP_CTkron_kron_Int_Int_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_bufchan_d;
  logic mergeHP_CTkron_kron_Int_Int_Int_bufchan_r;
  assign mergeHP_CTkron_kron_Int_Int_Int_r = ((! mergeHP_CTkron_kron_Int_Int_Int_bufchan_d[0]) || mergeHP_CTkron_kron_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTkron_kron_Int_Int_Int_r)
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_d <= mergeHP_CTkron_kron_Int_Int_Int_d;
  \Word16#_t  mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf;
  assign mergeHP_CTkron_kron_Int_Int_Int_bufchan_r = (! mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0]);
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_d = (mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0] ? mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf :
                                                  mergeHP_CTkron_kron_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTkron_kron_Int_Int_Int_buf_r && mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0]))
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTkron_kron_Int_Int_Int_buf_r) && (! mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf[0])))
        mergeHP_CTkron_kron_Int_Int_Int_bufchan_buf <= mergeHP_CTkron_kron_Int_Int_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTkron_kron_Int_Int_Int_buf,Word16#) > [(forkHP1_CTkron_kron_Int_Int_Int,Word16#),
                                                                     (forkHP1_CTkron_kron_Int_Int_In2,Word16#),
                                                                     (forkHP1_CTkron_kron_Int_Int_In3,Word16#)] */
  logic [2:0] mergeHP_CTkron_kron_Int_Int_Int_buf_emitted;
  logic [2:0] mergeHP_CTkron_kron_Int_Int_Int_buf_done;
  assign forkHP1_CTkron_kron_Int_Int_Int_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[0]))};
  assign forkHP1_CTkron_kron_Int_Int_In2_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[1]))};
  assign forkHP1_CTkron_kron_Int_Int_In3_d = {mergeHP_CTkron_kron_Int_Int_Int_buf_d[16:1],
                                              (mergeHP_CTkron_kron_Int_Int_Int_buf_d[0] && (! mergeHP_CTkron_kron_Int_Int_Int_buf_emitted[2]))};
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_done = (mergeHP_CTkron_kron_Int_Int_Int_buf_emitted | ({forkHP1_CTkron_kron_Int_Int_In3_d[0],
                                                                                                     forkHP1_CTkron_kron_Int_Int_In2_d[0],
                                                                                                     forkHP1_CTkron_kron_Int_Int_Int_d[0]} & {forkHP1_CTkron_kron_Int_Int_In3_r,
                                                                                                                                              forkHP1_CTkron_kron_Int_Int_In2_r,
                                                                                                                                              forkHP1_CTkron_kron_Int_Int_Int_r}));
  assign mergeHP_CTkron_kron_Int_Int_Int_buf_r = (& mergeHP_CTkron_kron_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Int_Int_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTkron_kron_Int_Int_Int_buf_emitted <= (mergeHP_CTkron_kron_Int_Int_Int_buf_r ? 3'd0 :
                                                      mergeHP_CTkron_kron_Int_Int_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTkron_kron_Int_Int_Int) : [(dconReadIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int),
                                                (dconWriteIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int)] > (memMergeChoice_CTkron_kron_Int_Int_Int,C2) (memMergeIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_select_d;
  assign dconReadIn_CTkron_kron_Int_Int_Int_select_d = ((| dconReadIn_CTkron_kron_Int_Int_Int_select_q) ? dconReadIn_CTkron_kron_Int_Int_Int_select_q :
                                                        (dconReadIn_CTkron_kron_Int_Int_Int_d[0] ? 2'd1 :
                                                         (dconWriteIn_CTkron_kron_Int_Int_Int_d[0] ? 2'd2 :
                                                          2'd0)));
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Int_Int_Int_select_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Int_Int_Int_select_q <= (dconReadIn_CTkron_kron_Int_Int_Int_done ? 2'd0 :
                                                      dconReadIn_CTkron_kron_Int_Int_Int_select_d);
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Int_Int_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Int_Int_Int_emit_q <= (dconReadIn_CTkron_kron_Int_Int_Int_done ? 2'd0 :
                                                    dconReadIn_CTkron_kron_Int_Int_Int_emit_d);
  logic [1:0] dconReadIn_CTkron_kron_Int_Int_Int_emit_d;
  assign dconReadIn_CTkron_kron_Int_Int_Int_emit_d = (dconReadIn_CTkron_kron_Int_Int_Int_emit_q | ({memMergeChoice_CTkron_kron_Int_Int_Int_d[0],
                                                                                                    memMergeIn_CTkron_kron_Int_Int_Int_d[0]} & {memMergeChoice_CTkron_kron_Int_Int_Int_r,
                                                                                                                                                memMergeIn_CTkron_kron_Int_Int_Int_r}));
  logic dconReadIn_CTkron_kron_Int_Int_Int_done;
  assign dconReadIn_CTkron_kron_Int_Int_Int_done = (& dconReadIn_CTkron_kron_Int_Int_Int_emit_d);
  assign {dconWriteIn_CTkron_kron_Int_Int_Int_r,
          dconReadIn_CTkron_kron_Int_Int_Int_r} = (dconReadIn_CTkron_kron_Int_Int_Int_done ? dconReadIn_CTkron_kron_Int_Int_Int_select_d :
                                                   2'd0);
  assign memMergeIn_CTkron_kron_Int_Int_Int_d = ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[0] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[0])) ? dconReadIn_CTkron_kron_Int_Int_Int_d :
                                                 ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[1] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[0])) ? dconWriteIn_CTkron_kron_Int_Int_Int_d :
                                                  {100'd0, 1'd0}));
  assign memMergeChoice_CTkron_kron_Int_Int_Int_d = ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[0] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                                     ((dconReadIn_CTkron_kron_Int_Int_Int_select_d[1] && (! dconReadIn_CTkron_kron_Int_Int_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTkron_kron_Int_Int_Int,
      Ty MemOut_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int_dbuf,MemIn_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) */
  logic [82:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address;
  logic [82:0] memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
  logic [82:0] memOut_CTkron_kron_Int_Int_Int_q;
  logic memOut_CTkron_kron_Int_Int_Int_valid;
  logic memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we;
  logic memOut_CTkron_kron_Int_Int_Int_we;
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din = memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[100:18];
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address = memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[17:2];
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we = (memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[1:1] && memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTkron_kron_Int_Int_Int_we <= 1'd0;
        memOut_CTkron_kron_Int_Int_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTkron_kron_Int_Int_Int_we <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we;
        memOut_CTkron_kron_Int_Int_Int_valid <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0];
        if (memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we)
          begin
            memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address] <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
            memOut_CTkron_kron_Int_Int_Int_q <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_din;
          end
        else
          memOut_CTkron_kron_Int_Int_Int_q <= memMergeIn_CTkron_kron_Int_Int_Int_dbuf_mem[memMergeIn_CTkron_kron_Int_Int_Int_dbuf_address];
      end
  assign memOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_q,
                                             memOut_CTkron_kron_Int_Int_Int_we,
                                             memOut_CTkron_kron_Int_Int_Int_valid};
  assign memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r = ((! memOut_CTkron_kron_Int_Int_Int_valid) || memOut_CTkron_kron_Int_Int_Int_r);
  logic [31:0] profiling_MemIn_CTkron_kron_Int_Int_Int_read;
  logic [31:0] profiling_MemIn_CTkron_kron_Int_Int_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTkron_kron_Int_Int_Int_write <= 0;
        profiling_MemIn_CTkron_kron_Int_Int_Int_read <= 0;
      end
    else
      if ((memMergeIn_CTkron_kron_Int_Int_Int_dbuf_we == 1'd1))
        profiling_MemIn_CTkron_kron_Int_Int_Int_write <= (profiling_MemIn_CTkron_kron_Int_Int_Int_write + 1);
      else
        if ((memOut_CTkron_kron_Int_Int_Int_valid == 1'd1))
          profiling_MemIn_CTkron_kron_Int_Int_Int_read <= (profiling_MemIn_CTkron_kron_Int_Int_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTkron_kron_Int_Int_Int) : (memMergeChoice_CTkron_kron_Int_Int_Int,C2) (memOut_CTkron_kron_Int_Int_Int_dbuf,MemOut_CTkron_kron_Int_Int_Int) > [(memReadOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int),
                                                                                                                                                                (memWriteOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int)] */
  logic [1:0] memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTkron_kron_Int_Int_Int_d[0] && memOut_CTkron_kron_Int_Int_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTkron_kron_Int_Int_Int_d[1:1])
        1'd0: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_dbuf_d[84:1],
                                                 memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTkron_kron_Int_Int_Int_d = {memOut_CTkron_kron_Int_Int_Int_dbuf_d[84:1],
                                                  memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd[1]};
  assign memOut_CTkron_kron_Int_Int_Int_dbuf_r = (| (memOut_CTkron_kron_Int_Int_Int_dbuf_onehotd & {memWriteOut_CTkron_kron_Int_Int_Int_r,
                                                                                                    memReadOut_CTkron_kron_Int_Int_Int_r}));
  assign memMergeChoice_CTkron_kron_Int_Int_Int_r = memOut_CTkron_kron_Int_Int_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int_rbuf,MemIn_CTkron_kron_Int_Int_Int) > (memMergeIn_CTkron_kron_Int_Int_Int_dbuf,MemIn_CTkron_kron_Int_Int_Int) */
  assign memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r = ((! memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d[0]) || memMergeIn_CTkron_kron_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d <= {100'd0, 1'd0};
    else
      if (memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r)
        memMergeIn_CTkron_kron_Int_Int_Int_dbuf_d <= memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTkron_kron_Int_Int_Int) : (memMergeIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) > (memMergeIn_CTkron_kron_Int_Int_Int_rbuf,MemIn_CTkron_kron_Int_Int_Int) */
  MemIn_CTkron_kron_Int_Int_Int_t memMergeIn_CTkron_kron_Int_Int_Int_buf;
  assign memMergeIn_CTkron_kron_Int_Int_Int_r = (! memMergeIn_CTkron_kron_Int_Int_Int_buf[0]);
  assign memMergeIn_CTkron_kron_Int_Int_Int_rbuf_d = (memMergeIn_CTkron_kron_Int_Int_Int_buf[0] ? memMergeIn_CTkron_kron_Int_Int_Int_buf :
                                                      memMergeIn_CTkron_kron_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Int_Int_Int_buf <= {100'd0, 1'd0};
    else
      if ((memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r && memMergeIn_CTkron_kron_Int_Int_Int_buf[0]))
        memMergeIn_CTkron_kron_Int_Int_Int_buf <= {100'd0, 1'd0};
      else if (((! memMergeIn_CTkron_kron_Int_Int_Int_rbuf_r) && (! memMergeIn_CTkron_kron_Int_Int_Int_buf[0])))
        memMergeIn_CTkron_kron_Int_Int_Int_buf <= memMergeIn_CTkron_kron_Int_Int_Int_d;
  
  /* dbuf (Ty MemOut_CTkron_kron_Int_Int_Int) : (memOut_CTkron_kron_Int_Int_Int_rbuf,MemOut_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int_dbuf,MemOut_CTkron_kron_Int_Int_Int) */
  assign memOut_CTkron_kron_Int_Int_Int_rbuf_r = ((! memOut_CTkron_kron_Int_Int_Int_dbuf_d[0]) || memOut_CTkron_kron_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Int_Int_Int_dbuf_d <= {84'd0, 1'd0};
    else
      if (memOut_CTkron_kron_Int_Int_Int_rbuf_r)
        memOut_CTkron_kron_Int_Int_Int_dbuf_d <= memOut_CTkron_kron_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTkron_kron_Int_Int_Int) : (memOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) > (memOut_CTkron_kron_Int_Int_Int_rbuf,MemOut_CTkron_kron_Int_Int_Int) */
  MemOut_CTkron_kron_Int_Int_Int_t memOut_CTkron_kron_Int_Int_Int_buf;
  assign memOut_CTkron_kron_Int_Int_Int_r = (! memOut_CTkron_kron_Int_Int_Int_buf[0]);
  assign memOut_CTkron_kron_Int_Int_Int_rbuf_d = (memOut_CTkron_kron_Int_Int_Int_buf[0] ? memOut_CTkron_kron_Int_Int_Int_buf :
                                                  memOut_CTkron_kron_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Int_Int_Int_buf <= {84'd0, 1'd0};
    else
      if ((memOut_CTkron_kron_Int_Int_Int_rbuf_r && memOut_CTkron_kron_Int_Int_Int_buf[0]))
        memOut_CTkron_kron_Int_Int_Int_buf <= {84'd0, 1'd0};
      else if (((! memOut_CTkron_kron_Int_Int_Int_rbuf_r) && (! memOut_CTkron_kron_Int_Int_Int_buf[0])))
        memOut_CTkron_kron_Int_Int_Int_buf <= memOut_CTkron_kron_Int_Int_Int_d;
  
  /* destruct (Ty Pointer_CTkron_kron_Int_Int_Int,
          Dcon Pointer_CTkron_kron_Int_Int_Int) : (scfarg_0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > [(destructReadIn_CTkron_kron_Int_Int_Int,Word16#)] */
  assign destructReadIn_CTkron_kron_Int_Int_Int_d = {scfarg_0_1_1_argbuf_d[16:1],
                                                     scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CTkron_kron_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Int_Int_Int,
      Dcon ReadIn_CTkron_kron_Int_Int_Int) : [(destructReadIn_CTkron_kron_Int_Int_Int,Word16#)] > (dconReadIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  assign dconReadIn_CTkron_kron_Int_Int_Int_d = ReadIn_CTkron_kron_Int_Int_Int_dc((& {destructReadIn_CTkron_kron_Int_Int_Int_d[0]}), destructReadIn_CTkron_kron_Int_Int_Int_d);
  assign {destructReadIn_CTkron_kron_Int_Int_Int_r} = {1 {(dconReadIn_CTkron_kron_Int_Int_Int_r && dconReadIn_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTkron_kron_Int_Int_Int,
          Dcon ReadOut_CTkron_kron_Int_Int_Int) : (memReadOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) > [(readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf,CTkron_kron_Int_Int_Int)] */
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d = {memReadOut_CTkron_kron_Int_Int_Int_d[84:2],
                                                                     memReadOut_CTkron_kron_Int_Int_Int_d[0]};
  assign memReadOut_CTkron_kron_Int_Int_Int_r = readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTkron_kron_Int_Int_Int) : [(lizzieLet23_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet31_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet32_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet33_1_argbuf,CTkron_kron_Int_Int_Int),
                                          (lizzieLet8_1_argbuf,CTkron_kron_Int_Int_Int)] > (writeMerge_choice_CTkron_kron_Int_Int_Int,C5) (writeMerge_data_CTkron_kron_Int_Int_Int,CTkron_kron_Int_Int_Int) */
  logic [4:0] lizzieLet23_1_argbuf_select_d;
  assign lizzieLet23_1_argbuf_select_d = ((| lizzieLet23_1_argbuf_select_q) ? lizzieLet23_1_argbuf_select_q :
                                          (lizzieLet23_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet31_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet32_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet33_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet8_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet23_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet23_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet23_1_argbuf_select_q <= (lizzieLet23_1_argbuf_done ? 5'd0 :
                                        lizzieLet23_1_argbuf_select_d);
  logic [1:0] lizzieLet23_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet23_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet23_1_argbuf_emit_q <= (lizzieLet23_1_argbuf_done ? 2'd0 :
                                      lizzieLet23_1_argbuf_emit_d);
  logic [1:0] lizzieLet23_1_argbuf_emit_d;
  assign lizzieLet23_1_argbuf_emit_d = (lizzieLet23_1_argbuf_emit_q | ({writeMerge_choice_CTkron_kron_Int_Int_Int_d[0],
                                                                        writeMerge_data_CTkron_kron_Int_Int_Int_d[0]} & {writeMerge_choice_CTkron_kron_Int_Int_Int_r,
                                                                                                                         writeMerge_data_CTkron_kron_Int_Int_Int_r}));
  logic lizzieLet23_1_argbuf_done;
  assign lizzieLet23_1_argbuf_done = (& lizzieLet23_1_argbuf_emit_d);
  assign {lizzieLet8_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet23_1_argbuf_r} = (lizzieLet23_1_argbuf_done ? lizzieLet23_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTkron_kron_Int_Int_Int_d = ((lizzieLet23_1_argbuf_select_d[0] && (! lizzieLet23_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                      ((lizzieLet23_1_argbuf_select_d[1] && (! lizzieLet23_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                       ((lizzieLet23_1_argbuf_select_d[2] && (! lizzieLet23_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                        ((lizzieLet23_1_argbuf_select_d[3] && (! lizzieLet23_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                         ((lizzieLet23_1_argbuf_select_d[4] && (! lizzieLet23_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                                          {83'd0, 1'd0})))));
  assign writeMerge_choice_CTkron_kron_Int_Int_Int_d = ((lizzieLet23_1_argbuf_select_d[0] && (! lizzieLet23_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                        ((lizzieLet23_1_argbuf_select_d[1] && (! lizzieLet23_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                         ((lizzieLet23_1_argbuf_select_d[2] && (! lizzieLet23_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                          ((lizzieLet23_1_argbuf_select_d[3] && (! lizzieLet23_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                           ((lizzieLet23_1_argbuf_select_d[4] && (! lizzieLet23_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (writeMerge_choice_CTkron_kron_Int_Int_Int,C5) (demuxWriteResult_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) > [(writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                          (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [4:0] demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTkron_kron_Int_Int_Int_d[0] && demuxWriteResult_CTkron_kron_Int_Int_Int_d[0]))
      unique case (writeMerge_choice_CTkron_kron_Int_Int_Int_d[3:1])
        3'd0: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd = 5'd0;
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[0]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[1]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[2]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                               demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[3]};
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d = {demuxWriteResult_CTkron_kron_Int_Int_Int_d[16:1],
                                                              demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd[4]};
  assign demuxWriteResult_CTkron_kron_Int_Int_Int_r = (| (demuxWriteResult_CTkron_kron_Int_Int_Int_onehotd & {writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r,
                                                                                                              writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_r}));
  assign writeMerge_choice_CTkron_kron_Int_Int_Int_r = demuxWriteResult_CTkron_kron_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Int_Int_Int,
      Dcon WriteIn_CTkron_kron_Int_Int_Int) : [(forkHP1_CTkron_kron_Int_Int_In2,Word16#),
                                               (writeMerge_data_CTkron_kron_Int_Int_Int,CTkron_kron_Int_Int_Int)] > (dconWriteIn_CTkron_kron_Int_Int_Int,MemIn_CTkron_kron_Int_Int_Int) */
  assign dconWriteIn_CTkron_kron_Int_Int_Int_d = WriteIn_CTkron_kron_Int_Int_Int_dc((& {forkHP1_CTkron_kron_Int_Int_In2_d[0],
                                                                                        writeMerge_data_CTkron_kron_Int_Int_Int_d[0]}), forkHP1_CTkron_kron_Int_Int_In2_d, writeMerge_data_CTkron_kron_Int_Int_Int_d);
  assign {forkHP1_CTkron_kron_Int_Int_In2_r,
          writeMerge_data_CTkron_kron_Int_Int_Int_r} = {2 {(dconWriteIn_CTkron_kron_Int_Int_Int_r && dconWriteIn_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTkron_kron_Int_Int_Int,
      Dcon Pointer_CTkron_kron_Int_Int_Int) : [(forkHP1_CTkron_kron_Int_Int_In3,Word16#)] > (dconPtr_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) */
  assign dconPtr_CTkron_kron_Int_Int_Int_d = Pointer_CTkron_kron_Int_Int_Int_dc((& {forkHP1_CTkron_kron_Int_Int_In3_d[0]}), forkHP1_CTkron_kron_Int_Int_In3_d);
  assign {forkHP1_CTkron_kron_Int_Int_In3_r} = {1 {(dconPtr_CTkron_kron_Int_Int_Int_r && dconPtr_CTkron_kron_Int_Int_Int_d[0])}};
  
  /* demux (Ty MemOut_CTkron_kron_Int_Int_Int,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (memWriteOut_CTkron_kron_Int_Int_Int,MemOut_CTkron_kron_Int_Int_Int) (dconPtr_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int) > [(_50,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                                                                                       (demuxWriteResult_CTkron_kron_Int_Int_Int,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [1:0] dconPtr_CTkron_kron_Int_Int_Int_onehotd;
  always_comb
    if ((memWriteOut_CTkron_kron_Int_Int_Int_d[0] && dconPtr_CTkron_kron_Int_Int_Int_d[0]))
      unique case (memWriteOut_CTkron_kron_Int_Int_Int_d[1:1])
        1'd0: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd2;
        default: dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTkron_kron_Int_Int_Int_onehotd = 2'd0;
  assign _50_d = {dconPtr_CTkron_kron_Int_Int_Int_d[16:1],
                  dconPtr_CTkron_kron_Int_Int_Int_onehotd[0]};
  assign demuxWriteResult_CTkron_kron_Int_Int_Int_d = {dconPtr_CTkron_kron_Int_Int_Int_d[16:1],
                                                       dconPtr_CTkron_kron_Int_Int_Int_onehotd[1]};
  assign dconPtr_CTkron_kron_Int_Int_Int_r = (| (dconPtr_CTkron_kron_Int_Int_Int_onehotd & {demuxWriteResult_CTkron_kron_Int_Int_Int_r,
                                                                                            _50_r}));
  assign memWriteOut_CTkron_kron_Int_Int_Int_r = dconPtr_CTkron_kron_Int_Int_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  logic [31:0] profiling_MemIn_MaskQTree_read;
  logic [31:0] profiling_MemIn_MaskQTree_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_MaskQTree_write <= 0;
        profiling_MemIn_MaskQTree_read <= 0;
      end
    else
      if ((memMergeIn_MaskQTree_dbuf_we == 1'd1))
        profiling_MemIn_MaskQTree_write <= (profiling_MemIn_MaskQTree_write + 1);
      else
        if ((memOut_MaskQTree_valid == 1'd1))
          profiling_MemIn_MaskQTree_read <= (profiling_MemIn_MaskQTree_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (mskacl_1_argbuf,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {mskacl_1_argbuf_d[16:1],
                                       mskacl_1_argbuf_d[0]};
  assign mskacl_1_argbuf_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(readPointer_MaskQTreemskacl_1_argbuf,MaskQTree)] */
  assign readPointer_MaskQTreemskacl_1_argbuf_d = {memReadOut_MaskQTree_d[67:2],
                                                   memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = readPointer_MaskQTreemskacl_1_argbuf_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_49,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _49_d = {dconPtr_MaskQTree_d[16:1],
                  dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _49_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1adl_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2adm_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m3adn_2,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnz_IntTupGo___Pointer_QTree_Intgo_6,Go),
                                                                                                                ($wnnz_IntTupGo___Pointer_QTree_Intwsxl,Pointer_QTree_Int)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_d  = {\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [16:1],
                                                       (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_done  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnz_IntTupGo___Pointer_QTree_Intwsxl_d [0],
                                                                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0]} & {\$wnnz_IntTupGo___Pointer_QTree_Intwsxl_r ,
                                                                                                                                                             \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r }));
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                         \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnz_IntTupGo___Pointer_QTree_Intgo_6,Go) > [(go_6_1,Go),
                                                              (go_6_2,Go)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done ;
  assign go_6_1_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted [0]));
  assign go_6_2_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted [1]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done  = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  | ({go_6_2_d[0],
                                                                                                               go_6_1_d[0]} & {go_6_2_r,
                                                                                                                               go_6_1_r}));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r  ? 2'd0 :
                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Intwsxl,Pointer_QTree_Int) > (wsxl_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_r ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_r  = ((! \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d [0]) || \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d  <= {16'd0,
                                                             1'd0};
    else
      if (\$wnnz_IntTupGo___Pointer_QTree_Intwsxl_r )
        \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_d ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_r  = (! \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf [0]);
  assign wsxl_1_argbuf_d = (\$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf [0] ? \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf  :
                            \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf  <= {16'd0,
                                                               1'd0};
    else
      if ((wsxl_1_argbuf_r && \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf [0]))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf  <= {16'd0,
                                                                 1'd0};
      else if (((! wsxl_1_argbuf_r) && (! \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf [0])))
        \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_buf  <= \$wnnz_IntTupGo___Pointer_QTree_Intwsxl_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_Int_resbuf,Int#)] > (es_7_1I#,Int) */
  assign \es_7_1I#_d  = \I#_dc ((& {\$wnnz_Int_resbuf_d [0]}), \$wnnz_Int_resbuf_d );
  assign {\$wnnz_Int_resbuf_r } = {1 {(\es_7_1I#_r  && \es_7_1I#_d [0])}};
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go),
                                                                                                                           (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                                           (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[32:1],
                                                              (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[2]))};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                                                                         applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                                                                         applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r ? 3'd0 :
                                                                applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done);
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_0_2_1,MyBool),
                                                        (es_0_2_2,MyBool),
                                                        (es_0_2_3,MyBool)] */
  logic [2:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [2:0] applyfnInt_Bool_5_resbuf_done;
  assign es_0_2_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_0_2_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_0_2_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                       (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_0_2_3_d[0],
                                                                               es_0_2_2_d[0],
                                                                               es_0_2_1_d[0]} & {es_0_2_3_r,
                                                                                                 es_0_2_2_r,
                                                                                                 es_0_2_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 3'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[32:1],
                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[64:33],
                                                                       (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[2]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r ? 3'd0 :
                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int) > [(arg0_2_1,MyDTInt_Int_Int),
                                                                                                          (arg0_2_2,MyDTInt_Int_Int),
                                                                                                          (arg0_2_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                                               arg0_2_2_d[0],
                                                                                                                                               arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                                                 arg0_2_2_r,
                                                                                                                                                                 arg0_2_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  
  /* fork (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > [(xac0_1,Int),
                                                     (xac0_2,Int)] */
  logic [1:0] applyfnInt_Int_Int_5_resbuf_emitted;
  logic [1:0] applyfnInt_Int_Int_5_resbuf_done;
  assign xac0_1_d = {applyfnInt_Int_Int_5_resbuf_d[32:1],
                     (applyfnInt_Int_Int_5_resbuf_d[0] && (! applyfnInt_Int_Int_5_resbuf_emitted[0]))};
  assign xac0_2_d = {applyfnInt_Int_Int_5_resbuf_d[32:1],
                     (applyfnInt_Int_Int_5_resbuf_d[0] && (! applyfnInt_Int_Int_5_resbuf_emitted[1]))};
  assign applyfnInt_Int_Int_5_resbuf_done = (applyfnInt_Int_Int_5_resbuf_emitted | ({xac0_2_d[0],
                                                                                     xac0_1_d[0]} & {xac0_2_r,
                                                                                                     xac0_1_r}));
  assign applyfnInt_Int_Int_5_resbuf_r = (& applyfnInt_Int_Int_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_resbuf_emitted <= 2'd0;
    else
      applyfnInt_Int_Int_5_resbuf_emitted <= (applyfnInt_Int_Int_5_resbuf_r ? 2'd0 :
                                              applyfnInt_Int_Int_5_resbuf_done);
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_main1,Int)] */
  assign arg0_1Dcon_main1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                               (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_main1,Int) > [(arg0_1Dcon_main1_1,Int),
                                          (arg0_1Dcon_main1_2,Int),
                                          (arg0_1Dcon_main1_3,Int),
                                          (arg0_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_1Dcon_main1_emitted;
  logic [3:0] arg0_1Dcon_main1_done;
  assign arg0_1Dcon_main1_1_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[0]))};
  assign arg0_1Dcon_main1_2_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[1]))};
  assign arg0_1Dcon_main1_3_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[2]))};
  assign arg0_1Dcon_main1_4_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[3]))};
  assign arg0_1Dcon_main1_done = (arg0_1Dcon_main1_emitted | ({arg0_1Dcon_main1_4_d[0],
                                                               arg0_1Dcon_main1_3_d[0],
                                                               arg0_1Dcon_main1_2_d[0],
                                                               arg0_1Dcon_main1_1_d[0]} & {arg0_1Dcon_main1_4_r,
                                                                                           arg0_1Dcon_main1_3_r,
                                                                                           arg0_1Dcon_main1_2_r,
                                                                                           arg0_1Dcon_main1_1_r}));
  assign arg0_1Dcon_main1_r = (& arg0_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_1Dcon_main1_emitted <= (arg0_1Dcon_main1_r ? 4'd0 :
                                   arg0_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_main1_1I#,Int) > [(xase_destruct,Int#)] */
  assign xase_destruct_d = {\arg0_1Dcon_main1_1I#_d [32:1],
                            \arg0_1Dcon_main1_1I#_d [0]};
  assign \arg0_1Dcon_main1_1I#_r  = xase_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_main1_2,Int) (arg0_1Dcon_main1_1,Int) > [(arg0_1Dcon_main1_1I#,Int)] */
  assign \arg0_1Dcon_main1_1I#_d  = {arg0_1Dcon_main1_1_d[32:1],
                                     (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0])};
  assign arg0_1Dcon_main1_1_r = (\arg0_1Dcon_main1_1I#_r  && (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0]));
  assign arg0_1Dcon_main1_2_r = (\arg0_1Dcon_main1_1I#_r  && (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_main1_3,Int) (arg0_2Dcon_main1,Go) > [(arg0_1Dcon_main1_3I#,Go)] */
  assign \arg0_1Dcon_main1_3I#_d  = (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]);
  assign arg0_2Dcon_main1_r = (\arg0_1Dcon_main1_3I#_r  && (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]));
  assign arg0_1Dcon_main1_3_r = (\arg0_1Dcon_main1_3I#_r  && (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_main1_3I#,Go) > [(arg0_1Dcon_main1_3I#_1,Go),
                                            (arg0_1Dcon_main1_3I#_2,Go),
                                            (arg0_1Dcon_main1_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_main1_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_main1_3I#_done ;
  assign \arg0_1Dcon_main1_3I#_1_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [0]));
  assign \arg0_1Dcon_main1_3I#_2_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [1]));
  assign \arg0_1Dcon_main1_3I#_3_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [2]));
  assign \arg0_1Dcon_main1_3I#_done  = (\arg0_1Dcon_main1_3I#_emitted  | ({\arg0_1Dcon_main1_3I#_3_d [0],
                                                                           \arg0_1Dcon_main1_3I#_2_d [0],
                                                                           \arg0_1Dcon_main1_3I#_1_d [0]} & {\arg0_1Dcon_main1_3I#_3_r ,
                                                                                                             \arg0_1Dcon_main1_3I#_2_r ,
                                                                                                             \arg0_1Dcon_main1_3I#_1_r }));
  assign \arg0_1Dcon_main1_3I#_r  = (& \arg0_1Dcon_main1_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_main1_3I#_emitted  <= (\arg0_1Dcon_main1_3I#_r  ? 3'd0 :
                                         \arg0_1Dcon_main1_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_main1_3I#_1,Go) > (arg0_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_main1_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_main1_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_main1_3I#_1_r  = ((! \arg0_1Dcon_main1_3I#_1_bufchan_d [0]) || \arg0_1Dcon_main1_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_main1_3I#_1_r )
        \arg0_1Dcon_main1_3I#_1_bufchan_d  <= \arg0_1Dcon_main1_3I#_1_d ;
  Go_t \arg0_1Dcon_main1_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_main1_3I#_1_bufchan_r  = (! \arg0_1Dcon_main1_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_1Dcon_main1_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_main1_3I#_1_bufchan_buf  :
                                              \arg0_1Dcon_main1_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_main1_3I#_1_argbuf_r  && \arg0_1Dcon_main1_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_1Dcon_main1_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= \arg0_1Dcon_main1_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_1Dcon_main1_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_main1_3I#_1_argbuf_0_d  = {32'd0,
                                                \arg0_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_main1_3I#_1_argbuf_r  = \arg0_1Dcon_main1_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_main1_3I#_1_argbuf_0,Int#) (xase_destruct,Int#) > (lizzieLet1_1wild1X1j_1_Eq,Bool) */
  assign lizzieLet1_1wild1X1j_1_Eq_d = {(\arg0_1Dcon_main1_3I#_1_argbuf_0_d [32:1] == xase_destruct_d[32:1]),
                                        (\arg0_1Dcon_main1_3I#_1_argbuf_0_d [0] && xase_destruct_d[0])};
  assign {\arg0_1Dcon_main1_3I#_1_argbuf_0_r ,
          xase_destruct_r} = {2 {(lizzieLet1_1wild1X1j_1_Eq_r && lizzieLet1_1wild1X1j_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_main1_3I#_2,Go) > (arg0_1Dcon_main1_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_main1_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_main1_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_main1_3I#_2_r  = ((! \arg0_1Dcon_main1_3I#_2_bufchan_d [0]) || \arg0_1Dcon_main1_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_main1_3I#_2_r )
        \arg0_1Dcon_main1_3I#_2_bufchan_d  <= \arg0_1Dcon_main1_3I#_2_d ;
  Go_t \arg0_1Dcon_main1_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_main1_3I#_2_bufchan_r  = (! \arg0_1Dcon_main1_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_main1_3I#_2_argbuf_d  = (\arg0_1Dcon_main1_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_main1_3I#_2_bufchan_buf  :
                                              \arg0_1Dcon_main1_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_main1_3I#_2_argbuf_r  && \arg0_1Dcon_main1_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_main1_3I#_2_argbuf_r ) && (! \arg0_1Dcon_main1_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= \arg0_1Dcon_main1_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_main1_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_main1_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_main1_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_main1_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_main1_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_main1_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go) > [(arg0_2Dcon_main1,Go)] */
  assign arg0_2Dcon_main1_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  assign arg0_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int) > [(arg0_2_1Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_2_1Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[32:1],
                                              (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r = (\arg0_2_1Dcon_$fNumInt_$ctimes_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (\arg0_2_1Dcon_$fNumInt_$ctimes_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_2_2Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                              (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_2_2Dcon_$fNumInt_$ctimes_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_2_2_r = (\arg0_2_2Dcon_$fNumInt_$ctimes_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*,Int) > [(arg0_2_2Dcon_$fNumInt_$c*_1,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c*_2,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c*_3,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c*_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$ctimes_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$ctimes_done ;
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_1_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_2_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_4_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_done  = (\arg0_2_2Dcon_$fNumInt_$ctimes_emitted  | ({\arg0_2_2Dcon_$fNumInt_$ctimes_4_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$ctimes_3_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$ctimes_2_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$ctimes_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$ctimes_4_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$ctimes_3_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$ctimes_2_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$ctimes_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_r  = (& \arg0_2_2Dcon_$fNumInt_$ctimes_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_$fNumInt_$ctimes_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$ctimes_emitted  <= (\arg0_2_2Dcon_$fNumInt_$ctimes_r  ? 4'd0 :
                                                  \arg0_2_2Dcon_$fNumInt_$ctimes_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c*_1I#,Int) > [(xa1m0_destruct,Int#)] */
  assign xa1m0_destruct_d = {\arg0_2_2Dcon_$fNumInt_$ctimes_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$ctimes_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_1I#_r  = xa1m0_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_2,Int) (arg0_2_2Dcon_$fNumInt_$c*_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c*_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_1_d [32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_1_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_2_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_3,Int) (arg0_2_1Dcon_$fNumInt_$c*,Int) > [(arg0_2_2Dcon_$fNumInt_$c*_3I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d  = {\arg0_2_1Dcon_$fNumInt_$ctimes_d [32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_2_1Dcon_$fNumInt_$ctimes_d [0])};
  assign \arg0_2_1Dcon_$fNumInt_$ctimes_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_2_1Dcon_$fNumInt_$ctimes_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_2_1Dcon_$fNumInt_$ctimes_d [0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_3I#,Int) > [(arg0_2_2Dcon_$fNumInt_$c*_3I#_1,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c*_3I#_2,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c*_3I#_3,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c*_3I#_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_done ;
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_done  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted  | ({\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d [0],
                                                                                                     \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d [0],
                                                                                                     \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d [0],
                                                                                                     \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_r ,
                                                                                                                                                    \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_r ,
                                                                                                                                                    \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_r ,
                                                                                                                                                    \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_r  = (& \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_r  ? 4'd0 :
                                                      \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c*_3I#_1I#,Int) > [(ya1m1_destruct,Int#)] */
  assign ya1m1_destruct_d = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  = ya1m1_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_3I#_2,Int) (arg0_2_2Dcon_$fNumInt_$c*_3I#_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c*_3I#_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d [32:1],
                                                      (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c*_3I#_3,Int) (xa1m0_destruct,Int#) > [(arg0_2_2Dcon_$fNumInt_$c*_3I#_3I#,Int#)] */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_d  = {xa1m0_destruct_d[32:1],
                                                      (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0])};
  assign xa1m0_destruct_r = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_r  = (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  
  /* op_mul (Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c*_3I#_3I#,Int#) (ya1m1_destruct,Int#) > (arg0_2_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#) */
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d  = {(\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [32:1] * ya1m1_destruct_d[32:1]),
                                                                     (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [0] && ya1m1_destruct_d[0])};
  assign {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ,
          ya1m1_destruct_r} = {2 {(\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r  && \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_2_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0]}), \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d );
  assign {\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r } = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_3I#_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c*_4,Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (\arg0_2_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_1_1I#_mux_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$ctimes_4_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int_Int) [(es_0_1_1I#_mux_mux,Int)] > (es_0_1_1I#_mux_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_mux_d  = {\es_0_1_1I#_mux_mux_d [32:1],
                                       (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0])};
  assign \es_0_1_1I#_mux_mux_r  = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  assign arg0_2_3_r = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) > [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8,Go),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1,Pointer_QTree_Int),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] */
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted;
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done;
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[0]));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[16:1],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[1]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[32:17],
                                                                                (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[2]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted | ({call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]} & {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r}));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r = (& call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= 3'd0;
    else
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r ? 3'd0 :
                                                                                  call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_Int_goConst,Go) > (call_$wnnz_Int_initBufi,Go) */
  Go_t call_$wnnz_Int_goConst_buf;
  assign call_$wnnz_Int_goConst_r = (! call_$wnnz_Int_goConst_buf[0]);
  assign call_$wnnz_Int_initBufi_d = (call_$wnnz_Int_goConst_buf[0] ? call_$wnnz_Int_goConst_buf :
                                      call_$wnnz_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_Int_initBufi_r && call_$wnnz_Int_goConst_buf[0]))
        call_$wnnz_Int_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_Int_initBufi_r) && (! call_$wnnz_Int_goConst_buf[0])))
        call_$wnnz_Int_goConst_buf <= call_$wnnz_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_Int_goMux1,Go),
                           (lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf,Go),
                           (lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf,Go),
                           (lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_8_goMux_choice,C5) (go_8_goMux_data,Go) */
  logic [4:0] call_$wnnz_Int_goMux1_select_d;
  assign call_$wnnz_Int_goMux1_select_d = ((| call_$wnnz_Int_goMux1_select_q) ? call_$wnnz_Int_goMux1_select_q :
                                           (call_$wnnz_Int_goMux1_d[0] ? 5'd1 :
                                            (lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_d[0] ? 5'd2 :
                                             (lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_d[0] ? 5'd4 :
                                              (lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_d[0] ? 5'd8 :
                                               (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                5'd0))))));
  logic [4:0] call_$wnnz_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_Int_goMux1_select_q <= (call_$wnnz_Int_goMux1_done ? 5'd0 :
                                         call_$wnnz_Int_goMux1_select_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_Int_goMux1_emit_q <= (call_$wnnz_Int_goMux1_done ? 2'd0 :
                                       call_$wnnz_Int_goMux1_emit_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_d;
  assign call_$wnnz_Int_goMux1_emit_d = (call_$wnnz_Int_goMux1_emit_q | ({go_8_goMux_choice_d[0],
                                                                          go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                   go_8_goMux_data_r}));
  logic call_$wnnz_Int_goMux1_done;
  assign call_$wnnz_Int_goMux1_done = (& call_$wnnz_Int_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_r,
          lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_r,
          lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_r,
          call_$wnnz_Int_goMux1_r} = (call_$wnnz_Int_goMux1_done ? call_$wnnz_Int_goMux1_select_d :
                                      5'd0);
  assign go_8_goMux_data_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? call_$wnnz_Int_goMux1_d :
                              ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_d :
                               ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_d :
                                ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_d :
                                 ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_8_goMux_choice_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_Int_initBuf,Go) > [(call_$wnnz_Int_unlockFork1,Go),
                                              (call_$wnnz_Int_unlockFork2,Go),
                                              (call_$wnnz_Int_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_Int_initBuf_emitted;
  logic [2:0] call_$wnnz_Int_initBuf_done;
  assign call_$wnnz_Int_unlockFork1_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[0]));
  assign call_$wnnz_Int_unlockFork2_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[1]));
  assign call_$wnnz_Int_unlockFork3_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[2]));
  assign call_$wnnz_Int_initBuf_done = (call_$wnnz_Int_initBuf_emitted | ({call_$wnnz_Int_unlockFork3_d[0],
                                                                           call_$wnnz_Int_unlockFork2_d[0],
                                                                           call_$wnnz_Int_unlockFork1_d[0]} & {call_$wnnz_Int_unlockFork3_r,
                                                                                                               call_$wnnz_Int_unlockFork2_r,
                                                                                                               call_$wnnz_Int_unlockFork1_r}));
  assign call_$wnnz_Int_initBuf_r = (& call_$wnnz_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_Int_initBuf_emitted <= (call_$wnnz_Int_initBuf_r ? 3'd0 :
                                         call_$wnnz_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_Int_initBufi,Go) > (call_$wnnz_Int_initBuf,Go) */
  assign call_$wnnz_Int_initBufi_r = ((! call_$wnnz_Int_initBuf_d[0]) || call_$wnnz_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_Int_initBufi_r)
        call_$wnnz_Int_initBuf_d <= call_$wnnz_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_Int_unlockFork1,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8,Go)] > (call_$wnnz_Int_goMux1,Go) */
  assign call_$wnnz_Int_goMux1_d = (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]);
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]));
  assign call_$wnnz_Int_unlockFork1_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_Int_unlockFork2,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1,Pointer_QTree_Int)] > (call_$wnnz_Int_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_Int_goMux2_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d[0]));
  assign call_$wnnz_Int_unlockFork2_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intwsxl_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz_Int) : (call_$wnnz_Int_unlockFork3,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] > (call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int) */
  assign call_$wnnz_Int_goMux3_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[16:1],
                                    (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  assign call_$wnnz_Int_unlockFork3_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) : (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) > [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9,Go),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                      (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [5:0] call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted;
  logic [5:0] call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done;
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[0]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[1]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[2]));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[16:1],
                                                                                                                                                              (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[3]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[32:17],
                                                                                                                                                              (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[4]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[48:33],
                                                                                                                                                               (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0] && (! call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted[5]))};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done = (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted | ({call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d[0],
                                                                                                                                                                                                                                                                                                                       call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d[0]} & {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_r}));
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r = (& call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted <= 6'd0;
    else
      call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_emitted <= (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r ? 6'd0 :
                                                                                                                                                               call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_done);
  
  /* rbuf (Ty Go) : (call_kron_kron_Int_Int_Int_goConst,Go) > (call_kron_kron_Int_Int_Int_initBufi,Go) */
  Go_t call_kron_kron_Int_Int_Int_goConst_buf;
  assign call_kron_kron_Int_Int_Int_goConst_r = (! call_kron_kron_Int_Int_Int_goConst_buf[0]);
  assign call_kron_kron_Int_Int_Int_initBufi_d = (call_kron_kron_Int_Int_Int_goConst_buf[0] ? call_kron_kron_Int_Int_Int_goConst_buf :
                                                  call_kron_kron_Int_Int_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goConst_buf <= 1'd0;
    else
      if ((call_kron_kron_Int_Int_Int_initBufi_r && call_kron_kron_Int_Int_Int_goConst_buf[0]))
        call_kron_kron_Int_Int_Int_goConst_buf <= 1'd0;
      else if (((! call_kron_kron_Int_Int_Int_initBufi_r) && (! call_kron_kron_Int_Int_Int_goConst_buf[0])))
        call_kron_kron_Int_Int_Int_goConst_buf <= call_kron_kron_Int_Int_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_kron_kron_Int_Int_Int_goMux1,Go),
                           (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf,Go),
                           (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf,Go),
                           (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf,Go),
                           (lizzieLet6_4QNode_Int_1_argbuf,Go)] > (go_9_goMux_choice,C5) (go_9_goMux_data,Go) */
  logic [4:0] call_kron_kron_Int_Int_Int_goMux1_select_d;
  assign call_kron_kron_Int_Int_Int_goMux1_select_d = ((| call_kron_kron_Int_Int_Int_goMux1_select_q) ? call_kron_kron_Int_Int_Int_goMux1_select_q :
                                                       (call_kron_kron_Int_Int_Int_goMux1_d[0] ? 5'd1 :
                                                        (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d[0] ? 5'd2 :
                                                         (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d[0] ? 5'd4 :
                                                          (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d[0] ? 5'd8 :
                                                           (lizzieLet6_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                            5'd0))))));
  logic [4:0] call_kron_kron_Int_Int_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goMux1_select_q <= 5'd0;
    else
      call_kron_kron_Int_Int_Int_goMux1_select_q <= (call_kron_kron_Int_Int_Int_goMux1_done ? 5'd0 :
                                                     call_kron_kron_Int_Int_Int_goMux1_select_d);
  logic [1:0] call_kron_kron_Int_Int_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_goMux1_emit_q <= 2'd0;
    else
      call_kron_kron_Int_Int_Int_goMux1_emit_q <= (call_kron_kron_Int_Int_Int_goMux1_done ? 2'd0 :
                                                   call_kron_kron_Int_Int_Int_goMux1_emit_d);
  logic [1:0] call_kron_kron_Int_Int_Int_goMux1_emit_d;
  assign call_kron_kron_Int_Int_Int_goMux1_emit_d = (call_kron_kron_Int_Int_Int_goMux1_emit_q | ({go_9_goMux_choice_d[0],
                                                                                                  go_9_goMux_data_d[0]} & {go_9_goMux_choice_r,
                                                                                                                           go_9_goMux_data_r}));
  logic call_kron_kron_Int_Int_Int_goMux1_done;
  assign call_kron_kron_Int_Int_Int_goMux1_done = (& call_kron_kron_Int_Int_Int_goMux1_emit_d);
  assign {lizzieLet6_4QNode_Int_1_argbuf_r,
          lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r,
          lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r,
          lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux1_r} = (call_kron_kron_Int_Int_Int_goMux1_done ? call_kron_kron_Int_Int_Int_goMux1_select_d :
                                                  5'd0);
  assign go_9_goMux_data_d = ((call_kron_kron_Int_Int_Int_goMux1_select_d[0] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? call_kron_kron_Int_Int_Int_goMux1_d :
                              ((call_kron_kron_Int_Int_Int_goMux1_select_d[1] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d :
                               ((call_kron_kron_Int_Int_Int_goMux1_select_d[2] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d :
                                ((call_kron_kron_Int_Int_Int_goMux1_select_d[3] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d :
                                 ((call_kron_kron_Int_Int_Int_goMux1_select_d[4] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet6_4QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_9_goMux_choice_d = ((call_kron_kron_Int_Int_Int_goMux1_select_d[0] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_kron_kron_Int_Int_Int_goMux1_select_d[1] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_kron_kron_Int_Int_Int_goMux1_select_d[2] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_kron_kron_Int_Int_Int_goMux1_select_d[3] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_kron_kron_Int_Int_Int_goMux1_select_d[4] && (! call_kron_kron_Int_Int_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_kron_kron_Int_Int_Int_initBuf,Go) > [(call_kron_kron_Int_Int_Int_unlockFork1,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork2,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork3,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork4,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork5,Go),
                                                          (call_kron_kron_Int_Int_Int_unlockFork6,Go)] */
  logic [5:0] call_kron_kron_Int_Int_Int_initBuf_emitted;
  logic [5:0] call_kron_kron_Int_Int_Int_initBuf_done;
  assign call_kron_kron_Int_Int_Int_unlockFork1_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork2_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[1]));
  assign call_kron_kron_Int_Int_Int_unlockFork3_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[2]));
  assign call_kron_kron_Int_Int_Int_unlockFork4_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[3]));
  assign call_kron_kron_Int_Int_Int_unlockFork5_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[4]));
  assign call_kron_kron_Int_Int_Int_unlockFork6_d = (call_kron_kron_Int_Int_Int_initBuf_d[0] && (! call_kron_kron_Int_Int_Int_initBuf_emitted[5]));
  assign call_kron_kron_Int_Int_Int_initBuf_done = (call_kron_kron_Int_Int_Int_initBuf_emitted | ({call_kron_kron_Int_Int_Int_unlockFork6_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork5_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork4_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork3_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork2_d[0],
                                                                                                   call_kron_kron_Int_Int_Int_unlockFork1_d[0]} & {call_kron_kron_Int_Int_Int_unlockFork6_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork5_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork4_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork3_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork2_r,
                                                                                                                                                   call_kron_kron_Int_Int_Int_unlockFork1_r}));
  assign call_kron_kron_Int_Int_Int_initBuf_r = (& call_kron_kron_Int_Int_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_initBuf_emitted <= 6'd0;
    else
      call_kron_kron_Int_Int_Int_initBuf_emitted <= (call_kron_kron_Int_Int_Int_initBuf_r ? 6'd0 :
                                                     call_kron_kron_Int_Int_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_kron_kron_Int_Int_Int_initBufi,Go) > (call_kron_kron_Int_Int_Int_initBuf,Go) */
  assign call_kron_kron_Int_Int_Int_initBufi_r = ((! call_kron_kron_Int_Int_Int_initBuf_d[0]) || call_kron_kron_Int_Int_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Int_Int_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_kron_kron_Int_Int_Int_initBufi_r)
        call_kron_kron_Int_Int_Int_initBuf_d <= call_kron_kron_Int_Int_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_kron_kron_Int_Int_Int_unlockFork1,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9,Go)] > (call_kron_kron_Int_Int_Int_goMux1,Go) */
  assign call_kron_kron_Int_Int_Int_goMux1_d = (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_r = (call_kron_kron_Int_Int_Int_goMux1_r && (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork1_r = (call_kron_kron_Int_Int_Int_goMux1_r && (call_kron_kron_Int_Int_Int_unlockFork1_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intgo_9_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_kron_kron_Int_Int_Int_unlockFork2,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL,MyDTInt_Bool)] > (call_kron_kron_Int_Int_Int_goMux2,MyDTInt_Bool) */
  assign call_kron_kron_Int_Int_Int_goMux2_d = (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_r = (call_kron_kron_Int_Int_Int_goMux2_r && (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork2_r = (call_kron_kron_Int_Int_Int_goMux2_r && (call_kron_kron_Int_Int_Int_unlockFork2_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntisZacL_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_kron_kron_Int_Int_Int_unlockFork3,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM,MyDTInt_Int_Int)] > (call_kron_kron_Int_Int_Int_goMux3,MyDTInt_Int_Int) */
  assign call_kron_kron_Int_Int_Int_goMux3_d = (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d[0]);
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_r = (call_kron_kron_Int_Int_Int_goMux3_r && (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork3_r = (call_kron_kron_Int_Int_Int_goMux3_r && (call_kron_kron_Int_Int_Int_unlockFork3_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_IntgacM_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_kron_kron_Int_Int_Int_unlockFork4,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN,Pointer_QTree_Int)] > (call_kron_kron_Int_Int_Int_goMux4,Pointer_QTree_Int) */
  assign call_kron_kron_Int_Int_Int_goMux4_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_r = (call_kron_kron_Int_Int_Int_goMux4_r && (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork4_r = (call_kron_kron_Int_Int_Int_goMux4_r && (call_kron_kron_Int_Int_Int_unlockFork4_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm1acN_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_kron_kron_Int_Int_Int_unlockFork5,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO,Pointer_QTree_Int)] > (call_kron_kron_Int_Int_Int_goMux5,Pointer_QTree_Int) */
  assign call_kron_kron_Int_Int_Int_goMux5_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_r = (call_kron_kron_Int_Int_Int_goMux5_r && (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork5_r = (call_kron_kron_Int_Int_Int_goMux5_r && (call_kron_kron_Int_Int_Int_unlockFork5_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intm2acO_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (call_kron_kron_Int_Int_Int_unlockFork6,Go) [(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1,Pointer_CTkron_kron_Int_Int_Int)] > (call_kron_kron_Int_Int_Int_goMux6,Pointer_CTkron_kron_Int_Int_Int) */
  assign call_kron_kron_Int_Int_Int_goMux6_d = {call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[16:1],
                                                (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0])};
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_r = (call_kron_kron_Int_Int_Int_goMux6_r && (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0]));
  assign call_kron_kron_Int_Int_Int_unlockFork6_r = (call_kron_kron_Int_Int_Int_goMux6_r && (call_kron_kron_Int_Int_Int_unlockFork6_d[0] && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Intsc_0_1_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) : (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) > [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10,Go),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                   (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2,Pointer_CTmain_mask_Int)] */
  logic [3:0] call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted;
  logic [3:0] call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done;
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d = (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[0]));
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[16:1],
                                                                                                            (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[1]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[32:17],
                                                                                                              (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[2]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[48:33],
                                                                                                              (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0] && (! call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted[3]))};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done = (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted | ({call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d[0],
                                                                                                                                                                                                                     call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d[0]} & {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r,
                                                                                                                                                                                                                                                                                                                             call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_r,
                                                                                                                                                                                                                                                                                                                             call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_r,
                                                                                                                                                                                                                                                                                                                             call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_r}));
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r = (& call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted <= 4'd0;
    else
      call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_emitted <= (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r ? 4'd0 :
                                                                                                              call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_done);
  
  /* rbuf (Ty Go) : (call_main_mask_Int_goConst,Go) > (call_main_mask_Int_initBufi,Go) */
  Go_t call_main_mask_Int_goConst_buf;
  assign call_main_mask_Int_goConst_r = (! call_main_mask_Int_goConst_buf[0]);
  assign call_main_mask_Int_initBufi_d = (call_main_mask_Int_goConst_buf[0] ? call_main_mask_Int_goConst_buf :
                                          call_main_mask_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goConst_buf <= 1'd0;
    else
      if ((call_main_mask_Int_initBufi_r && call_main_mask_Int_goConst_buf[0]))
        call_main_mask_Int_goConst_buf <= 1'd0;
      else if (((! call_main_mask_Int_initBufi_r) && (! call_main_mask_Int_goConst_buf[0])))
        call_main_mask_Int_goConst_buf <= call_main_mask_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_mask_Int_goMux1,Go),
                           (lizzieLet35_3Lcall_main_mask_Int3_1_argbuf,Go),
                           (lizzieLet35_3Lcall_main_mask_Int2_1_argbuf,Go),
                           (lizzieLet35_3Lcall_main_mask_Int1_1_argbuf,Go),
                           (lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf,Go)] > (go_10_goMux_choice,C5) (go_10_goMux_data,Go) */
  logic [4:0] call_main_mask_Int_goMux1_select_d;
  assign call_main_mask_Int_goMux1_select_d = ((| call_main_mask_Int_goMux1_select_q) ? call_main_mask_Int_goMux1_select_q :
                                               (call_main_mask_Int_goMux1_d[0] ? 5'd1 :
                                                (lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_d[0] ? 5'd2 :
                                                 (lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_d[0] ? 5'd4 :
                                                  (lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_d[0] ? 5'd8 :
                                                   (lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                    5'd0))))));
  logic [4:0] call_main_mask_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goMux1_select_q <= 5'd0;
    else
      call_main_mask_Int_goMux1_select_q <= (call_main_mask_Int_goMux1_done ? 5'd0 :
                                             call_main_mask_Int_goMux1_select_d);
  logic [1:0] call_main_mask_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_goMux1_emit_q <= 2'd0;
    else
      call_main_mask_Int_goMux1_emit_q <= (call_main_mask_Int_goMux1_done ? 2'd0 :
                                           call_main_mask_Int_goMux1_emit_d);
  logic [1:0] call_main_mask_Int_goMux1_emit_d;
  assign call_main_mask_Int_goMux1_emit_d = (call_main_mask_Int_goMux1_emit_q | ({go_10_goMux_choice_d[0],
                                                                                  go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                            go_10_goMux_data_r}));
  logic call_main_mask_Int_goMux1_done;
  assign call_main_mask_Int_goMux1_done = (& call_main_mask_Int_goMux1_emit_d);
  assign {lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_r,
          lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_r,
          lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_r,
          lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_r,
          call_main_mask_Int_goMux1_r} = (call_main_mask_Int_goMux1_done ? call_main_mask_Int_goMux1_select_d :
                                          5'd0);
  assign go_10_goMux_data_d = ((call_main_mask_Int_goMux1_select_d[0] && (! call_main_mask_Int_goMux1_emit_q[0])) ? call_main_mask_Int_goMux1_d :
                               ((call_main_mask_Int_goMux1_select_d[1] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_d :
                                ((call_main_mask_Int_goMux1_select_d[2] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_d :
                                 ((call_main_mask_Int_goMux1_select_d[3] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_d :
                                  ((call_main_mask_Int_goMux1_select_d[4] && (! call_main_mask_Int_goMux1_emit_q[0])) ? lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_10_goMux_choice_d = ((call_main_mask_Int_goMux1_select_d[0] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_main_mask_Int_goMux1_select_d[1] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_main_mask_Int_goMux1_select_d[2] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_main_mask_Int_goMux1_select_d[3] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_main_mask_Int_goMux1_select_d[4] && (! call_main_mask_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_mask_Int_initBuf,Go) > [(call_main_mask_Int_unlockFork1,Go),
                                                  (call_main_mask_Int_unlockFork2,Go),
                                                  (call_main_mask_Int_unlockFork3,Go),
                                                  (call_main_mask_Int_unlockFork4,Go)] */
  logic [3:0] call_main_mask_Int_initBuf_emitted;
  logic [3:0] call_main_mask_Int_initBuf_done;
  assign call_main_mask_Int_unlockFork1_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[0]));
  assign call_main_mask_Int_unlockFork2_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[1]));
  assign call_main_mask_Int_unlockFork3_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[2]));
  assign call_main_mask_Int_unlockFork4_d = (call_main_mask_Int_initBuf_d[0] && (! call_main_mask_Int_initBuf_emitted[3]));
  assign call_main_mask_Int_initBuf_done = (call_main_mask_Int_initBuf_emitted | ({call_main_mask_Int_unlockFork4_d[0],
                                                                                   call_main_mask_Int_unlockFork3_d[0],
                                                                                   call_main_mask_Int_unlockFork2_d[0],
                                                                                   call_main_mask_Int_unlockFork1_d[0]} & {call_main_mask_Int_unlockFork4_r,
                                                                                                                           call_main_mask_Int_unlockFork3_r,
                                                                                                                           call_main_mask_Int_unlockFork2_r,
                                                                                                                           call_main_mask_Int_unlockFork1_r}));
  assign call_main_mask_Int_initBuf_r = (& call_main_mask_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_initBuf_emitted <= 4'd0;
    else
      call_main_mask_Int_initBuf_emitted <= (call_main_mask_Int_initBuf_r ? 4'd0 :
                                             call_main_mask_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_mask_Int_initBufi,Go) > (call_main_mask_Int_initBuf,Go) */
  assign call_main_mask_Int_initBufi_r = ((! call_main_mask_Int_initBuf_d[0]) || call_main_mask_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_main_mask_Int_initBufi_r)
        call_main_mask_Int_initBuf_d <= call_main_mask_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_mask_Int_unlockFork1,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10,Go)] > (call_main_mask_Int_goMux1,Go) */
  assign call_main_mask_Int_goMux1_d = (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d[0]);
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_r = (call_main_mask_Int_goMux1_r && (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d[0]));
  assign call_main_mask_Int_unlockFork1_r = (call_main_mask_Int_goMux1_r && (call_main_mask_Int_unlockFork1_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intgo_10_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_main_mask_Int_unlockFork2,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack,Pointer_QTree_Int)] > (call_main_mask_Int_goMux2,Pointer_QTree_Int) */
  assign call_main_mask_Int_goMux2_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d[16:1],
                                        (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_r = (call_main_mask_Int_goMux2_r && (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d[0]));
  assign call_main_mask_Int_unlockFork2_r = (call_main_mask_Int_goMux2_r && (call_main_mask_Int_unlockFork2_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmack_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_main_mask_Int_unlockFork3,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl,Pointer_MaskQTree)] > (call_main_mask_Int_goMux3,Pointer_MaskQTree) */
  assign call_main_mask_Int_goMux3_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d[16:1],
                                        (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_r = (call_main_mask_Int_goMux3_r && (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d[0]));
  assign call_main_mask_Int_unlockFork3_r = (call_main_mask_Int_goMux3_r && (call_main_mask_Int_unlockFork3_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intmskacl_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_mask_Int) : (call_main_mask_Int_unlockFork4,Go) [(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2,Pointer_CTmain_mask_Int)] > (call_main_mask_Int_goMux4,Pointer_CTmain_mask_Int) */
  assign call_main_mask_Int_goMux4_d = {call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[16:1],
                                        (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0])};
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_r = (call_main_mask_Int_goMux4_r && (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0]));
  assign call_main_mask_Int_unlockFork4_r = (call_main_mask_Int_goMux4_r && (call_main_mask_Int_unlockFork4_d[0] && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Intsc_0_2_d[0]));
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) : (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) > [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11,Go),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE,Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                    (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [5:0] \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted ;
  logic [5:0] \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done ;
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [0]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [1]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [2]));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [32:1],
                                                                                                                                                      (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [3]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [48:33],
                                                                                                                                                     (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [4]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [64:49],
                                                                                                                                                       (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0] && (! \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted [5]))};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done  = (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  | ({\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d [0],
                                                                                                                                                                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d [0]} & {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_r }));
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  = (& \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  <= 6'd0;
    else
      \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_emitted  <= (\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  ? 6'd0 :
                                                                                                                                                       \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_done );
  
  /* rbuf (Ty Go) : (call_map''_map''_Int_Int_Int_goConst,Go) > (call_map''_map''_Int_Int_Int_initBufi,Go) */
  Go_t \call_map''_map''_Int_Int_Int_goConst_buf ;
  assign \call_map''_map''_Int_Int_Int_goConst_r  = (! \call_map''_map''_Int_Int_Int_goConst_buf [0]);
  assign \call_map''_map''_Int_Int_Int_initBufi_d  = (\call_map''_map''_Int_Int_Int_goConst_buf [0] ? \call_map''_map''_Int_Int_Int_goConst_buf  :
                                                      \call_map''_map''_Int_Int_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_map''_map''_Int_Int_Int_initBufi_r  && \call_map''_map''_Int_Int_Int_goConst_buf [0]))
        \call_map''_map''_Int_Int_Int_goConst_buf  <= 1'd0;
      else if (((! \call_map''_map''_Int_Int_Int_initBufi_r ) && (! \call_map''_map''_Int_Int_Int_goConst_buf [0])))
        \call_map''_map''_Int_Int_Int_goConst_buf  <= \call_map''_map''_Int_Int_Int_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_map''_map''_Int_Int_Int_goMux1,Go),
                     (lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf,Go),
                     (lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf,Go),
                     (lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf,Go),
                     (lizzieLet17_4QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] \call_map''_map''_Int_Int_Int_goMux1_select_d ;
  assign \call_map''_map''_Int_Int_Int_goMux1_select_d  = ((| \call_map''_map''_Int_Int_Int_goMux1_select_q ) ? \call_map''_map''_Int_Int_Int_goMux1_select_q  :
                                                           (\call_map''_map''_Int_Int_Int_goMux1_d [0] ? 5'd1 :
                                                            (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d [0] ? 5'd2 :
                                                             (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d [0] ? 5'd4 :
                                                              (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d [0] ? 5'd8 :
                                                               (lizzieLet17_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                                5'd0))))));
  logic [4:0] \call_map''_map''_Int_Int_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goMux1_select_q  <= 5'd0;
    else
      \call_map''_map''_Int_Int_Int_goMux1_select_q  <= (\call_map''_map''_Int_Int_Int_goMux1_done  ? 5'd0 :
                                                         \call_map''_map''_Int_Int_Int_goMux1_select_d );
  logic [1:0] \call_map''_map''_Int_Int_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_map''_map''_Int_Int_Int_goMux1_emit_q  <= (\call_map''_map''_Int_Int_Int_goMux1_done  ? 2'd0 :
                                                       \call_map''_map''_Int_Int_Int_goMux1_emit_d );
  logic [1:0] \call_map''_map''_Int_Int_Int_goMux1_emit_d ;
  assign \call_map''_map''_Int_Int_Int_goMux1_emit_d  = (\call_map''_map''_Int_Int_Int_goMux1_emit_q  | ({go_11_goMux_choice_d[0],
                                                                                                          go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                                    go_11_goMux_data_r}));
  logic \call_map''_map''_Int_Int_Int_goMux1_done ;
  assign \call_map''_map''_Int_Int_Int_goMux1_done  = (& \call_map''_map''_Int_Int_Int_goMux1_emit_d );
  assign {lizzieLet17_4QNode_Int_1_argbuf_r,
          \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ,
          \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ,
          \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ,
          \call_map''_map''_Int_Int_Int_goMux1_r } = (\call_map''_map''_Int_Int_Int_goMux1_done  ? \call_map''_map''_Int_Int_Int_goMux1_select_d  :
                                                      5'd0);
  assign go_11_goMux_data_d = ((\call_map''_map''_Int_Int_Int_goMux1_select_d [0] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \call_map''_map''_Int_Int_Int_goMux1_d  :
                               ((\call_map''_map''_Int_Int_Int_goMux1_select_d [1] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d  :
                                ((\call_map''_map''_Int_Int_Int_goMux1_select_d [2] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d  :
                                 ((\call_map''_map''_Int_Int_Int_goMux1_select_d [3] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d  :
                                  ((\call_map''_map''_Int_Int_Int_goMux1_select_d [4] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [0])) ? lizzieLet17_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((\call_map''_map''_Int_Int_Int_goMux1_select_d [0] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_map''_map''_Int_Int_Int_goMux1_select_d [1] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_map''_map''_Int_Int_Int_goMux1_select_d [2] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_map''_map''_Int_Int_Int_goMux1_select_d [3] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_map''_map''_Int_Int_Int_goMux1_select_d [4] && (! \call_map''_map''_Int_Int_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_map''_map''_Int_Int_Int_initBuf,Go) > [(call_map''_map''_Int_Int_Int_unlockFork1,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork2,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork3,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork4,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork5,Go),
                                                            (call_map''_map''_Int_Int_Int_unlockFork6,Go)] */
  logic [5:0] \call_map''_map''_Int_Int_Int_initBuf_emitted ;
  logic [5:0] \call_map''_map''_Int_Int_Int_initBuf_done ;
  assign \call_map''_map''_Int_Int_Int_unlockFork1_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork2_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [1]));
  assign \call_map''_map''_Int_Int_Int_unlockFork3_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [2]));
  assign \call_map''_map''_Int_Int_Int_unlockFork4_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [3]));
  assign \call_map''_map''_Int_Int_Int_unlockFork5_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [4]));
  assign \call_map''_map''_Int_Int_Int_unlockFork6_d  = (\call_map''_map''_Int_Int_Int_initBuf_d [0] && (! \call_map''_map''_Int_Int_Int_initBuf_emitted [5]));
  assign \call_map''_map''_Int_Int_Int_initBuf_done  = (\call_map''_map''_Int_Int_Int_initBuf_emitted  | ({\call_map''_map''_Int_Int_Int_unlockFork6_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork5_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork4_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork3_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork2_d [0],
                                                                                                           \call_map''_map''_Int_Int_Int_unlockFork1_d [0]} & {\call_map''_map''_Int_Int_Int_unlockFork6_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork5_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork4_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork3_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork2_r ,
                                                                                                                                                               \call_map''_map''_Int_Int_Int_unlockFork1_r }));
  assign \call_map''_map''_Int_Int_Int_initBuf_r  = (& \call_map''_map''_Int_Int_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_initBuf_emitted  <= 6'd0;
    else
      \call_map''_map''_Int_Int_Int_initBuf_emitted  <= (\call_map''_map''_Int_Int_Int_initBuf_r  ? 6'd0 :
                                                         \call_map''_map''_Int_Int_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_map''_map''_Int_Int_Int_initBufi,Go) > (call_map''_map''_Int_Int_Int_initBuf,Go) */
  assign \call_map''_map''_Int_Int_Int_initBufi_r  = ((! \call_map''_map''_Int_Int_Int_initBuf_d [0]) || \call_map''_map''_Int_Int_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Int_Int_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_map''_map''_Int_Int_Int_initBufi_r )
        \call_map''_map''_Int_Int_Int_initBuf_d  <= \call_map''_map''_Int_Int_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_map''_map''_Int_Int_Int_unlockFork1,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11,Go)] > (call_map''_map''_Int_Int_Int_goMux1,Go) */
  assign \call_map''_map''_Int_Int_Int_goMux1_d  = (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_r  = (\call_map''_map''_Int_Int_Int_goMux1_r  && (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork1_r  = (\call_map''_map''_Int_Int_Int_goMux1_r  && (\call_map''_map''_Int_Int_Int_unlockFork1_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intgo_11_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_map''_map''_Int_Int_Int_unlockFork2,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC,MyDTInt_Bool)] > (call_map''_map''_Int_Int_Int_goMux2,MyDTInt_Bool) */
  assign \call_map''_map''_Int_Int_Int_goMux2_d  = (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_r  = (\call_map''_map''_Int_Int_Int_goMux2_r  && (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork2_r  = (\call_map''_map''_Int_Int_Int_goMux2_r  && (\call_map''_map''_Int_Int_Int_unlockFork2_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntisZacC_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_map''_map''_Int_Int_Int_unlockFork3,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD,MyDTInt_Int_Int)] > (call_map''_map''_Int_Int_Int_goMux3,MyDTInt_Int_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux3_d  = (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d [0]);
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_r  = (\call_map''_map''_Int_Int_Int_goMux3_r  && (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork3_r  = (\call_map''_map''_Int_Int_Int_goMux3_r  && (\call_map''_map''_Int_Int_Int_unlockFork3_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntgacD_d [0]));
  
  /* mux (Ty Go,
     Ty Int) : (call_map''_map''_Int_Int_Int_unlockFork4,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE,Int)] > (call_map''_map''_Int_Int_Int_goMux4,Int) */
  assign \call_map''_map''_Int_Int_Int_goMux4_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d [32:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_r  = (\call_map''_map''_Int_Int_Int_goMux4_r  && (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork4_r  = (\call_map''_map''_Int_Int_Int_goMux4_r  && (\call_map''_map''_Int_Int_Int_unlockFork4_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intv'acE_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_map''_map''_Int_Int_Int_unlockFork5,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF,Pointer_QTree_Int)] > (call_map''_map''_Int_Int_Int_goMux5,Pointer_QTree_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux5_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d [16:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_r  = (\call_map''_map''_Int_Int_Int_goMux5_r  && (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork5_r  = (\call_map''_map''_Int_Int_Int_goMux5_r  && (\call_map''_map''_Int_Int_Int_unlockFork5_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_IntmacF_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (call_map''_map''_Int_Int_Int_unlockFork6,Go) [(call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3,Pointer_CTmap''_map''_Int_Int_Int)] > (call_map''_map''_Int_Int_Int_goMux6,Pointer_CTmap''_map''_Int_Int_Int) */
  assign \call_map''_map''_Int_Int_Int_goMux6_d  = {\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [16:1],
                                                    (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0])};
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_r  = (\call_map''_map''_Int_Int_Int_goMux6_r  && (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0]));
  assign \call_map''_map''_Int_Int_Int_unlockFork6_r  = (\call_map''_map''_Int_Int_Int_goMux6_r  && (\call_map''_map''_Int_Int_Int_unlockFork6_d [0] && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Intsc_0_3_d [0]));
  
  /* buf (Ty Int) : (es_0_1_1I#_mux_mux_mux,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t \es_0_1_1I#_mux_mux_mux_bufchan_d ;
  logic \es_0_1_1I#_mux_mux_mux_bufchan_r ;
  assign \es_0_1_1I#_mux_mux_mux_r  = ((! \es_0_1_1I#_mux_mux_mux_bufchan_d [0]) || \es_0_1_1I#_mux_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_1_1I#_mux_mux_mux_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\es_0_1_1I#_mux_mux_mux_r )
        \es_0_1_1I#_mux_mux_mux_bufchan_d  <= \es_0_1_1I#_mux_mux_mux_d ;
  Int_t \es_0_1_1I#_mux_mux_mux_bufchan_buf ;
  assign \es_0_1_1I#_mux_mux_mux_bufchan_r  = (! \es_0_1_1I#_mux_mux_mux_bufchan_buf [0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (\es_0_1_1I#_mux_mux_mux_bufchan_buf [0] ? \es_0_1_1I#_mux_mux_mux_bufchan_buf  :
                                          \es_0_1_1I#_mux_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && \es_0_1_1I#_mux_mux_mux_bufchan_buf [0]))
        \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! \es_0_1_1I#_mux_mux_mux_bufchan_buf [0])))
        \es_0_1_1I#_mux_mux_mux_bufchan_buf  <= \es_0_1_1I#_mux_mux_mux_bufchan_d ;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_2_1,MyBool) (lizzieLet17_4QVal_Int_2,Go) > [(es_0_2_1MyFalse,Go),
                                                                  (es_0_2_1MyTrue,Go)] */
  logic [1:0] lizzieLet17_4QVal_Int_2_onehotd;
  always_comb
    if ((es_0_2_1_d[0] && lizzieLet17_4QVal_Int_2_d[0]))
      unique case (es_0_2_1_d[1:1])
        1'd0: lizzieLet17_4QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet17_4QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet17_4QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet17_4QVal_Int_2_onehotd = 2'd0;
  assign es_0_2_1MyFalse_d = lizzieLet17_4QVal_Int_2_onehotd[0];
  assign es_0_2_1MyTrue_d = lizzieLet17_4QVal_Int_2_onehotd[1];
  assign lizzieLet17_4QVal_Int_2_r = (| (lizzieLet17_4QVal_Int_2_onehotd & {es_0_2_1MyTrue_r,
                                                                            es_0_2_1MyFalse_r}));
  assign es_0_2_1_r = lizzieLet17_4QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_0_2_1MyFalse,Go) > (es_0_2_1MyFalse_1_argbuf,Go) */
  Go_t es_0_2_1MyFalse_bufchan_d;
  logic es_0_2_1MyFalse_bufchan_r;
  assign es_0_2_1MyFalse_r = ((! es_0_2_1MyFalse_bufchan_d[0]) || es_0_2_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_2_1MyFalse_r)
        es_0_2_1MyFalse_bufchan_d <= es_0_2_1MyFalse_d;
  Go_t es_0_2_1MyFalse_bufchan_buf;
  assign es_0_2_1MyFalse_bufchan_r = (! es_0_2_1MyFalse_bufchan_buf[0]);
  assign es_0_2_1MyFalse_1_argbuf_d = (es_0_2_1MyFalse_bufchan_buf[0] ? es_0_2_1MyFalse_bufchan_buf :
                                       es_0_2_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_2_1MyFalse_1_argbuf_r && es_0_2_1MyFalse_bufchan_buf[0]))
        es_0_2_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_2_1MyFalse_1_argbuf_r) && (! es_0_2_1MyFalse_bufchan_buf[0])))
        es_0_2_1MyFalse_bufchan_buf <= es_0_2_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_2_1MyTrue,Go) > [(es_0_2_1MyTrue_1,Go),
                                      (es_0_2_1MyTrue_2,Go)] */
  logic [1:0] es_0_2_1MyTrue_emitted;
  logic [1:0] es_0_2_1MyTrue_done;
  assign es_0_2_1MyTrue_1_d = (es_0_2_1MyTrue_d[0] && (! es_0_2_1MyTrue_emitted[0]));
  assign es_0_2_1MyTrue_2_d = (es_0_2_1MyTrue_d[0] && (! es_0_2_1MyTrue_emitted[1]));
  assign es_0_2_1MyTrue_done = (es_0_2_1MyTrue_emitted | ({es_0_2_1MyTrue_2_d[0],
                                                           es_0_2_1MyTrue_1_d[0]} & {es_0_2_1MyTrue_2_r,
                                                                                     es_0_2_1MyTrue_1_r}));
  assign es_0_2_1MyTrue_r = (& es_0_2_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_emitted <= 2'd0;
    else
      es_0_2_1MyTrue_emitted <= (es_0_2_1MyTrue_r ? 2'd0 :
                                 es_0_2_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_0_2_1MyTrue_1,Go)] > (es_0_2_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_0_2_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_0_2_1MyTrue_1_d[0]}), es_0_2_1MyTrue_1_d);
  assign {es_0_2_1MyTrue_1_r} = {1 {(es_0_2_1MyTrue_1QNone_Int_r && es_0_2_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_2_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet20_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_2_1MyTrue_1QNone_Int_bufchan_d;
  logic es_0_2_1MyTrue_1QNone_Int_bufchan_r;
  assign es_0_2_1MyTrue_1QNone_Int_r = ((! es_0_2_1MyTrue_1QNone_Int_bufchan_d[0]) || es_0_2_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_2_1MyTrue_1QNone_Int_r)
        es_0_2_1MyTrue_1QNone_Int_bufchan_d <= es_0_2_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_0_2_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_0_2_1MyTrue_1QNone_Int_bufchan_r = (! es_0_2_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (es_0_2_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_0_2_1MyTrue_1QNone_Int_bufchan_buf :
                                   es_0_2_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && es_0_2_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_0_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! es_0_2_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_0_2_1MyTrue_1QNone_Int_bufchan_buf <= es_0_2_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_0_2_1MyTrue_2,Go) > (es_0_2_1MyTrue_2_argbuf,Go) */
  Go_t es_0_2_1MyTrue_2_bufchan_d;
  logic es_0_2_1MyTrue_2_bufchan_r;
  assign es_0_2_1MyTrue_2_r = ((! es_0_2_1MyTrue_2_bufchan_d[0]) || es_0_2_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_2_1MyTrue_2_r)
        es_0_2_1MyTrue_2_bufchan_d <= es_0_2_1MyTrue_2_d;
  Go_t es_0_2_1MyTrue_2_bufchan_buf;
  assign es_0_2_1MyTrue_2_bufchan_r = (! es_0_2_1MyTrue_2_bufchan_buf[0]);
  assign es_0_2_1MyTrue_2_argbuf_d = (es_0_2_1MyTrue_2_bufchan_buf[0] ? es_0_2_1MyTrue_2_bufchan_buf :
                                      es_0_2_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_2_1MyTrue_2_argbuf_r && es_0_2_1MyTrue_2_bufchan_buf[0]))
        es_0_2_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_2_1MyTrue_2_argbuf_r) && (! es_0_2_1MyTrue_2_bufchan_buf[0])))
        es_0_2_1MyTrue_2_bufchan_buf <= es_0_2_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_2_2,MyBool) (lizzieLet17_6QVal_Int,Pointer_CTmap''_map''_Int_Int_Int) > [(es_0_2_2MyFalse,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                              (es_0_2_2MyTrue,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [1:0] lizzieLet17_6QVal_Int_onehotd;
  always_comb
    if ((es_0_2_2_d[0] && lizzieLet17_6QVal_Int_d[0]))
      unique case (es_0_2_2_d[1:1])
        1'd0: lizzieLet17_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_6QVal_Int_onehotd = 2'd0;
  assign es_0_2_2MyFalse_d = {lizzieLet17_6QVal_Int_d[16:1],
                              lizzieLet17_6QVal_Int_onehotd[0]};
  assign es_0_2_2MyTrue_d = {lizzieLet17_6QVal_Int_d[16:1],
                             lizzieLet17_6QVal_Int_onehotd[1]};
  assign lizzieLet17_6QVal_Int_r = (| (lizzieLet17_6QVal_Int_onehotd & {es_0_2_2MyTrue_r,
                                                                        es_0_2_2MyFalse_r}));
  assign es_0_2_2_r = lizzieLet17_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_2_2MyFalse,Pointer_CTmap''_map''_Int_Int_Int) > (es_0_2_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyFalse_bufchan_d;
  logic es_0_2_2MyFalse_bufchan_r;
  assign es_0_2_2MyFalse_r = ((! es_0_2_2MyFalse_bufchan_d[0]) || es_0_2_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_2_2MyFalse_r)
        es_0_2_2MyFalse_bufchan_d <= es_0_2_2MyFalse_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyFalse_bufchan_buf;
  assign es_0_2_2MyFalse_bufchan_r = (! es_0_2_2MyFalse_bufchan_buf[0]);
  assign es_0_2_2MyFalse_1_argbuf_d = (es_0_2_2MyFalse_bufchan_buf[0] ? es_0_2_2MyFalse_bufchan_buf :
                                       es_0_2_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_2_2MyFalse_1_argbuf_r && es_0_2_2MyFalse_bufchan_buf[0]))
        es_0_2_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_2_2MyFalse_1_argbuf_r) && (! es_0_2_2MyFalse_bufchan_buf[0])))
        es_0_2_2MyFalse_bufchan_buf <= es_0_2_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (es_0_2_2MyTrue,Pointer_CTmap''_map''_Int_Int_Int) > (es_0_2_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyTrue_bufchan_d;
  logic es_0_2_2MyTrue_bufchan_r;
  assign es_0_2_2MyTrue_r = ((! es_0_2_2MyTrue_bufchan_d[0]) || es_0_2_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_2_2MyTrue_r) es_0_2_2MyTrue_bufchan_d <= es_0_2_2MyTrue_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  es_0_2_2MyTrue_bufchan_buf;
  assign es_0_2_2MyTrue_bufchan_r = (! es_0_2_2MyTrue_bufchan_buf[0]);
  assign es_0_2_2MyTrue_1_argbuf_d = (es_0_2_2MyTrue_bufchan_buf[0] ? es_0_2_2MyTrue_bufchan_buf :
                                      es_0_2_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_2_2MyTrue_1_argbuf_r && es_0_2_2MyTrue_bufchan_buf[0]))
        es_0_2_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_2_2MyTrue_1_argbuf_r) && (! es_0_2_2MyTrue_bufchan_buf[0])))
        es_0_2_2MyTrue_bufchan_buf <= es_0_2_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_0_2_3,MyBool) (xac0_2,Int) > [(es_0_2_3MyFalse,Int),
                                                   (_48,Int)] */
  logic [1:0] xac0_2_onehotd;
  always_comb
    if ((es_0_2_3_d[0] && xac0_2_d[0]))
      unique case (es_0_2_3_d[1:1])
        1'd0: xac0_2_onehotd = 2'd1;
        1'd1: xac0_2_onehotd = 2'd2;
        default: xac0_2_onehotd = 2'd0;
      endcase
    else xac0_2_onehotd = 2'd0;
  assign es_0_2_3MyFalse_d = {xac0_2_d[32:1], xac0_2_onehotd[0]};
  assign _48_d = {xac0_2_d[32:1], xac0_2_onehotd[1]};
  assign xac0_2_r = (| (xac0_2_onehotd & {_48_r,
                                          es_0_2_3MyFalse_r}));
  assign es_0_2_3_r = xac0_2_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(es_0_2_3MyFalse,Int)] > (es_0_2_3MyFalse_1QVal_Int,QTree_Int) */
  assign es_0_2_3MyFalse_1QVal_Int_d = QVal_Int_dc((& {es_0_2_3MyFalse_d[0]}), es_0_2_3MyFalse_d);
  assign {es_0_2_3MyFalse_r} = {1 {(es_0_2_3MyFalse_1QVal_Int_r && es_0_2_3MyFalse_1QVal_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_0_2_3MyFalse_1QVal_Int,QTree_Int) > (lizzieLet19_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_2_3MyFalse_1QVal_Int_bufchan_d;
  logic es_0_2_3MyFalse_1QVal_Int_bufchan_r;
  assign es_0_2_3MyFalse_1QVal_Int_r = ((! es_0_2_3MyFalse_1QVal_Int_bufchan_d[0]) || es_0_2_3MyFalse_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_3MyFalse_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_2_3MyFalse_1QVal_Int_r)
        es_0_2_3MyFalse_1QVal_Int_bufchan_d <= es_0_2_3MyFalse_1QVal_Int_d;
  QTree_Int_t es_0_2_3MyFalse_1QVal_Int_bufchan_buf;
  assign es_0_2_3MyFalse_1QVal_Int_bufchan_r = (! es_0_2_3MyFalse_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (es_0_2_3MyFalse_1QVal_Int_bufchan_buf[0] ? es_0_2_3MyFalse_1QVal_Int_bufchan_buf :
                                   es_0_2_3MyFalse_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && es_0_2_3MyFalse_1QVal_Int_bufchan_buf[0]))
        es_0_2_3MyFalse_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! es_0_2_3MyFalse_1QVal_Int_bufchan_buf[0])))
        es_0_2_3MyFalse_1QVal_Int_bufchan_buf <= es_0_2_3MyFalse_1QVal_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  logic es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_r;
  assign es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_r = ((! es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d[0]) || es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= {32'd0,
                                                                  1'd0};
    else
      if (es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_r)
        es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_d;
  \Int#_t  es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf;
  assign es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_r = (! es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0] ? es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf :
                                 es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                    1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]))
        es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                      1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0])))
        es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_1ww2XyF_1_1_Add32,Int#) (lizzieLet26_4Lcall_$wnnz_Int0,Int#) > (es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32,Int#) */
  assign es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_d = {(es_6_1ww2XyF_1_1_Add32_d[32:1] + lizzieLet26_4Lcall_$wnnz_Int0_d[32:1]),
                                                            (es_6_1ww2XyF_1_1_Add32_d[0] && lizzieLet26_4Lcall_$wnnz_Int0_d[0])};
  assign {es_6_1ww2XyF_1_1_Add32_r,
          lizzieLet26_4Lcall_$wnnz_Int0_r} = {2 {(es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_r && es_4_1_1lizzieLet26_4Lcall_$wnnz_Int0_1_Add32_d[0])}};
  
  /* sink (Ty Int) : (es_7_1I#,Int) > */
  assign {\es_7_1I#_r , \es_7_1I#_dout } = {\es_7_1I#_rout ,
                                            \es_7_1I#_d };
  
  /* buf (Ty MyDTInt_Int_Int) : (gacD_2_2,MyDTInt_Int_Int) > (gacD_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacD_2_2_bufchan_d;
  logic gacD_2_2_bufchan_r;
  assign gacD_2_2_r = ((! gacD_2_2_bufchan_d[0]) || gacD_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_2_2_bufchan_d <= 1'd0;
    else if (gacD_2_2_r) gacD_2_2_bufchan_d <= gacD_2_2_d;
  MyDTInt_Int_Int_t gacD_2_2_bufchan_buf;
  assign gacD_2_2_bufchan_r = (! gacD_2_2_bufchan_buf[0]);
  assign gacD_2_2_argbuf_d = (gacD_2_2_bufchan_buf[0] ? gacD_2_2_bufchan_buf :
                              gacD_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacD_2_2_argbuf_r && gacD_2_2_bufchan_buf[0]))
        gacD_2_2_bufchan_buf <= 1'd0;
      else if (((! gacD_2_2_argbuf_r) && (! gacD_2_2_bufchan_buf[0])))
        gacD_2_2_bufchan_buf <= gacD_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacD_2_destruct,MyDTInt_Int_Int) > [(gacD_2_1,MyDTInt_Int_Int),
                                                                 (gacD_2_2,MyDTInt_Int_Int)] */
  logic [1:0] gacD_2_destruct_emitted;
  logic [1:0] gacD_2_destruct_done;
  assign gacD_2_1_d = (gacD_2_destruct_d[0] && (! gacD_2_destruct_emitted[0]));
  assign gacD_2_2_d = (gacD_2_destruct_d[0] && (! gacD_2_destruct_emitted[1]));
  assign gacD_2_destruct_done = (gacD_2_destruct_emitted | ({gacD_2_2_d[0],
                                                             gacD_2_1_d[0]} & {gacD_2_2_r,
                                                                               gacD_2_1_r}));
  assign gacD_2_destruct_r = (& gacD_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_2_destruct_emitted <= 2'd0;
    else
      gacD_2_destruct_emitted <= (gacD_2_destruct_r ? 2'd0 :
                                  gacD_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacD_3_2,MyDTInt_Int_Int) > (gacD_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacD_3_2_bufchan_d;
  logic gacD_3_2_bufchan_r;
  assign gacD_3_2_r = ((! gacD_3_2_bufchan_d[0]) || gacD_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_3_2_bufchan_d <= 1'd0;
    else if (gacD_3_2_r) gacD_3_2_bufchan_d <= gacD_3_2_d;
  MyDTInt_Int_Int_t gacD_3_2_bufchan_buf;
  assign gacD_3_2_bufchan_r = (! gacD_3_2_bufchan_buf[0]);
  assign gacD_3_2_argbuf_d = (gacD_3_2_bufchan_buf[0] ? gacD_3_2_bufchan_buf :
                              gacD_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacD_3_2_argbuf_r && gacD_3_2_bufchan_buf[0]))
        gacD_3_2_bufchan_buf <= 1'd0;
      else if (((! gacD_3_2_argbuf_r) && (! gacD_3_2_bufchan_buf[0])))
        gacD_3_2_bufchan_buf <= gacD_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacD_3_destruct,MyDTInt_Int_Int) > [(gacD_3_1,MyDTInt_Int_Int),
                                                                 (gacD_3_2,MyDTInt_Int_Int)] */
  logic [1:0] gacD_3_destruct_emitted;
  logic [1:0] gacD_3_destruct_done;
  assign gacD_3_1_d = (gacD_3_destruct_d[0] && (! gacD_3_destruct_emitted[0]));
  assign gacD_3_2_d = (gacD_3_destruct_d[0] && (! gacD_3_destruct_emitted[1]));
  assign gacD_3_destruct_done = (gacD_3_destruct_emitted | ({gacD_3_2_d[0],
                                                             gacD_3_1_d[0]} & {gacD_3_2_r,
                                                                               gacD_3_1_r}));
  assign gacD_3_destruct_r = (& gacD_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_3_destruct_emitted <= 2'd0;
    else
      gacD_3_destruct_emitted <= (gacD_3_destruct_r ? 2'd0 :
                                  gacD_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacD_4_destruct,MyDTInt_Int_Int) > (gacD_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacD_4_destruct_bufchan_d;
  logic gacD_4_destruct_bufchan_r;
  assign gacD_4_destruct_r = ((! gacD_4_destruct_bufchan_d[0]) || gacD_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacD_4_destruct_r)
        gacD_4_destruct_bufchan_d <= gacD_4_destruct_d;
  MyDTInt_Int_Int_t gacD_4_destruct_bufchan_buf;
  assign gacD_4_destruct_bufchan_r = (! gacD_4_destruct_bufchan_buf[0]);
  assign gacD_4_1_argbuf_d = (gacD_4_destruct_bufchan_buf[0] ? gacD_4_destruct_bufchan_buf :
                              gacD_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacD_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacD_4_1_argbuf_r && gacD_4_destruct_bufchan_buf[0]))
        gacD_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacD_4_1_argbuf_r) && (! gacD_4_destruct_bufchan_buf[0])))
        gacD_4_destruct_bufchan_buf <= gacD_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (gacM_2_2,MyDTInt_Int_Int) > (gacM_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacM_2_2_bufchan_d;
  logic gacM_2_2_bufchan_r;
  assign gacM_2_2_r = ((! gacM_2_2_bufchan_d[0]) || gacM_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_2_bufchan_d <= 1'd0;
    else if (gacM_2_2_r) gacM_2_2_bufchan_d <= gacM_2_2_d;
  MyDTInt_Int_Int_t gacM_2_2_bufchan_buf;
  assign gacM_2_2_bufchan_r = (! gacM_2_2_bufchan_buf[0]);
  assign gacM_2_2_argbuf_d = (gacM_2_2_bufchan_buf[0] ? gacM_2_2_bufchan_buf :
                              gacM_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacM_2_2_argbuf_r && gacM_2_2_bufchan_buf[0]))
        gacM_2_2_bufchan_buf <= 1'd0;
      else if (((! gacM_2_2_argbuf_r) && (! gacM_2_2_bufchan_buf[0])))
        gacM_2_2_bufchan_buf <= gacM_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacM_2_destruct,MyDTInt_Int_Int) > [(gacM_2_1,MyDTInt_Int_Int),
                                                                 (gacM_2_2,MyDTInt_Int_Int)] */
  logic [1:0] gacM_2_destruct_emitted;
  logic [1:0] gacM_2_destruct_done;
  assign gacM_2_1_d = (gacM_2_destruct_d[0] && (! gacM_2_destruct_emitted[0]));
  assign gacM_2_2_d = (gacM_2_destruct_d[0] && (! gacM_2_destruct_emitted[1]));
  assign gacM_2_destruct_done = (gacM_2_destruct_emitted | ({gacM_2_2_d[0],
                                                             gacM_2_1_d[0]} & {gacM_2_2_r,
                                                                               gacM_2_1_r}));
  assign gacM_2_destruct_r = (& gacM_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_2_destruct_emitted <= 2'd0;
    else
      gacM_2_destruct_emitted <= (gacM_2_destruct_r ? 2'd0 :
                                  gacM_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacM_3_2,MyDTInt_Int_Int) > (gacM_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacM_3_2_bufchan_d;
  logic gacM_3_2_bufchan_r;
  assign gacM_3_2_r = ((! gacM_3_2_bufchan_d[0]) || gacM_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_2_bufchan_d <= 1'd0;
    else if (gacM_3_2_r) gacM_3_2_bufchan_d <= gacM_3_2_d;
  MyDTInt_Int_Int_t gacM_3_2_bufchan_buf;
  assign gacM_3_2_bufchan_r = (! gacM_3_2_bufchan_buf[0]);
  assign gacM_3_2_argbuf_d = (gacM_3_2_bufchan_buf[0] ? gacM_3_2_bufchan_buf :
                              gacM_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacM_3_2_argbuf_r && gacM_3_2_bufchan_buf[0]))
        gacM_3_2_bufchan_buf <= 1'd0;
      else if (((! gacM_3_2_argbuf_r) && (! gacM_3_2_bufchan_buf[0])))
        gacM_3_2_bufchan_buf <= gacM_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (gacM_3_destruct,MyDTInt_Int_Int) > [(gacM_3_1,MyDTInt_Int_Int),
                                                                 (gacM_3_2,MyDTInt_Int_Int)] */
  logic [1:0] gacM_3_destruct_emitted;
  logic [1:0] gacM_3_destruct_done;
  assign gacM_3_1_d = (gacM_3_destruct_d[0] && (! gacM_3_destruct_emitted[0]));
  assign gacM_3_2_d = (gacM_3_destruct_d[0] && (! gacM_3_destruct_emitted[1]));
  assign gacM_3_destruct_done = (gacM_3_destruct_emitted | ({gacM_3_2_d[0],
                                                             gacM_3_1_d[0]} & {gacM_3_2_r,
                                                                               gacM_3_1_r}));
  assign gacM_3_destruct_r = (& gacM_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_3_destruct_emitted <= 2'd0;
    else
      gacM_3_destruct_emitted <= (gacM_3_destruct_r ? 2'd0 :
                                  gacM_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (gacM_4_destruct,MyDTInt_Int_Int) > (gacM_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t gacM_4_destruct_bufchan_d;
  logic gacM_4_destruct_bufchan_r;
  assign gacM_4_destruct_r = ((! gacM_4_destruct_bufchan_d[0]) || gacM_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacM_4_destruct_r)
        gacM_4_destruct_bufchan_d <= gacM_4_destruct_d;
  MyDTInt_Int_Int_t gacM_4_destruct_bufchan_buf;
  assign gacM_4_destruct_bufchan_r = (! gacM_4_destruct_bufchan_buf[0]);
  assign gacM_4_1_argbuf_d = (gacM_4_destruct_bufchan_buf[0] ? gacM_4_destruct_bufchan_buf :
                              gacM_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacM_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacM_4_1_argbuf_r && gacM_4_destruct_bufchan_buf[0]))
        gacM_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacM_4_1_argbuf_r) && (! gacM_4_destruct_bufchan_buf[0])))
        gacM_4_destruct_bufchan_buf <= gacM_4_destruct_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c*) : [(go_1,Go)] > (go_1Dcon_$fNumInt_$c*,MyDTInt_Int_Int) */
  assign \go_1Dcon_$fNumInt_$ctimes_d  = \Dcon_$fNumInt_$ctimes_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_$fNumInt_$ctimes_r  && \go_1Dcon_$fNumInt_$ctimes_d [0])}};
  
  /* fork (Ty C5) : (go_10_goMux_choice,C5) > [(go_10_goMux_choice_1,C5),
                                          (go_10_goMux_choice_2,C5),
                                          (go_10_goMux_choice_3,C5)] */
  logic [2:0] go_10_goMux_choice_emitted;
  logic [2:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_3_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[2]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_3_d[0],
                                                                   go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_3_r,
                                                                                                 go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 3'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 3'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C5) [(call_main_mask_Int_goMux2,Pointer_QTree_Int),
                                                        (t3act_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2acs_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1acr_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4acu_1_argbuf,Pointer_QTree_Int)] > (mack_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] mack_goMux_mux_mux;
  logic [4:0] mack_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[3:1])
      3'd0:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd1,
                                                       call_main_mask_Int_goMux2_d};
      3'd1:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd2,
                                                       t3act_1_1_argbuf_d};
      3'd2:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd4,
                                                       t2acs_2_1_argbuf_d};
      3'd3:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd8,
                                                       t1acr_3_1_argbuf_d};
      3'd4:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd16,
                                                       t4acu_1_argbuf_d};
      default:
        {mack_goMux_mux_onehot, mack_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign mack_goMux_mux_d = {mack_goMux_mux_mux[16:1],
                             (mack_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (mack_goMux_mux_d[0] && mack_goMux_mux_r);
  assign {t4acu_1_argbuf_r,
          t1acr_3_1_argbuf_r,
          t2acs_2_1_argbuf_r,
          t3act_1_1_argbuf_r,
          call_main_mask_Int_goMux2_r} = (go_10_goMux_choice_1_r ? mack_goMux_mux_onehot :
                                          5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_10_goMux_choice_2,C5) [(call_main_mask_Int_goMux3,Pointer_MaskQTree),
                                                        (q3aco_1_1_argbuf,Pointer_MaskQTree),
                                                        (q2acn_2_1_argbuf,Pointer_MaskQTree),
                                                        (q1acm_3_1_argbuf,Pointer_MaskQTree),
                                                        (lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree)] > (mskacl_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] mskacl_goMux_mux_mux;
  logic [4:0] mskacl_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[3:1])
      3'd0:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Int_goMux3_d};
      3'd1:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd2,
                                                           q3aco_1_1_argbuf_d};
      3'd2:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd4,
                                                           q2acn_2_1_argbuf_d};
      3'd3:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd8,
                                                           q1acm_3_1_argbuf_d};
      3'd4:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd16,
                                                           lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_d};
      default:
        {mskacl_goMux_mux_onehot, mskacl_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign mskacl_goMux_mux_d = {mskacl_goMux_mux_mux[16:1],
                               (mskacl_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (mskacl_goMux_mux_d[0] && mskacl_goMux_mux_r);
  assign {lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_r,
          q1acm_3_1_argbuf_r,
          q2acn_2_1_argbuf_r,
          q3aco_1_1_argbuf_r,
          call_main_mask_Int_goMux3_r} = (go_10_goMux_choice_2_r ? mskacl_goMux_mux_onehot :
                                          5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_mask_Int) : (go_10_goMux_choice_3,C5) [(call_main_mask_Int_goMux4,Pointer_CTmain_mask_Int),
                                                              (sca2_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (sca1_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (sca0_2_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (sca3_2_1_argbuf,Pointer_CTmain_mask_Int)] > (sc_0_2_goMux_mux,Pointer_CTmain_mask_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Int_goMux4_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_10_goMux_choice_3_d[0])};
  assign go_10_goMux_choice_3_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_main_mask_Int_goMux4_r} = (go_10_goMux_choice_3_r ? sc_0_2_goMux_mux_onehot :
                                          5'd0);
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5),
                                          (go_11_goMux_choice_3,C5),
                                          (go_11_goMux_choice_4,C5),
                                          (go_11_goMux_choice_5,C5)] */
  logic [4:0] go_11_goMux_choice_emitted;
  logic [4:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_3_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[2]))};
  assign go_11_goMux_choice_4_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[3]))};
  assign go_11_goMux_choice_5_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[4]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_5_d[0],
                                                                   go_11_goMux_choice_4_d[0],
                                                                   go_11_goMux_choice_3_d[0],
                                                                   go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_5_r,
                                                                                                 go_11_goMux_choice_4_r,
                                                                                                 go_11_goMux_choice_3_r,
                                                                                                 go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 5'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 5'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_11_goMux_choice_1,C5) [(call_map''_map''_Int_Int_Int_goMux2,MyDTInt_Bool),
                                                   (isZacC_2_2_argbuf,MyDTInt_Bool),
                                                   (isZacC_3_2_argbuf,MyDTInt_Bool),
                                                   (isZacC_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet17_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (isZacC_goMux_mux,MyDTInt_Bool) */
  logic [0:0] isZacC_goMux_mux_mux;
  logic [4:0] isZacC_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Int_Int_Int_goMux2_d };
      3'd1:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd2,
                                                           isZacC_2_2_argbuf_d};
      3'd2:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd4,
                                                           isZacC_3_2_argbuf_d};
      3'd3:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd8,
                                                           isZacC_4_1_argbuf_d};
      3'd4:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd16,
                                                           lizzieLet17_5QNode_Int_2_argbuf_d};
      default:
        {isZacC_goMux_mux_onehot, isZacC_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacC_goMux_mux_d = (isZacC_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0]);
  assign go_11_goMux_choice_1_r = (isZacC_goMux_mux_d[0] && isZacC_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_2_argbuf_r,
          isZacC_4_1_argbuf_r,
          isZacC_3_2_argbuf_r,
          isZacC_2_2_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux2_r } = (go_11_goMux_choice_1_r ? isZacC_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_11_goMux_choice_2,C5) [(call_map''_map''_Int_Int_Int_goMux3,MyDTInt_Int_Int),
                                                      (gacD_2_2_argbuf,MyDTInt_Int_Int),
                                                      (gacD_3_2_argbuf,MyDTInt_Int_Int),
                                                      (gacD_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet17_3QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (gacD_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] gacD_goMux_mux_mux;
  logic [4:0] gacD_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Int_Int_Int_goMux3_d };
      3'd1:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd2,
                                                       gacD_2_2_argbuf_d};
      3'd2:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd4,
                                                       gacD_3_2_argbuf_d};
      3'd3:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd8,
                                                       gacD_4_1_argbuf_d};
      3'd4:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd16,
                                                       lizzieLet17_3QNode_Int_2_argbuf_d};
      default:
        {gacD_goMux_mux_onehot, gacD_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacD_goMux_mux_d = (gacD_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0]);
  assign go_11_goMux_choice_2_r = (gacD_goMux_mux_d[0] && gacD_goMux_mux_r);
  assign {lizzieLet17_3QNode_Int_2_argbuf_r,
          gacD_4_1_argbuf_r,
          gacD_3_2_argbuf_r,
          gacD_2_2_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux3_r } = (go_11_goMux_choice_2_r ? gacD_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Int) : (go_11_goMux_choice_3,C5) [(call_map''_map''_Int_Int_Int_goMux4,Int),
                                          (v'acE_2_2_argbuf,Int),
                                          (v'acE_3_2_argbuf,Int),
                                          (v'acE_4_1_argbuf,Int),
                                          (lizzieLet17_7QNode_Int_2_argbuf,Int)] > (v'acE_goMux_mux,Int) */
  logic [32:0] \v'acE_goMux_mux_mux ;
  logic [4:0] \v'acE_goMux_mux_onehot ;
  always_comb
    unique case (go_11_goMux_choice_3_d[3:1])
      3'd0:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd1,
                                                             \call_map''_map''_Int_Int_Int_goMux4_d };
      3'd1:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd2,
                                                             \v'acE_2_2_argbuf_d };
      3'd2:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd4,
                                                             \v'acE_3_2_argbuf_d };
      3'd3:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd8,
                                                             \v'acE_4_1_argbuf_d };
      3'd4:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd16,
                                                             lizzieLet17_7QNode_Int_2_argbuf_d};
      default:
        {\v'acE_goMux_mux_onehot , \v'acE_goMux_mux_mux } = {5'd0,
                                                             {32'd0, 1'd0}};
    endcase
  assign \v'acE_goMux_mux_d  = {\v'acE_goMux_mux_mux [32:1],
                                (\v'acE_goMux_mux_mux [0] && go_11_goMux_choice_3_d[0])};
  assign go_11_goMux_choice_3_r = (\v'acE_goMux_mux_d [0] && \v'acE_goMux_mux_r );
  assign {lizzieLet17_7QNode_Int_2_argbuf_r,
          \v'acE_4_1_argbuf_r ,
          \v'acE_3_2_argbuf_r ,
          \v'acE_2_2_argbuf_r ,
          \call_map''_map''_Int_Int_Int_goMux4_r } = (go_11_goMux_choice_3_r ? \v'acE_goMux_mux_onehot  :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_4,C5) [(call_map''_map''_Int_Int_Int_goMux5,Pointer_QTree_Int),
                                                        (q3acJ_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2acI_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1acH_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4acK_1_argbuf,Pointer_QTree_Int)] > (macF_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] macF_goMux_mux_mux;
  logic [4:0] macF_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_4_d[3:1])
      3'd0:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Int_Int_Int_goMux5_d };
      3'd1:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd2,
                                                       q3acJ_1_1_argbuf_d};
      3'd2:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd4,
                                                       q2acI_2_1_argbuf_d};
      3'd3:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd8,
                                                       q1acH_3_1_argbuf_d};
      3'd4:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd16,
                                                       q4acK_1_argbuf_d};
      default:
        {macF_goMux_mux_onehot, macF_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign macF_goMux_mux_d = {macF_goMux_mux_mux[16:1],
                             (macF_goMux_mux_mux[0] && go_11_goMux_choice_4_d[0])};
  assign go_11_goMux_choice_4_r = (macF_goMux_mux_d[0] && macF_goMux_mux_r);
  assign {q4acK_1_argbuf_r,
          q1acH_3_1_argbuf_r,
          q2acI_2_1_argbuf_r,
          q3acJ_1_1_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux5_r } = (go_11_goMux_choice_4_r ? macF_goMux_mux_onehot :
                                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (go_11_goMux_choice_5,C5) [(call_map''_map''_Int_Int_Int_goMux6,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca2_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca1_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sca3_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (sc_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) */
  logic [16:0] sc_0_3_goMux_mux_mux;
  logic [4:0] sc_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Int_Int_Int_goMux6_d };
      3'd1:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd2,
                                                           sca2_3_1_argbuf_d};
      3'd2:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd4,
                                                           sca1_3_1_argbuf_d};
      3'd3:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd8,
                                                           sca0_3_1_argbuf_d};
      3'd4:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd16,
                                                           sca3_3_1_argbuf_d};
      default:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_3_goMux_mux_d = {sc_0_3_goMux_mux_mux[16:1],
                               (sc_0_3_goMux_mux_mux[0] && go_11_goMux_choice_5_d[0])};
  assign go_11_goMux_choice_5_r = (sc_0_3_goMux_mux_d[0] && sc_0_3_goMux_mux_r);
  assign {sca3_3_1_argbuf_r,
          sca0_3_1_argbuf_r,
          sca1_3_1_argbuf_r,
          sca2_3_1_argbuf_r,
          \call_map''_map''_Int_Int_Int_goMux6_r } = (go_11_goMux_choice_5_r ? sc_0_3_goMux_mux_onehot :
                                                      5'd0);
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lkron_kron_Int_Int_Intsbos) : [(go_12_1,Go)] > (go_12_1Lkron_kron_Int_Int_Intsbos,CTkron_kron_Int_Int_Int) */
  assign go_12_1Lkron_kron_Int_Int_Intsbos_d = Lkron_kron_Int_Int_Intsbos_dc((& {go_12_1_d[0]}), go_12_1_d);
  assign {go_12_1_r} = {1 {(go_12_1Lkron_kron_Int_Int_Intsbos_r && go_12_1Lkron_kron_Int_Int_Intsbos_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (go_12_1Lkron_kron_Int_Int_Intsbos,CTkron_kron_Int_Int_Int) > (lizzieLet23_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d;
  logic go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_r;
  assign go_12_1Lkron_kron_Int_Int_Intsbos_r = ((! go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d[0]) || go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d <= {83'd0, 1'd0};
    else
      if (go_12_1Lkron_kron_Int_Int_Intsbos_r)
        go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d <= go_12_1Lkron_kron_Int_Int_Intsbos_d;
  CTkron_kron_Int_Int_Int_t go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf;
  assign go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_r = (! go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0] ? go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf :
                                   go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0]))
        go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf[0])))
        go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_buf <= go_12_1Lkron_kron_Int_Int_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_12_2,Go) > (go_12_2_argbuf,Go) */
  Go_t go_12_2_bufchan_d;
  logic go_12_2_bufchan_r;
  assign go_12_2_r = ((! go_12_2_bufchan_d[0]) || go_12_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_d <= 1'd0;
    else if (go_12_2_r) go_12_2_bufchan_d <= go_12_2_d;
  Go_t go_12_2_bufchan_buf;
  assign go_12_2_bufchan_r = (! go_12_2_bufchan_buf[0]);
  assign go_12_2_argbuf_d = (go_12_2_bufchan_buf[0] ? go_12_2_bufchan_buf :
                             go_12_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_buf <= 1'd0;
    else
      if ((go_12_2_argbuf_r && go_12_2_bufchan_buf[0]))
        go_12_2_bufchan_buf <= 1'd0;
      else if (((! go_12_2_argbuf_r) && (! go_12_2_bufchan_buf[0])))
        go_12_2_bufchan_buf <= go_12_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) : [(go_12_2_argbuf,Go),
                                                                                                                                (isZacL_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                (gacM_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                (m1acN_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                (m2acO_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                (lizzieLet13_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int) */
  assign call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_dc((& {go_12_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                  isZacL_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  gacM_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  m1acN_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  m2acO_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                  lizzieLet13_1_1_argbuf_d[0]}), go_12_2_argbuf_d, isZacL_1_1_argbuf_d, gacM_1_1_argbuf_d, m1acN_1_1_argbuf_d, m2acO_1_1_argbuf_d, lizzieLet13_1_1_argbuf_d);
  assign {go_12_2_argbuf_r,
          isZacL_1_1_argbuf_r,
          gacM_1_1_argbuf_r,
          m1acN_1_1_argbuf_r,
          m2acO_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r} = {6 {(call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_r && call_kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTkron_kron_Int_Int_Int_1_d[0])}};
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lmain_mask_Intsbos) : [(go_13_1,Go)] > (go_13_1Lmain_mask_Intsbos,CTmain_mask_Int) */
  assign go_13_1Lmain_mask_Intsbos_d = Lmain_mask_Intsbos_dc((& {go_13_1_d[0]}), go_13_1_d);
  assign {go_13_1_r} = {1 {(go_13_1Lmain_mask_Intsbos_r && go_13_1Lmain_mask_Intsbos_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (go_13_1Lmain_mask_Intsbos,CTmain_mask_Int) > (lizzieLet24_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t go_13_1Lmain_mask_Intsbos_bufchan_d;
  logic go_13_1Lmain_mask_Intsbos_bufchan_r;
  assign go_13_1Lmain_mask_Intsbos_r = ((! go_13_1Lmain_mask_Intsbos_bufchan_d[0]) || go_13_1Lmain_mask_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_13_1Lmain_mask_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_13_1Lmain_mask_Intsbos_r)
        go_13_1Lmain_mask_Intsbos_bufchan_d <= go_13_1Lmain_mask_Intsbos_d;
  CTmain_mask_Int_t go_13_1Lmain_mask_Intsbos_bufchan_buf;
  assign go_13_1Lmain_mask_Intsbos_bufchan_r = (! go_13_1Lmain_mask_Intsbos_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (go_13_1Lmain_mask_Intsbos_bufchan_buf[0] ? go_13_1Lmain_mask_Intsbos_bufchan_buf :
                                   go_13_1Lmain_mask_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_13_1Lmain_mask_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && go_13_1Lmain_mask_Intsbos_bufchan_buf[0]))
        go_13_1Lmain_mask_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! go_13_1Lmain_mask_Intsbos_bufchan_buf[0])))
        go_13_1Lmain_mask_Intsbos_bufchan_buf <= go_13_1Lmain_mask_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_13_2,Go) > (go_13_2_argbuf,Go) */
  Go_t go_13_2_bufchan_d;
  logic go_13_2_bufchan_r;
  assign go_13_2_r = ((! go_13_2_bufchan_d[0]) || go_13_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_d <= 1'd0;
    else if (go_13_2_r) go_13_2_bufchan_d <= go_13_2_d;
  Go_t go_13_2_bufchan_buf;
  assign go_13_2_bufchan_r = (! go_13_2_bufchan_buf[0]);
  assign go_13_2_argbuf_d = (go_13_2_bufchan_buf[0] ? go_13_2_bufchan_buf :
                             go_13_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_buf <= 1'd0;
    else
      if ((go_13_2_argbuf_r && go_13_2_bufchan_buf[0]))
        go_13_2_bufchan_buf <= 1'd0;
      else if (((! go_13_2_argbuf_r) && (! go_13_2_bufchan_buf[0])))
        go_13_2_bufchan_buf <= go_13_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) : [(go_13_2_argbuf,Go),
                                                                                       (mack_1_1_argbuf,Pointer_QTree_Int),
                                                                                       (mskacl_1_1_argbuf,Pointer_MaskQTree),
                                                                                       (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Int)] > (call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int) */
  assign call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_dc((& {go_13_2_argbuf_d[0],
                                                                                                                                                                                        mack_1_1_argbuf_d[0],
                                                                                                                                                                                        mskacl_1_1_argbuf_d[0],
                                                                                                                                                                                        lizzieLet4_1_1_argbuf_d[0]}), go_13_2_argbuf_d, mack_1_1_argbuf_d, mskacl_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_13_2_argbuf_r,
          mack_1_1_argbuf_r,
          mskacl_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {4 {(call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_r && call_main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree___Pointer_CTmain_mask_Int_1_d[0])}};
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lmap''_map''_Int_Int_Intsbos) : [(go_14_1,Go)] > (go_14_1Lmap''_map''_Int_Int_Intsbos,CTmap''_map''_Int_Int_Int) */
  assign \go_14_1Lmap''_map''_Int_Int_Intsbos_d  = \Lmap''_map''_Int_Int_Intsbos_dc ((& {go_14_1_d[0]}), go_14_1_d);
  assign {go_14_1_r} = {1 {(\go_14_1Lmap''_map''_Int_Int_Intsbos_r  && \go_14_1Lmap''_map''_Int_Int_Intsbos_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (go_14_1Lmap''_map''_Int_Int_Intsbos,CTmap''_map''_Int_Int_Int) > (lizzieLet25_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d ;
  logic \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_r ;
  assign \go_14_1Lmap''_map''_Int_Int_Intsbos_r  = ((! \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d [0]) || \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d  <= {99'd0, 1'd0};
    else
      if (\go_14_1Lmap''_map''_Int_Int_Intsbos_r )
        \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d  <= \go_14_1Lmap''_map''_Int_Int_Intsbos_d ;
  \CTmap''_map''_Int_Int_Int_t  \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf ;
  assign \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_r  = (! \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0]);
  assign lizzieLet25_1_argbuf_d = (\go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0] ? \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  :
                                   \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0]))
        \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf [0])))
        \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_buf  <= \go_14_1Lmap''_map''_Int_Int_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_14_2,Go) > (go_14_2_argbuf,Go) */
  Go_t go_14_2_bufchan_d;
  logic go_14_2_bufchan_r;
  assign go_14_2_r = ((! go_14_2_bufchan_d[0]) || go_14_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_d <= 1'd0;
    else if (go_14_2_r) go_14_2_bufchan_d <= go_14_2_d;
  Go_t go_14_2_bufchan_buf;
  assign go_14_2_bufchan_r = (! go_14_2_bufchan_buf[0]);
  assign go_14_2_argbuf_d = (go_14_2_bufchan_buf[0] ? go_14_2_bufchan_buf :
                             go_14_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_buf <= 1'd0;
    else
      if ((go_14_2_argbuf_r && go_14_2_bufchan_buf[0]))
        go_14_2_bufchan_buf <= 1'd0;
      else if (((! go_14_2_argbuf_r) && (! go_14_2_bufchan_buf[0])))
        go_14_2_bufchan_buf <= go_14_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) : [(go_14_2_argbuf,Go),
                                                                                                                    (isZacC_1_1_argbuf,MyDTInt_Bool),
                                                                                                                    (gacD_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                    (v'acE_1_1_argbuf,Int),
                                                                                                                    (macF_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                    (lizzieLet9_1_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int) */
  assign \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d  = \TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_dc ((& {go_14_2_argbuf_d[0],
                                                                                                                                                                                                                                                                isZacC_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                gacD_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                \v'acE_1_1_argbuf_d [0],
                                                                                                                                                                                                                                                                macF_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                lizzieLet9_1_1_argbuf_d[0]}), go_14_2_argbuf_d, isZacC_1_1_argbuf_d, gacD_1_1_argbuf_d, \v'acE_1_1_argbuf_d , macF_1_1_argbuf_d, lizzieLet9_1_1_argbuf_d);
  assign {go_14_2_argbuf_r,
          isZacC_1_1_argbuf_r,
          gacD_1_1_argbuf_r,
          \v'acE_1_1_argbuf_r ,
          macF_1_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r} = {6 {(\call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_r  && \call_map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int___Pointer_CTmap''_map''_Int_Int_Int_1_d [0])}};
  
  /* fork (Ty C4) : (go_15_goMux_choice,C4) > [(go_15_goMux_choice_1,C4),
                                          (go_15_goMux_choice_2,C4)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_15_goMux_choice_1,C4) [(lizzieLet14_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet15_1_argbuf,Int#),
                                           (lizzieLet14_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet14_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet15_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet14_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet14_1_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet14_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz_Int) : (go_15_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_7_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_7_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C4) : (go_16_goMux_choice,C4) > [(go_16_goMux_choice_1,C4),
                                          (go_16_goMux_choice_2,C4)] */
  logic [1:0] go_16_goMux_choice_emitted;
  logic [1:0] go_16_goMux_choice_done;
  assign go_16_goMux_choice_1_d = {go_16_goMux_choice_d[2:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[0]))};
  assign go_16_goMux_choice_2_d = {go_16_goMux_choice_d[2:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[1]))};
  assign go_16_goMux_choice_done = (go_16_goMux_choice_emitted | ({go_16_goMux_choice_2_d[0],
                                                                   go_16_goMux_choice_1_d[0]} & {go_16_goMux_choice_2_r,
                                                                                                 go_16_goMux_choice_1_r}));
  assign go_16_goMux_choice_r = (& go_16_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_goMux_choice_emitted <= 2'd0;
    else
      go_16_goMux_choice_emitted <= (go_16_goMux_choice_r ? 2'd0 :
                                     go_16_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Pointer_QTree_Int) : (go_16_goMux_choice_1,C4) [(lizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet12_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [3:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet10_1_argbuf_d};
      2'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   contRet_0_1_1_argbuf_d};
      2'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet11_1_argbuf_d};
      2'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet12_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_1_d[0])};
  assign go_16_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet12_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (go_16_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (go_16_goMux_choice_2,C4) [(lizzieLet6_7QNone_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (sc_0_11_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (lizzieLet6_7QVal_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                      (lizzieLet6_7QError_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [3:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet6_7QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   sc_0_11_1_argbuf_d};
      2'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet6_7QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet6_7QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_2_d[0])};
  assign go_16_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_7QError_Int_1_argbuf_r,
          lizzieLet6_7QVal_Int_1_argbuf_r,
          sc_0_11_1_argbuf_r,
          lizzieLet6_7QNone_Int_1_argbuf_r} = (go_16_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C6) : (go_17_goMux_choice,C6) > [(go_17_goMux_choice_1,C6),
                                          (go_17_goMux_choice_2,C6)] */
  logic [1:0] go_17_goMux_choice_emitted;
  logic [1:0] go_17_goMux_choice_done;
  assign go_17_goMux_choice_1_d = {go_17_goMux_choice_d[3:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[0]))};
  assign go_17_goMux_choice_2_d = {go_17_goMux_choice_d[3:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[1]))};
  assign go_17_goMux_choice_done = (go_17_goMux_choice_emitted | ({go_17_goMux_choice_2_d[0],
                                                                   go_17_goMux_choice_1_d[0]} & {go_17_goMux_choice_2_r,
                                                                                                 go_17_goMux_choice_1_r}));
  assign go_17_goMux_choice_r = (& go_17_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_goMux_choice_emitted <= 2'd0;
    else
      go_17_goMux_choice_emitted <= (go_17_goMux_choice_r ? 2'd0 :
                                     go_17_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Int) : (go_17_goMux_choice_1,C6) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet10_1_5MQVal_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [5:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet10_1_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_1_d[0])};
  assign go_17_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet10_1_5MQVal_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_17_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTmain_mask_Int) : (go_17_goMux_choice_2,C6) [(lizzieLet10_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (sc_0_15_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet10_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf,Pointer_CTmain_mask_Int),
                                                              (lizzieLet10_1_4MQNode_4QError_Int_1_argbuf,Pointer_CTmain_mask_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTmain_mask_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [5:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet10_1_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd2,
                                                                   sc_0_15_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet10_1_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_d};
      3'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_2_d[0])};
  assign go_17_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_r,
          lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_r,
          lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_r,
          lizzieLet10_1_6MQVal_1_argbuf_r,
          sc_0_15_1_argbuf_r,
          lizzieLet10_1_6MQNone_1_argbuf_r} = (go_17_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                               6'd0);
  
  /* fork (Ty C5) : (go_18_goMux_choice,C5) > [(go_18_goMux_choice_1,C5),
                                          (go_18_goMux_choice_2,C5)] */
  logic [1:0] go_18_goMux_choice_emitted;
  logic [1:0] go_18_goMux_choice_done;
  assign go_18_goMux_choice_1_d = {go_18_goMux_choice_d[3:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[0]))};
  assign go_18_goMux_choice_2_d = {go_18_goMux_choice_d[3:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[1]))};
  assign go_18_goMux_choice_done = (go_18_goMux_choice_emitted | ({go_18_goMux_choice_2_d[0],
                                                                   go_18_goMux_choice_1_d[0]} & {go_18_goMux_choice_2_r,
                                                                                                 go_18_goMux_choice_1_r}));
  assign go_18_goMux_choice_r = (& go_18_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_goMux_choice_emitted <= 2'd0;
    else
      go_18_goMux_choice_emitted <= (go_18_goMux_choice_r ? 2'd0 :
                                     go_18_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_18_goMux_choice_1,C5) [(lizzieLet5_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet6_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet8_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_3_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_3_goMux_mux_mux;
  logic [4:0] srtarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet5_1_1_argbuf_d};
      3'd1:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_3_1_argbuf_d};
      3'd2:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet6_1_1_argbuf_d};
      3'd3:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet7_1_1_argbuf_d};
      3'd4:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet8_1_1_argbuf_d};
      default:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_3_goMux_mux_d = {srtarg_0_3_goMux_mux_mux[16:1],
                                   (srtarg_0_3_goMux_mux_mux[0] && go_18_goMux_choice_1_d[0])};
  assign go_18_goMux_choice_1_r = (srtarg_0_3_goMux_mux_d[0] && srtarg_0_3_goMux_mux_r);
  assign {lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          contRet_0_3_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = (go_18_goMux_choice_1_r ? srtarg_0_3_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Int_Int_Int) : (go_18_goMux_choice_2,C5) [(lizzieLet17_6QNone_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (sc_0_19_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (es_0_2_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (es_0_2_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int),
                                                                        (lizzieLet17_6QError_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int)] > (scfarg_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) */
  logic [16:0] scfarg_0_3_goMux_mux_mux;
  logic [4:0] scfarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet17_6QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd2,
                                                                   sc_0_19_1_argbuf_d};
      3'd2:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd4,
                                                                   es_0_2_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd8,
                                                                   es_0_2_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet17_6QError_Int_1_argbuf_d};
      default:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_3_goMux_mux_d = {scfarg_0_3_goMux_mux_mux[16:1],
                                   (scfarg_0_3_goMux_mux_mux[0] && go_18_goMux_choice_2_d[0])};
  assign go_18_goMux_choice_2_r = (scfarg_0_3_goMux_mux_d[0] && scfarg_0_3_goMux_mux_r);
  assign {lizzieLet17_6QError_Int_1_argbuf_r,
          es_0_2_2MyTrue_1_argbuf_r,
          es_0_2_2MyFalse_1_argbuf_r,
          sc_0_19_1_argbuf_r,
          lizzieLet17_6QNone_Int_1_argbuf_r} = (go_18_goMux_choice_2_r ? scfarg_0_3_goMux_mux_onehot :
                                                5'd0);
  
  /* buf (Ty MyDTInt_Int_Int) : (go_1Dcon_$fNumInt_$c*,MyDTInt_Int_Int) > (es_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$ctimes_bufchan_d ;
  logic \go_1Dcon_$fNumInt_$ctimes_bufchan_r ;
  assign \go_1Dcon_$fNumInt_$ctimes_r  = ((! \go_1Dcon_$fNumInt_$ctimes_bufchan_d [0]) || \go_1Dcon_$fNumInt_$ctimes_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$ctimes_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_$fNumInt_$ctimes_r )
        \go_1Dcon_$fNumInt_$ctimes_bufchan_d  <= \go_1Dcon_$fNumInt_$ctimes_d ;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$ctimes_bufchan_buf ;
  assign \go_1Dcon_$fNumInt_$ctimes_bufchan_r  = (! \go_1Dcon_$fNumInt_$ctimes_bufchan_buf [0]);
  assign es_4_1_argbuf_d = (\go_1Dcon_$fNumInt_$ctimes_bufchan_buf [0] ? \go_1Dcon_$fNumInt_$ctimes_bufchan_buf  :
                            \go_1Dcon_$fNumInt_$ctimes_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_1Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
    else
      if ((es_4_1_argbuf_r && \go_1Dcon_$fNumInt_$ctimes_bufchan_buf [0]))
        \go_1Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! \go_1Dcon_$fNumInt_$ctimes_bufchan_buf [0])))
        \go_1Dcon_$fNumInt_$ctimes_bufchan_buf  <= \go_1Dcon_$fNumInt_$ctimes_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_main1) : [(go_2,Go)] > (go_2Dcon_main1,MyDTInt_Bool) */
  assign go_2Dcon_main1_d = Dcon_main1_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_main1_r && go_2Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_2Dcon_main1,MyDTInt_Bool) > (es_3_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_2Dcon_main1_bufchan_d;
  logic go_2Dcon_main1_bufchan_r;
  assign go_2Dcon_main1_r = ((! go_2Dcon_main1_bufchan_d[0]) || go_2Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_main1_r) go_2Dcon_main1_bufchan_d <= go_2Dcon_main1_d;
  MyDTInt_Bool_t go_2Dcon_main1_bufchan_buf;
  assign go_2Dcon_main1_bufchan_r = (! go_2Dcon_main1_bufchan_buf[0]);
  assign es_3_1_argbuf_d = (go_2Dcon_main1_bufchan_buf[0] ? go_2Dcon_main1_bufchan_buf :
                            go_2Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_3_1_argbuf_r && go_2Dcon_main1_bufchan_buf[0]))
        go_2Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! go_2Dcon_main1_bufchan_buf[0])))
        go_2Dcon_main1_bufchan_buf <= go_2Dcon_main1_bufchan_d;
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_3_argbuf,Go),
                                                                                              (es_3_1_argbuf,MyDTInt_Bool),
                                                                                              (es_4_1_argbuf,MyDTInt_Int_Int),
                                                                                              (m2adm_1,Pointer_QTree_Int),
                                                                                              (m3adn_2,Pointer_QTree_Int)] > (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_3_argbuf_d[0],
                                                                                                                                                                                                         es_3_1_argbuf_d[0],
                                                                                                                                                                                                         es_4_1_argbuf_d[0],
                                                                                                                                                                                                         m2adm_1_d[0],
                                                                                                                                                                                                         m3adn_2_d[0]}), go_3_argbuf_d, es_3_1_argbuf_d, es_4_1_argbuf_d, m2adm_1_d, m3adn_2_d);
  assign {go_3_argbuf_r,
          es_3_1_argbuf_r,
          es_4_1_argbuf_r,
          m2adm_1_r,
          m3adn_2_r} = {5 {(kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_4,Go) > (go_4_argbuf,Go) */
  Go_t go_4_bufchan_d;
  logic go_4_bufchan_r;
  assign go_4_r = ((! go_4_bufchan_d[0]) || go_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_d <= 1'd0;
    else if (go_4_r) go_4_bufchan_d <= go_4_d;
  Go_t go_4_bufchan_buf;
  assign go_4_bufchan_r = (! go_4_bufchan_buf[0]);
  assign go_4_argbuf_d = (go_4_bufchan_buf[0] ? go_4_bufchan_buf :
                          go_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_buf <= 1'd0;
    else
      if ((go_4_argbuf_r && go_4_bufchan_buf[0]))
        go_4_bufchan_buf <= 1'd0;
      else if (((! go_4_argbuf_r) && (! go_4_bufchan_buf[0])))
        go_4_bufchan_buf <= go_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree,
      Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree) : [(go_4_argbuf,Go),
                                                             (es_1_1_argbuf,Pointer_QTree_Int),
                                                             (m1adl_0,Pointer_MaskQTree)] > (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree) */
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d = TupGo___Pointer_QTree_Int___Pointer_MaskQTree_dc((& {go_4_argbuf_d[0],
                                                                                                                               es_1_1_argbuf_d[0],
                                                                                                                               m1adl_0_d[0]}), go_4_argbuf_d, es_1_1_argbuf_d, m1adl_0_d);
  assign {go_4_argbuf_r,
          es_1_1_argbuf_r,
          m1adl_0_r} = {3 {(main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0])}};
  
  /* buf (Ty Go) : (go_5,Go) > (go_5_argbuf,Go) */
  Go_t go_5_bufchan_d;
  logic go_5_bufchan_r;
  assign go_5_r = ((! go_5_bufchan_d[0]) || go_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_d <= 1'd0;
    else if (go_5_r) go_5_bufchan_d <= go_5_d;
  Go_t go_5_bufchan_buf;
  assign go_5_bufchan_r = (! go_5_bufchan_buf[0]);
  assign go_5_argbuf_d = (go_5_bufchan_buf[0] ? go_5_bufchan_buf :
                          go_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_buf <= 1'd0;
    else
      if ((go_5_argbuf_r && go_5_bufchan_buf[0]))
        go_5_bufchan_buf <= 1'd0;
      else if (((! go_5_argbuf_r) && (! go_5_bufchan_buf[0])))
        go_5_bufchan_buf <= go_5_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_5_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_5_argbuf_d[0],
                                                                                     es_0_1_argbuf_d[0]}), go_5_argbuf_d, es_0_1_argbuf_d);
  assign {go_5_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  && \$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon L$wnnz_Intsbos) : [(go_6_1,Go)] > (go_6_1L$wnnz_Intsbos,CT$wnnz_Int) */
  assign go_6_1L$wnnz_Intsbos_d = L$wnnz_Intsbos_dc((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(go_6_1L$wnnz_Intsbos_r && go_6_1L$wnnz_Intsbos_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (go_6_1L$wnnz_Intsbos,CT$wnnz_Int) > (lizzieLet0_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_bufchan_d;
  logic go_6_1L$wnnz_Intsbos_bufchan_r;
  assign go_6_1L$wnnz_Intsbos_r = ((! go_6_1L$wnnz_Intsbos_bufchan_d[0]) || go_6_1L$wnnz_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wnnz_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_6_1L$wnnz_Intsbos_r)
        go_6_1L$wnnz_Intsbos_bufchan_d <= go_6_1L$wnnz_Intsbos_d;
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_bufchan_buf;
  assign go_6_1L$wnnz_Intsbos_bufchan_r = (! go_6_1L$wnnz_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_6_1L$wnnz_Intsbos_bufchan_buf[0] ? go_6_1L$wnnz_Intsbos_bufchan_buf :
                                  go_6_1L$wnnz_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_6_1L$wnnz_Intsbos_bufchan_buf[0]))
        go_6_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_6_1L$wnnz_Intsbos_bufchan_buf[0])))
        go_6_1L$wnnz_Intsbos_bufchan_buf <= go_6_1L$wnnz_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : [(go_6_2_argbuf,Go),
                                                               (wsxl_1_argbuf,Pointer_QTree_Int),
                                                               (lizzieLet16_1_argbuf,Pointer_CT$wnnz_Int)] > (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) */
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_dc((& {go_6_2_argbuf_d[0],
                                                                                                                                    wsxl_1_argbuf_d[0],
                                                                                                                                    lizzieLet16_1_argbuf_d[0]}), go_6_2_argbuf_d, wsxl_1_argbuf_d, lizzieLet16_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          wsxl_1_argbuf_r,
          lizzieLet16_1_argbuf_r} = {3 {(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0])}};
  
  /* fork (Ty C5) : (go_8_goMux_choice,C5) > [(go_8_goMux_choice_1,C5),
                                         (go_8_goMux_choice_2,C5)] */
  logic [1:0] go_8_goMux_choice_emitted;
  logic [1:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 2'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 2'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_8_goMux_choice_1,C5) [(call_$wnnz_Int_goMux2,Pointer_QTree_Int),
                                                       (q2acW_1_1_argbuf,Pointer_QTree_Int),
                                                       (q3acX_2_1_argbuf,Pointer_QTree_Int),
                                                       (q4acY_3_1_argbuf,Pointer_QTree_Int),
                                                       (q1acV_1_argbuf,Pointer_QTree_Int)] > (wsxl_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsxl_1_goMux_mux_mux;
  logic [4:0] wsxl_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux2_d};
      3'd1:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd2,
                                                           q2acW_1_1_argbuf_d};
      3'd2:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd4,
                                                           q3acX_2_1_argbuf_d};
      3'd3:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd8,
                                                           q4acY_3_1_argbuf_d};
      3'd4:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd16,
                                                           q1acV_1_argbuf_d};
      default:
        {wsxl_1_goMux_mux_onehot, wsxl_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsxl_1_goMux_mux_d = {wsxl_1_goMux_mux_mux[16:1],
                               (wsxl_1_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (wsxl_1_goMux_mux_d[0] && wsxl_1_goMux_mux_r);
  assign {q1acV_1_argbuf_r,
          q4acY_3_1_argbuf_r,
          q3acX_2_1_argbuf_r,
          q2acW_1_1_argbuf_r,
          call_$wnnz_Int_goMux2_r} = (go_8_goMux_choice_1_r ? wsxl_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz_Int) : (go_8_goMux_choice_2,C5) [(call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int),
                                                         (sca2_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca1_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca0_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca3_1_argbuf,Pointer_CT$wnnz_Int)] > (sc_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_Int_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_Int_goMux3_r} = (go_8_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                      5'd0);
  
  /* fork (Ty C5) : (go_9_goMux_choice,C5) > [(go_9_goMux_choice_1,C5),
                                         (go_9_goMux_choice_2,C5),
                                         (go_9_goMux_choice_3,C5),
                                         (go_9_goMux_choice_4,C5),
                                         (go_9_goMux_choice_5,C5)] */
  logic [4:0] go_9_goMux_choice_emitted;
  logic [4:0] go_9_goMux_choice_done;
  assign go_9_goMux_choice_1_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[0]))};
  assign go_9_goMux_choice_2_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[1]))};
  assign go_9_goMux_choice_3_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[2]))};
  assign go_9_goMux_choice_4_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[3]))};
  assign go_9_goMux_choice_5_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[4]))};
  assign go_9_goMux_choice_done = (go_9_goMux_choice_emitted | ({go_9_goMux_choice_5_d[0],
                                                                 go_9_goMux_choice_4_d[0],
                                                                 go_9_goMux_choice_3_d[0],
                                                                 go_9_goMux_choice_2_d[0],
                                                                 go_9_goMux_choice_1_d[0]} & {go_9_goMux_choice_5_r,
                                                                                              go_9_goMux_choice_4_r,
                                                                                              go_9_goMux_choice_3_r,
                                                                                              go_9_goMux_choice_2_r,
                                                                                              go_9_goMux_choice_1_r}));
  assign go_9_goMux_choice_r = (& go_9_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_goMux_choice_emitted <= 5'd0;
    else
      go_9_goMux_choice_emitted <= (go_9_goMux_choice_r ? 5'd0 :
                                    go_9_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_9_goMux_choice_1,C5) [(call_kron_kron_Int_Int_Int_goMux2,MyDTInt_Bool),
                                                  (isZacL_2_2_argbuf,MyDTInt_Bool),
                                                  (isZacL_3_2_argbuf,MyDTInt_Bool),
                                                  (isZacL_4_1_argbuf,MyDTInt_Bool),
                                                  (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (isZacL_goMux_mux,MyDTInt_Bool) */
  logic [0:0] isZacL_goMux_mux_mux;
  logic [4:0] isZacL_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_1_d[3:1])
      3'd0:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Int_Int_Int_goMux2_d};
      3'd1:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd2,
                                                           isZacL_2_2_argbuf_d};
      3'd2:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd4,
                                                           isZacL_3_2_argbuf_d};
      3'd3:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd8,
                                                           isZacL_4_1_argbuf_d};
      3'd4:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd16,
                                                           lizzieLet6_5QNode_Int_2_argbuf_d};
      default:
        {isZacL_goMux_mux_onehot, isZacL_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacL_goMux_mux_d = (isZacL_goMux_mux_mux[0] && go_9_goMux_choice_1_d[0]);
  assign go_9_goMux_choice_1_r = (isZacL_goMux_mux_d[0] && isZacL_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_2_argbuf_r,
          isZacL_4_1_argbuf_r,
          isZacL_3_2_argbuf_r,
          isZacL_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux2_r} = (go_9_goMux_choice_1_r ? isZacL_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_9_goMux_choice_2,C5) [(call_kron_kron_Int_Int_Int_goMux3,MyDTInt_Int_Int),
                                                     (gacM_2_2_argbuf,MyDTInt_Int_Int),
                                                     (gacM_3_2_argbuf,MyDTInt_Int_Int),
                                                     (gacM_4_1_argbuf,MyDTInt_Int_Int),
                                                     (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (gacM_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] gacM_goMux_mux_mux;
  logic [4:0] gacM_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_2_d[3:1])
      3'd0:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Int_Int_Int_goMux3_d};
      3'd1:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd2,
                                                       gacM_2_2_argbuf_d};
      3'd2:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd4,
                                                       gacM_3_2_argbuf_d};
      3'd3:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd8,
                                                       gacM_4_1_argbuf_d};
      3'd4:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd16,
                                                       lizzieLet6_3QNode_Int_2_argbuf_d};
      default:
        {gacM_goMux_mux_onehot, gacM_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacM_goMux_mux_d = (gacM_goMux_mux_mux[0] && go_9_goMux_choice_2_d[0]);
  assign go_9_goMux_choice_2_r = (gacM_goMux_mux_d[0] && gacM_goMux_mux_r);
  assign {lizzieLet6_3QNode_Int_2_argbuf_r,
          gacM_4_1_argbuf_r,
          gacM_3_2_argbuf_r,
          gacM_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux3_r} = (go_9_goMux_choice_2_r ? gacM_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_9_goMux_choice_3,C5) [(call_kron_kron_Int_Int_Int_goMux4,Pointer_QTree_Int),
                                                       (q3acS_1_1_argbuf,Pointer_QTree_Int),
                                                       (q2acR_2_1_argbuf,Pointer_QTree_Int),
                                                       (q1acQ_3_1_argbuf,Pointer_QTree_Int),
                                                       (q4acT_1_argbuf,Pointer_QTree_Int)] > (m1acN_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1acN_goMux_mux_mux;
  logic [4:0] m1acN_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_3_d[3:1])
      3'd0:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Int_Int_Int_goMux4_d};
      3'd1:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd2,
                                                         q3acS_1_1_argbuf_d};
      3'd2:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd4,
                                                         q2acR_2_1_argbuf_d};
      3'd3:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd8,
                                                         q1acQ_3_1_argbuf_d};
      3'd4:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd16,
                                                         q4acT_1_argbuf_d};
      default:
        {m1acN_goMux_mux_onehot, m1acN_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1acN_goMux_mux_d = {m1acN_goMux_mux_mux[16:1],
                              (m1acN_goMux_mux_mux[0] && go_9_goMux_choice_3_d[0])};
  assign go_9_goMux_choice_3_r = (m1acN_goMux_mux_d[0] && m1acN_goMux_mux_r);
  assign {q4acT_1_argbuf_r,
          q1acQ_3_1_argbuf_r,
          q2acR_2_1_argbuf_r,
          q3acS_1_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux4_r} = (go_9_goMux_choice_3_r ? m1acN_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_9_goMux_choice_4,C5) [(call_kron_kron_Int_Int_Int_goMux5,Pointer_QTree_Int),
                                                       (m2acO_2_2_argbuf,Pointer_QTree_Int),
                                                       (m2acO_3_2_argbuf,Pointer_QTree_Int),
                                                       (m2acO_4_1_argbuf,Pointer_QTree_Int),
                                                       (lizzieLet6_6QNode_Int_2_argbuf,Pointer_QTree_Int)] > (m2acO_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2acO_goMux_mux_mux;
  logic [4:0] m2acO_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_4_d[3:1])
      3'd0:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Int_Int_Int_goMux5_d};
      3'd1:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd2,
                                                         m2acO_2_2_argbuf_d};
      3'd2:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd4,
                                                         m2acO_3_2_argbuf_d};
      3'd3:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd8,
                                                         m2acO_4_1_argbuf_d};
      3'd4:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd16,
                                                         lizzieLet6_6QNode_Int_2_argbuf_d};
      default:
        {m2acO_goMux_mux_onehot, m2acO_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2acO_goMux_mux_d = {m2acO_goMux_mux_mux[16:1],
                              (m2acO_goMux_mux_mux[0] && go_9_goMux_choice_4_d[0])};
  assign go_9_goMux_choice_4_r = (m2acO_goMux_mux_d[0] && m2acO_goMux_mux_r);
  assign {lizzieLet6_6QNode_Int_2_argbuf_r,
          m2acO_4_1_argbuf_r,
          m2acO_3_2_argbuf_r,
          m2acO_2_2_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux5_r} = (go_9_goMux_choice_4_r ? m2acO_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTkron_kron_Int_Int_Int) : (go_9_goMux_choice_5,C5) [(call_kron_kron_Int_Int_Int_goMux6,Pointer_CTkron_kron_Int_Int_Int),
                                                                     (sca2_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                     (sca1_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                     (sca0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int),
                                                                     (sca3_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int)] > (sc_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Int_Int_Int_goMux6_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_9_goMux_choice_5_d[0])};
  assign go_9_goMux_choice_5_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_kron_kron_Int_Int_Int_goMux6_r} = (go_9_goMux_choice_5_r ? sc_0_1_goMux_mux_onehot :
                                                  5'd0);
  
  /* buf (Ty MyDTInt_Bool) : (isZacC_2_2,MyDTInt_Bool) > (isZacC_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacC_2_2_bufchan_d;
  logic isZacC_2_2_bufchan_r;
  assign isZacC_2_2_r = ((! isZacC_2_2_bufchan_d[0]) || isZacC_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_2_2_bufchan_d <= 1'd0;
    else if (isZacC_2_2_r) isZacC_2_2_bufchan_d <= isZacC_2_2_d;
  MyDTInt_Bool_t isZacC_2_2_bufchan_buf;
  assign isZacC_2_2_bufchan_r = (! isZacC_2_2_bufchan_buf[0]);
  assign isZacC_2_2_argbuf_d = (isZacC_2_2_bufchan_buf[0] ? isZacC_2_2_bufchan_buf :
                                isZacC_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacC_2_2_argbuf_r && isZacC_2_2_bufchan_buf[0]))
        isZacC_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacC_2_2_argbuf_r) && (! isZacC_2_2_bufchan_buf[0])))
        isZacC_2_2_bufchan_buf <= isZacC_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacC_2_destruct,MyDTInt_Bool) > [(isZacC_2_1,MyDTInt_Bool),
                                                             (isZacC_2_2,MyDTInt_Bool)] */
  logic [1:0] isZacC_2_destruct_emitted;
  logic [1:0] isZacC_2_destruct_done;
  assign isZacC_2_1_d = (isZacC_2_destruct_d[0] && (! isZacC_2_destruct_emitted[0]));
  assign isZacC_2_2_d = (isZacC_2_destruct_d[0] && (! isZacC_2_destruct_emitted[1]));
  assign isZacC_2_destruct_done = (isZacC_2_destruct_emitted | ({isZacC_2_2_d[0],
                                                                 isZacC_2_1_d[0]} & {isZacC_2_2_r,
                                                                                     isZacC_2_1_r}));
  assign isZacC_2_destruct_r = (& isZacC_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_2_destruct_emitted <= 2'd0;
    else
      isZacC_2_destruct_emitted <= (isZacC_2_destruct_r ? 2'd0 :
                                    isZacC_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacC_3_2,MyDTInt_Bool) > (isZacC_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacC_3_2_bufchan_d;
  logic isZacC_3_2_bufchan_r;
  assign isZacC_3_2_r = ((! isZacC_3_2_bufchan_d[0]) || isZacC_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_3_2_bufchan_d <= 1'd0;
    else if (isZacC_3_2_r) isZacC_3_2_bufchan_d <= isZacC_3_2_d;
  MyDTInt_Bool_t isZacC_3_2_bufchan_buf;
  assign isZacC_3_2_bufchan_r = (! isZacC_3_2_bufchan_buf[0]);
  assign isZacC_3_2_argbuf_d = (isZacC_3_2_bufchan_buf[0] ? isZacC_3_2_bufchan_buf :
                                isZacC_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacC_3_2_argbuf_r && isZacC_3_2_bufchan_buf[0]))
        isZacC_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacC_3_2_argbuf_r) && (! isZacC_3_2_bufchan_buf[0])))
        isZacC_3_2_bufchan_buf <= isZacC_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacC_3_destruct,MyDTInt_Bool) > [(isZacC_3_1,MyDTInt_Bool),
                                                             (isZacC_3_2,MyDTInt_Bool)] */
  logic [1:0] isZacC_3_destruct_emitted;
  logic [1:0] isZacC_3_destruct_done;
  assign isZacC_3_1_d = (isZacC_3_destruct_d[0] && (! isZacC_3_destruct_emitted[0]));
  assign isZacC_3_2_d = (isZacC_3_destruct_d[0] && (! isZacC_3_destruct_emitted[1]));
  assign isZacC_3_destruct_done = (isZacC_3_destruct_emitted | ({isZacC_3_2_d[0],
                                                                 isZacC_3_1_d[0]} & {isZacC_3_2_r,
                                                                                     isZacC_3_1_r}));
  assign isZacC_3_destruct_r = (& isZacC_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_3_destruct_emitted <= 2'd0;
    else
      isZacC_3_destruct_emitted <= (isZacC_3_destruct_r ? 2'd0 :
                                    isZacC_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacC_4_destruct,MyDTInt_Bool) > (isZacC_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacC_4_destruct_bufchan_d;
  logic isZacC_4_destruct_bufchan_r;
  assign isZacC_4_destruct_r = ((! isZacC_4_destruct_bufchan_d[0]) || isZacC_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacC_4_destruct_r)
        isZacC_4_destruct_bufchan_d <= isZacC_4_destruct_d;
  MyDTInt_Bool_t isZacC_4_destruct_bufchan_buf;
  assign isZacC_4_destruct_bufchan_r = (! isZacC_4_destruct_bufchan_buf[0]);
  assign isZacC_4_1_argbuf_d = (isZacC_4_destruct_bufchan_buf[0] ? isZacC_4_destruct_bufchan_buf :
                                isZacC_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacC_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacC_4_1_argbuf_r && isZacC_4_destruct_bufchan_buf[0]))
        isZacC_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacC_4_1_argbuf_r) && (! isZacC_4_destruct_bufchan_buf[0])))
        isZacC_4_destruct_bufchan_buf <= isZacC_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_2_2,MyDTInt_Bool) > (isZacL_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_2_2_bufchan_d;
  logic isZacL_2_2_bufchan_r;
  assign isZacL_2_2_r = ((! isZacL_2_2_bufchan_d[0]) || isZacL_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_2_bufchan_d <= 1'd0;
    else if (isZacL_2_2_r) isZacL_2_2_bufchan_d <= isZacL_2_2_d;
  MyDTInt_Bool_t isZacL_2_2_bufchan_buf;
  assign isZacL_2_2_bufchan_r = (! isZacL_2_2_bufchan_buf[0]);
  assign isZacL_2_2_argbuf_d = (isZacL_2_2_bufchan_buf[0] ? isZacL_2_2_bufchan_buf :
                                isZacL_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacL_2_2_argbuf_r && isZacL_2_2_bufchan_buf[0]))
        isZacL_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacL_2_2_argbuf_r) && (! isZacL_2_2_bufchan_buf[0])))
        isZacL_2_2_bufchan_buf <= isZacL_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacL_2_destruct,MyDTInt_Bool) > [(isZacL_2_1,MyDTInt_Bool),
                                                             (isZacL_2_2,MyDTInt_Bool)] */
  logic [1:0] isZacL_2_destruct_emitted;
  logic [1:0] isZacL_2_destruct_done;
  assign isZacL_2_1_d = (isZacL_2_destruct_d[0] && (! isZacL_2_destruct_emitted[0]));
  assign isZacL_2_2_d = (isZacL_2_destruct_d[0] && (! isZacL_2_destruct_emitted[1]));
  assign isZacL_2_destruct_done = (isZacL_2_destruct_emitted | ({isZacL_2_2_d[0],
                                                                 isZacL_2_1_d[0]} & {isZacL_2_2_r,
                                                                                     isZacL_2_1_r}));
  assign isZacL_2_destruct_r = (& isZacL_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_2_destruct_emitted <= 2'd0;
    else
      isZacL_2_destruct_emitted <= (isZacL_2_destruct_r ? 2'd0 :
                                    isZacL_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_3_2,MyDTInt_Bool) > (isZacL_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_3_2_bufchan_d;
  logic isZacL_3_2_bufchan_r;
  assign isZacL_3_2_r = ((! isZacL_3_2_bufchan_d[0]) || isZacL_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_2_bufchan_d <= 1'd0;
    else if (isZacL_3_2_r) isZacL_3_2_bufchan_d <= isZacL_3_2_d;
  MyDTInt_Bool_t isZacL_3_2_bufchan_buf;
  assign isZacL_3_2_bufchan_r = (! isZacL_3_2_bufchan_buf[0]);
  assign isZacL_3_2_argbuf_d = (isZacL_3_2_bufchan_buf[0] ? isZacL_3_2_bufchan_buf :
                                isZacL_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacL_3_2_argbuf_r && isZacL_3_2_bufchan_buf[0]))
        isZacL_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacL_3_2_argbuf_r) && (! isZacL_3_2_bufchan_buf[0])))
        isZacL_3_2_bufchan_buf <= isZacL_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (isZacL_3_destruct,MyDTInt_Bool) > [(isZacL_3_1,MyDTInt_Bool),
                                                             (isZacL_3_2,MyDTInt_Bool)] */
  logic [1:0] isZacL_3_destruct_emitted;
  logic [1:0] isZacL_3_destruct_done;
  assign isZacL_3_1_d = (isZacL_3_destruct_d[0] && (! isZacL_3_destruct_emitted[0]));
  assign isZacL_3_2_d = (isZacL_3_destruct_d[0] && (! isZacL_3_destruct_emitted[1]));
  assign isZacL_3_destruct_done = (isZacL_3_destruct_emitted | ({isZacL_3_2_d[0],
                                                                 isZacL_3_1_d[0]} & {isZacL_3_2_r,
                                                                                     isZacL_3_1_r}));
  assign isZacL_3_destruct_r = (& isZacL_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_3_destruct_emitted <= 2'd0;
    else
      isZacL_3_destruct_emitted <= (isZacL_3_destruct_r ? 2'd0 :
                                    isZacL_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (isZacL_4_destruct,MyDTInt_Bool) > (isZacL_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t isZacL_4_destruct_bufchan_d;
  logic isZacL_4_destruct_bufchan_r;
  assign isZacL_4_destruct_r = ((! isZacL_4_destruct_bufchan_d[0]) || isZacL_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacL_4_destruct_r)
        isZacL_4_destruct_bufchan_d <= isZacL_4_destruct_d;
  MyDTInt_Bool_t isZacL_4_destruct_bufchan_buf;
  assign isZacL_4_destruct_bufchan_r = (! isZacL_4_destruct_bufchan_buf[0]);
  assign isZacL_4_1_argbuf_d = (isZacL_4_destruct_bufchan_buf[0] ? isZacL_4_destruct_bufchan_buf :
                                isZacL_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacL_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacL_4_1_argbuf_r && isZacL_4_destruct_bufchan_buf[0]))
        isZacL_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacL_4_1_argbuf_r) && (! isZacL_4_destruct_bufchan_buf[0])))
        isZacL_4_destruct_bufchan_buf <= isZacL_4_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) > [(kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12,Go),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                           (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1,Pointer_QTree_Int)] */
  logic [4:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted;
  logic [4:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[0]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[1]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[2]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_d = {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[16:1],
                                                                                                                         (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[3]))};
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_d = {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[32:17],
                                                                                                                         (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[4]))};
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted | ({kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_d[0],
                                                                                                                                                                                                                                         kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_d[0]} & {kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_r,
                                                                                                                                                                                                                                                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_r}));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r = (& kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= 5'd0;
    else
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r ? 5'd0 :
                                                                                                                        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1,MyDTInt_Int_Int) > (gacM_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_d;
  MyDTInt_Int_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf[0]);
  assign gacM_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf :
                              kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf <= 1'd0;
    else
      if ((gacM_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf <= 1'd0;
      else if (((! gacM_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntgacM_1_bufchan_d;
  
  /* fork (Ty Go) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12,Go) > [(go_12_1,Go),
                                                                                                                                (go_12_2,Go)] */
  logic [1:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted;
  logic [1:0] kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_done;
  assign go_12_1_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted[0]));
  assign go_12_2_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_d[0] && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted[1]));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_done = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted | ({go_12_2_d[0],
                                                                                                                                                                                                                                               go_12_1_d[0]} & {go_12_2_r,
                                                                                                                                                                                                                                                                go_12_1_r}));
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_r = (& kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted <= 2'd0;
    else
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_emitted <= (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_r ? 2'd0 :
                                                                                                                           kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_12_done);
  
  /* buf (Ty MyDTInt_Bool) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1,MyDTInt_Bool) > (isZacL_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_d;
  MyDTInt_Bool_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf[0]);
  assign isZacL_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf :
                                kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf <= 1'd0;
    else
      if ((isZacL_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf <= 1'd0;
      else if (((! isZacL_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntisZacL_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1,Pointer_QTree_Int) > (m1acN_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d <= {16'd0,
                                                                                                                               1'd0};
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf[0]);
  assign m1acN_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf :
                               kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((m1acN_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! m1acN_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm1acN_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1,Pointer_QTree_Int) > (m2acO_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d;
  logic kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_r;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_r = ((! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d[0]) || kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d <= {16'd0,
                                                                                                                               1'd0};
    else
      if (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_r)
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf;
  assign kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_r = (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf[0]);
  assign m2acO_1_1_argbuf_d = (kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf[0] ? kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf :
                               kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((m2acO_1_1_argbuf_r && kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf[0]))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! m2acO_1_1_argbuf_r) && (! kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf[0])))
        kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_buf <= kron_kron_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intm2acO_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (kron_kron_Int_Int_Int_resbuf,Pointer_QTree_Int) > (es_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_bufchan_d;
  logic kron_kron_Int_Int_Int_resbuf_bufchan_r;
  assign kron_kron_Int_Int_Int_resbuf_r = ((! kron_kron_Int_Int_Int_resbuf_bufchan_d[0]) || kron_kron_Int_Int_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (kron_kron_Int_Int_Int_resbuf_r)
        kron_kron_Int_Int_Int_resbuf_bufchan_d <= kron_kron_Int_Int_Int_resbuf_d;
  Pointer_QTree_Int_t kron_kron_Int_Int_Int_resbuf_bufchan_buf;
  assign kron_kron_Int_Int_Int_resbuf_bufchan_r = (! kron_kron_Int_Int_Int_resbuf_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (kron_kron_Int_Int_Int_resbuf_bufchan_buf[0] ? kron_kron_Int_Int_Int_resbuf_bufchan_buf :
                            kron_kron_Int_Int_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && kron_kron_Int_Int_Int_resbuf_bufchan_buf[0]))
        kron_kron_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! kron_kron_Int_Int_Int_resbuf_bufchan_buf[0])))
        kron_kron_Int_Int_Int_resbuf_bufchan_buf <= kron_kron_Int_Int_Int_resbuf_bufchan_d;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet10_1_1MQNode,MaskQTree) > [(q1acm_destruct,Pointer_MaskQTree),
                                                              (q2acn_destruct,Pointer_MaskQTree),
                                                              (q3aco_destruct,Pointer_MaskQTree),
                                                              (q4acp_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet10_1_1MQNode_emitted;
  logic [3:0] lizzieLet10_1_1MQNode_done;
  assign q1acm_destruct_d = {lizzieLet10_1_1MQNode_d[18:3],
                             (lizzieLet10_1_1MQNode_d[0] && (! lizzieLet10_1_1MQNode_emitted[0]))};
  assign q2acn_destruct_d = {lizzieLet10_1_1MQNode_d[34:19],
                             (lizzieLet10_1_1MQNode_d[0] && (! lizzieLet10_1_1MQNode_emitted[1]))};
  assign q3aco_destruct_d = {lizzieLet10_1_1MQNode_d[50:35],
                             (lizzieLet10_1_1MQNode_d[0] && (! lizzieLet10_1_1MQNode_emitted[2]))};
  assign q4acp_destruct_d = {lizzieLet10_1_1MQNode_d[66:51],
                             (lizzieLet10_1_1MQNode_d[0] && (! lizzieLet10_1_1MQNode_emitted[3]))};
  assign lizzieLet10_1_1MQNode_done = (lizzieLet10_1_1MQNode_emitted | ({q4acp_destruct_d[0],
                                                                         q3aco_destruct_d[0],
                                                                         q2acn_destruct_d[0],
                                                                         q1acm_destruct_d[0]} & {q4acp_destruct_r,
                                                                                                 q3aco_destruct_r,
                                                                                                 q2acn_destruct_r,
                                                                                                 q1acm_destruct_r}));
  assign lizzieLet10_1_1MQNode_r = (& lizzieLet10_1_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1MQNode_emitted <= 4'd0;
    else
      lizzieLet10_1_1MQNode_emitted <= (lizzieLet10_1_1MQNode_r ? 4'd0 :
                                        lizzieLet10_1_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet10_1_2,MaskQTree) (lizzieLet10_1_1,MaskQTree) > [(_47,MaskQTree),
                                                                                  (_46,MaskQTree),
                                                                                  (lizzieLet10_1_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet10_1_1_onehotd;
  always_comb
    if ((lizzieLet10_1_2_d[0] && lizzieLet10_1_1_d[0]))
      unique case (lizzieLet10_1_2_d[2:1])
        2'd0: lizzieLet10_1_1_onehotd = 3'd1;
        2'd1: lizzieLet10_1_1_onehotd = 3'd2;
        2'd2: lizzieLet10_1_1_onehotd = 3'd4;
        default: lizzieLet10_1_1_onehotd = 3'd0;
      endcase
    else lizzieLet10_1_1_onehotd = 3'd0;
  assign _47_d = {lizzieLet10_1_1_d[66:1],
                  lizzieLet10_1_1_onehotd[0]};
  assign _46_d = {lizzieLet10_1_1_d[66:1],
                  lizzieLet10_1_1_onehotd[1]};
  assign lizzieLet10_1_1MQNode_d = {lizzieLet10_1_1_d[66:1],
                                    lizzieLet10_1_1_onehotd[2]};
  assign lizzieLet10_1_1_r = (| (lizzieLet10_1_1_onehotd & {lizzieLet10_1_1MQNode_r,
                                                            _46_r,
                                                            _47_r}));
  assign lizzieLet10_1_2_r = lizzieLet10_1_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet10_1_3,MaskQTree) (go_10_goMux_data,Go) > [(lizzieLet10_1_3MQNone,Go),
                                                                     (lizzieLet10_1_3MQVal,Go),
                                                                     (lizzieLet10_1_3MQNode,Go)] */
  logic [2:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet10_1_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet10_1_3_d[2:1])
        2'd0: go_10_goMux_data_onehotd = 3'd1;
        2'd1: go_10_goMux_data_onehotd = 3'd2;
        2'd2: go_10_goMux_data_onehotd = 3'd4;
        default: go_10_goMux_data_onehotd = 3'd0;
      endcase
    else go_10_goMux_data_onehotd = 3'd0;
  assign lizzieLet10_1_3MQNone_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet10_1_3MQVal_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet10_1_3MQNode_d = go_10_goMux_data_onehotd[2];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet10_1_3MQNode_r,
                                                              lizzieLet10_1_3MQVal_r,
                                                              lizzieLet10_1_3MQNone_r}));
  assign lizzieLet10_1_3_r = go_10_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet10_1_3MQNone,Go) > [(lizzieLet10_1_3MQNone_1,Go),
                                             (lizzieLet10_1_3MQNone_2,Go)] */
  logic [1:0] lizzieLet10_1_3MQNone_emitted;
  logic [1:0] lizzieLet10_1_3MQNone_done;
  assign lizzieLet10_1_3MQNone_1_d = (lizzieLet10_1_3MQNone_d[0] && (! lizzieLet10_1_3MQNone_emitted[0]));
  assign lizzieLet10_1_3MQNone_2_d = (lizzieLet10_1_3MQNone_d[0] && (! lizzieLet10_1_3MQNone_emitted[1]));
  assign lizzieLet10_1_3MQNone_done = (lizzieLet10_1_3MQNone_emitted | ({lizzieLet10_1_3MQNone_2_d[0],
                                                                         lizzieLet10_1_3MQNone_1_d[0]} & {lizzieLet10_1_3MQNone_2_r,
                                                                                                          lizzieLet10_1_3MQNone_1_r}));
  assign lizzieLet10_1_3MQNone_r = (& lizzieLet10_1_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQNone_emitted <= 2'd0;
    else
      lizzieLet10_1_3MQNone_emitted <= (lizzieLet10_1_3MQNone_r ? 2'd0 :
                                        lizzieLet10_1_3MQNone_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet10_1_3MQNone_1,Go)] > (lizzieLet10_1_3MQNone_1QNone_Int,QTree_Int) */
  assign lizzieLet10_1_3MQNone_1QNone_Int_d = QNone_Int_dc((& {lizzieLet10_1_3MQNone_1_d[0]}), lizzieLet10_1_3MQNone_1_d);
  assign {lizzieLet10_1_3MQNone_1_r} = {1 {(lizzieLet10_1_3MQNone_1QNone_Int_r && lizzieLet10_1_3MQNone_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_1_3MQNone_1QNone_Int,QTree_Int) > (lizzieLet11_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d;
  logic lizzieLet10_1_3MQNone_1QNone_Int_bufchan_r;
  assign lizzieLet10_1_3MQNone_1QNone_Int_r = ((! lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d[0]) || lizzieLet10_1_3MQNone_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet10_1_3MQNone_1QNone_Int_r)
        lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d <= lizzieLet10_1_3MQNone_1QNone_Int_d;
  QTree_Int_t lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf;
  assign lizzieLet10_1_3MQNone_1QNone_Int_bufchan_r = (! lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf[0] ? lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf :
                                     lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf[0]))
        lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf[0])))
        lizzieLet10_1_3MQNone_1QNone_Int_bufchan_buf <= lizzieLet10_1_3MQNone_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_1_3MQNone_2,Go) > (lizzieLet10_1_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet10_1_3MQNone_2_bufchan_d;
  logic lizzieLet10_1_3MQNone_2_bufchan_r;
  assign lizzieLet10_1_3MQNone_2_r = ((! lizzieLet10_1_3MQNone_2_bufchan_d[0]) || lizzieLet10_1_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_3MQNone_2_r)
        lizzieLet10_1_3MQNone_2_bufchan_d <= lizzieLet10_1_3MQNone_2_d;
  Go_t lizzieLet10_1_3MQNone_2_bufchan_buf;
  assign lizzieLet10_1_3MQNone_2_bufchan_r = (! lizzieLet10_1_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet10_1_3MQNone_2_argbuf_d = (lizzieLet10_1_3MQNone_2_bufchan_buf[0] ? lizzieLet10_1_3MQNone_2_bufchan_buf :
                                             lizzieLet10_1_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_3MQNone_2_argbuf_r && lizzieLet10_1_3MQNone_2_bufchan_buf[0]))
        lizzieLet10_1_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_3MQNone_2_argbuf_r) && (! lizzieLet10_1_3MQNone_2_bufchan_buf[0])))
        lizzieLet10_1_3MQNone_2_bufchan_buf <= lizzieLet10_1_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet10_1_3MQNone_2_argbuf,Go),
                           (lizzieLet35_3Lcall_main_mask_Int0_1_argbuf,Go),
                           (lizzieLet10_1_3MQVal_1_argbuf,Go),
                           (lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf,Go),
                           (lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf,Go),
                           (lizzieLet10_1_4MQNode_3QError_Int_2_argbuf,Go)] > (go_17_goMux_choice,C6) (go_17_goMux_data,Go) */
  logic [5:0] lizzieLet10_1_3MQNone_2_argbuf_select_d;
  assign lizzieLet10_1_3MQNone_2_argbuf_select_d = ((| lizzieLet10_1_3MQNone_2_argbuf_select_q) ? lizzieLet10_1_3MQNone_2_argbuf_select_q :
                                                    (lizzieLet10_1_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                     (lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_d[0] ? 6'd2 :
                                                      (lizzieLet10_1_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                       (lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_d[0] ? 6'd8 :
                                                        (lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_d[0] ? 6'd16 :
                                                         (lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_d[0] ? 6'd32 :
                                                          6'd0)))))));
  logic [5:0] lizzieLet10_1_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet10_1_3MQNone_2_argbuf_select_q <= (lizzieLet10_1_3MQNone_2_argbuf_done ? 6'd0 :
                                                  lizzieLet10_1_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet10_1_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_3MQNone_2_argbuf_emit_q <= (lizzieLet10_1_3MQNone_2_argbuf_done ? 2'd0 :
                                                lizzieLet10_1_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_3MQNone_2_argbuf_emit_d;
  assign lizzieLet10_1_3MQNone_2_argbuf_emit_d = (lizzieLet10_1_3MQNone_2_argbuf_emit_q | ({go_17_goMux_choice_d[0],
                                                                                            go_17_goMux_data_d[0]} & {go_17_goMux_choice_r,
                                                                                                                      go_17_goMux_data_r}));
  logic lizzieLet10_1_3MQNone_2_argbuf_done;
  assign lizzieLet10_1_3MQNone_2_argbuf_done = (& lizzieLet10_1_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_r,
          lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_r,
          lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_r,
          lizzieLet10_1_3MQVal_1_argbuf_r,
          lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_r,
          lizzieLet10_1_3MQNone_2_argbuf_r} = (lizzieLet10_1_3MQNone_2_argbuf_done ? lizzieLet10_1_3MQNone_2_argbuf_select_d :
                                               6'd0);
  assign go_17_goMux_data_d = ((lizzieLet10_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet10_1_3MQNone_2_argbuf_d :
                               ((lizzieLet10_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_d :
                                ((lizzieLet10_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet10_1_3MQVal_1_argbuf_d :
                                 ((lizzieLet10_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_d :
                                  ((lizzieLet10_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_d :
                                   ((lizzieLet10_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_d :
                                    1'd0))))));
  assign go_17_goMux_choice_d = ((lizzieLet10_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet10_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet10_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet10_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet10_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet10_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet10_1_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet10_1_3MQVal,Go) > (lizzieLet10_1_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet10_1_3MQVal_bufchan_d;
  logic lizzieLet10_1_3MQVal_bufchan_r;
  assign lizzieLet10_1_3MQVal_r = ((! lizzieLet10_1_3MQVal_bufchan_d[0]) || lizzieLet10_1_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_3MQVal_r)
        lizzieLet10_1_3MQVal_bufchan_d <= lizzieLet10_1_3MQVal_d;
  Go_t lizzieLet10_1_3MQVal_bufchan_buf;
  assign lizzieLet10_1_3MQVal_bufchan_r = (! lizzieLet10_1_3MQVal_bufchan_buf[0]);
  assign lizzieLet10_1_3MQVal_1_argbuf_d = (lizzieLet10_1_3MQVal_bufchan_buf[0] ? lizzieLet10_1_3MQVal_bufchan_buf :
                                            lizzieLet10_1_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_3MQVal_1_argbuf_r && lizzieLet10_1_3MQVal_bufchan_buf[0]))
        lizzieLet10_1_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_3MQVal_1_argbuf_r) && (! lizzieLet10_1_3MQVal_bufchan_buf[0])))
        lizzieLet10_1_3MQVal_bufchan_buf <= lizzieLet10_1_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Int) : (lizzieLet10_1_4,MaskQTree) (readPointer_QTree_Intmack_1_argbuf_rwb,QTree_Int) > [(_45,QTree_Int),
                                                                                                         (_44,QTree_Int),
                                                                                                         (lizzieLet10_1_4MQNode,QTree_Int)] */
  logic [2:0] readPointer_QTree_Intmack_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet10_1_4_d[0] && readPointer_QTree_Intmack_1_argbuf_rwb_d[0]))
      unique case (lizzieLet10_1_4_d[2:1])
        2'd0: readPointer_QTree_Intmack_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Intmack_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Intmack_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Intmack_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Intmack_1_argbuf_rwb_onehotd = 3'd0;
  assign _45_d = {readPointer_QTree_Intmack_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intmack_1_argbuf_rwb_onehotd[0]};
  assign _44_d = {readPointer_QTree_Intmack_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intmack_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet10_1_4MQNode_d = {readPointer_QTree_Intmack_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intmack_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Intmack_1_argbuf_rwb_r = (| (readPointer_QTree_Intmack_1_argbuf_rwb_onehotd & {lizzieLet10_1_4MQNode_r,
                                                                                                          _44_r,
                                                                                                          _45_r}));
  assign lizzieLet10_1_4_r = readPointer_QTree_Intmack_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet10_1_4MQNode,QTree_Int) > [(lizzieLet10_1_4MQNode_1,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_2,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_3,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_4,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_5,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_6,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_7,QTree_Int),
                                                           (lizzieLet10_1_4MQNode_8,QTree_Int)] */
  logic [7:0] lizzieLet10_1_4MQNode_emitted;
  logic [7:0] lizzieLet10_1_4MQNode_done;
  assign lizzieLet10_1_4MQNode_1_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[0]))};
  assign lizzieLet10_1_4MQNode_2_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[1]))};
  assign lizzieLet10_1_4MQNode_3_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[2]))};
  assign lizzieLet10_1_4MQNode_4_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[3]))};
  assign lizzieLet10_1_4MQNode_5_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[4]))};
  assign lizzieLet10_1_4MQNode_6_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[5]))};
  assign lizzieLet10_1_4MQNode_7_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[6]))};
  assign lizzieLet10_1_4MQNode_8_d = {lizzieLet10_1_4MQNode_d[66:1],
                                      (lizzieLet10_1_4MQNode_d[0] && (! lizzieLet10_1_4MQNode_emitted[7]))};
  assign lizzieLet10_1_4MQNode_done = (lizzieLet10_1_4MQNode_emitted | ({lizzieLet10_1_4MQNode_8_d[0],
                                                                         lizzieLet10_1_4MQNode_7_d[0],
                                                                         lizzieLet10_1_4MQNode_6_d[0],
                                                                         lizzieLet10_1_4MQNode_5_d[0],
                                                                         lizzieLet10_1_4MQNode_4_d[0],
                                                                         lizzieLet10_1_4MQNode_3_d[0],
                                                                         lizzieLet10_1_4MQNode_2_d[0],
                                                                         lizzieLet10_1_4MQNode_1_d[0]} & {lizzieLet10_1_4MQNode_8_r,
                                                                                                          lizzieLet10_1_4MQNode_7_r,
                                                                                                          lizzieLet10_1_4MQNode_6_r,
                                                                                                          lizzieLet10_1_4MQNode_5_r,
                                                                                                          lizzieLet10_1_4MQNode_4_r,
                                                                                                          lizzieLet10_1_4MQNode_3_r,
                                                                                                          lizzieLet10_1_4MQNode_2_r,
                                                                                                          lizzieLet10_1_4MQNode_1_r}));
  assign lizzieLet10_1_4MQNode_r = (& lizzieLet10_1_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_4MQNode_emitted <= 8'd0;
    else
      lizzieLet10_1_4MQNode_emitted <= (lizzieLet10_1_4MQNode_r ? 8'd0 :
                                        lizzieLet10_1_4MQNode_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet10_1_4MQNode_1QNode_Int,QTree_Int) > [(t1acr_destruct,Pointer_QTree_Int),
                                                                            (t2acs_destruct,Pointer_QTree_Int),
                                                                            (t3act_destruct,Pointer_QTree_Int),
                                                                            (t4acu_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet10_1_4MQNode_1QNode_Int_emitted;
  logic [3:0] lizzieLet10_1_4MQNode_1QNode_Int_done;
  assign t1acr_destruct_d = {lizzieLet10_1_4MQNode_1QNode_Int_d[18:3],
                             (lizzieLet10_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet10_1_4MQNode_1QNode_Int_emitted[0]))};
  assign t2acs_destruct_d = {lizzieLet10_1_4MQNode_1QNode_Int_d[34:19],
                             (lizzieLet10_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet10_1_4MQNode_1QNode_Int_emitted[1]))};
  assign t3act_destruct_d = {lizzieLet10_1_4MQNode_1QNode_Int_d[50:35],
                             (lizzieLet10_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet10_1_4MQNode_1QNode_Int_emitted[2]))};
  assign t4acu_destruct_d = {lizzieLet10_1_4MQNode_1QNode_Int_d[66:51],
                             (lizzieLet10_1_4MQNode_1QNode_Int_d[0] && (! lizzieLet10_1_4MQNode_1QNode_Int_emitted[3]))};
  assign lizzieLet10_1_4MQNode_1QNode_Int_done = (lizzieLet10_1_4MQNode_1QNode_Int_emitted | ({t4acu_destruct_d[0],
                                                                                               t3act_destruct_d[0],
                                                                                               t2acs_destruct_d[0],
                                                                                               t1acr_destruct_d[0]} & {t4acu_destruct_r,
                                                                                                                       t3act_destruct_r,
                                                                                                                       t2acs_destruct_r,
                                                                                                                       t1acr_destruct_r}));
  assign lizzieLet10_1_4MQNode_1QNode_Int_r = (& lizzieLet10_1_4MQNode_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet10_1_4MQNode_1QNode_Int_emitted <= (lizzieLet10_1_4MQNode_1QNode_Int_r ? 4'd0 :
                                                   lizzieLet10_1_4MQNode_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet10_1_4MQNode_2,QTree_Int) (lizzieLet10_1_4MQNode_1,QTree_Int) > [(_43,QTree_Int),
                                                                                                  (_42,QTree_Int),
                                                                                                  (lizzieLet10_1_4MQNode_1QNode_Int,QTree_Int),
                                                                                                  (_41,QTree_Int)] */
  logic [3:0] lizzieLet10_1_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_2_d[0] && lizzieLet10_1_4MQNode_1_d[0]))
      unique case (lizzieLet10_1_4MQNode_2_d[2:1])
        2'd0: lizzieLet10_1_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet10_1_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet10_1_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet10_1_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet10_1_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet10_1_4MQNode_1_onehotd = 4'd0;
  assign _43_d = {lizzieLet10_1_4MQNode_1_d[66:1],
                  lizzieLet10_1_4MQNode_1_onehotd[0]};
  assign _42_d = {lizzieLet10_1_4MQNode_1_d[66:1],
                  lizzieLet10_1_4MQNode_1_onehotd[1]};
  assign lizzieLet10_1_4MQNode_1QNode_Int_d = {lizzieLet10_1_4MQNode_1_d[66:1],
                                               lizzieLet10_1_4MQNode_1_onehotd[2]};
  assign _41_d = {lizzieLet10_1_4MQNode_1_d[66:1],
                  lizzieLet10_1_4MQNode_1_onehotd[3]};
  assign lizzieLet10_1_4MQNode_1_r = (| (lizzieLet10_1_4MQNode_1_onehotd & {_41_r,
                                                                            lizzieLet10_1_4MQNode_1QNode_Int_r,
                                                                            _42_r,
                                                                            _43_r}));
  assign lizzieLet10_1_4MQNode_2_r = lizzieLet10_1_4MQNode_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet10_1_4MQNode_3,QTree_Int) (lizzieLet10_1_3MQNode,Go) > [(lizzieLet10_1_4MQNode_3QNone_Int,Go),
                                                                                  (lizzieLet10_1_4MQNode_3QVal_Int,Go),
                                                                                  (lizzieLet10_1_4MQNode_3QNode_Int,Go),
                                                                                  (lizzieLet10_1_4MQNode_3QError_Int,Go)] */
  logic [3:0] lizzieLet10_1_3MQNode_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_3_d[0] && lizzieLet10_1_3MQNode_d[0]))
      unique case (lizzieLet10_1_4MQNode_3_d[2:1])
        2'd0: lizzieLet10_1_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet10_1_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet10_1_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet10_1_3MQNode_onehotd = 4'd8;
        default: lizzieLet10_1_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet10_1_3MQNode_onehotd = 4'd0;
  assign lizzieLet10_1_4MQNode_3QNone_Int_d = lizzieLet10_1_3MQNode_onehotd[0];
  assign lizzieLet10_1_4MQNode_3QVal_Int_d = lizzieLet10_1_3MQNode_onehotd[1];
  assign lizzieLet10_1_4MQNode_3QNode_Int_d = lizzieLet10_1_3MQNode_onehotd[2];
  assign lizzieLet10_1_4MQNode_3QError_Int_d = lizzieLet10_1_3MQNode_onehotd[3];
  assign lizzieLet10_1_3MQNode_r = (| (lizzieLet10_1_3MQNode_onehotd & {lizzieLet10_1_4MQNode_3QError_Int_r,
                                                                        lizzieLet10_1_4MQNode_3QNode_Int_r,
                                                                        lizzieLet10_1_4MQNode_3QVal_Int_r,
                                                                        lizzieLet10_1_4MQNode_3QNone_Int_r}));
  assign lizzieLet10_1_4MQNode_3_r = lizzieLet10_1_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet10_1_4MQNode_3QError_Int,Go) > [(lizzieLet10_1_4MQNode_3QError_Int_1,Go),
                                                         (lizzieLet10_1_4MQNode_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet10_1_4MQNode_3QError_Int_emitted;
  logic [1:0] lizzieLet10_1_4MQNode_3QError_Int_done;
  assign lizzieLet10_1_4MQNode_3QError_Int_1_d = (lizzieLet10_1_4MQNode_3QError_Int_d[0] && (! lizzieLet10_1_4MQNode_3QError_Int_emitted[0]));
  assign lizzieLet10_1_4MQNode_3QError_Int_2_d = (lizzieLet10_1_4MQNode_3QError_Int_d[0] && (! lizzieLet10_1_4MQNode_3QError_Int_emitted[1]));
  assign lizzieLet10_1_4MQNode_3QError_Int_done = (lizzieLet10_1_4MQNode_3QError_Int_emitted | ({lizzieLet10_1_4MQNode_3QError_Int_2_d[0],
                                                                                                 lizzieLet10_1_4MQNode_3QError_Int_1_d[0]} & {lizzieLet10_1_4MQNode_3QError_Int_2_r,
                                                                                                                                              lizzieLet10_1_4MQNode_3QError_Int_1_r}));
  assign lizzieLet10_1_4MQNode_3QError_Int_r = (& lizzieLet10_1_4MQNode_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet10_1_4MQNode_3QError_Int_emitted <= (lizzieLet10_1_4MQNode_3QError_Int_r ? 2'd0 :
                                                    lizzieLet10_1_4MQNode_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet10_1_4MQNode_3QError_Int_1,Go)] > (lizzieLet10_1_4MQNode_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet10_1_4MQNode_3QError_Int_1_d[0]}), lizzieLet10_1_4MQNode_3QError_Int_1_d);
  assign {lizzieLet10_1_4MQNode_3QError_Int_1_r} = {1 {(lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_r && lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_1_4MQNode_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet16_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_r = ((! lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_r)
        lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d <= lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet10_1_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_1_4MQNode_3QError_Int_2,Go) > (lizzieLet10_1_4MQNode_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QError_Int_2_r = ((! lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_4MQNode_3QError_Int_2_r)
        lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d <= lizzieLet10_1_4MQNode_3QError_Int_2_d;
  Go_t lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_r = (! lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_d = (lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf :
                                                         lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_r && lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_4MQNode_3QError_Int_2_argbuf_r) && (! lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_buf <= lizzieLet10_1_4MQNode_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_1_4MQNode_3QNode_Int,Go) > (lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QNode_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QNode_Int_r = ((! lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_4MQNode_3QNode_Int_r)
        lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d <= lizzieLet10_1_4MQNode_3QNode_Int_d;
  Go_t lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QNode_Int_bufchan_r = (! lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_d = (lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf :
                                                        lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_r && lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_4MQNode_3QNode_Int_1_argbuf_r) && (! lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QNode_Int_bufchan_buf <= lizzieLet10_1_4MQNode_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet10_1_4MQNode_3QNone_Int,Go) > [(lizzieLet10_1_4MQNode_3QNone_Int_1,Go),
                                                        (lizzieLet10_1_4MQNode_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet10_1_4MQNode_3QNone_Int_emitted;
  logic [1:0] lizzieLet10_1_4MQNode_3QNone_Int_done;
  assign lizzieLet10_1_4MQNode_3QNone_Int_1_d = (lizzieLet10_1_4MQNode_3QNone_Int_d[0] && (! lizzieLet10_1_4MQNode_3QNone_Int_emitted[0]));
  assign lizzieLet10_1_4MQNode_3QNone_Int_2_d = (lizzieLet10_1_4MQNode_3QNone_Int_d[0] && (! lizzieLet10_1_4MQNode_3QNone_Int_emitted[1]));
  assign lizzieLet10_1_4MQNode_3QNone_Int_done = (lizzieLet10_1_4MQNode_3QNone_Int_emitted | ({lizzieLet10_1_4MQNode_3QNone_Int_2_d[0],
                                                                                               lizzieLet10_1_4MQNode_3QNone_Int_1_d[0]} & {lizzieLet10_1_4MQNode_3QNone_Int_2_r,
                                                                                                                                           lizzieLet10_1_4MQNode_3QNone_Int_1_r}));
  assign lizzieLet10_1_4MQNode_3QNone_Int_r = (& lizzieLet10_1_4MQNode_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet10_1_4MQNode_3QNone_Int_emitted <= (lizzieLet10_1_4MQNode_3QNone_Int_r ? 2'd0 :
                                                   lizzieLet10_1_4MQNode_3QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet10_1_4MQNode_3QNone_Int_1,Go)] > (lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet10_1_4MQNode_3QNone_Int_1_d[0]}), lizzieLet10_1_4MQNode_3QNone_Int_1_d);
  assign {lizzieLet10_1_4MQNode_3QNone_Int_1_r} = {1 {(lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_r && lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet13_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_r = ((! lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_r)
        lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf :
                                   lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet10_1_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_1_4MQNode_3QNone_Int_2,Go) > (lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QNone_Int_2_r = ((! lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_4MQNode_3QNone_Int_2_r)
        lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d <= lizzieLet10_1_4MQNode_3QNone_Int_2_d;
  Go_t lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_r = (! lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_d = (lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf :
                                                        lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_r && lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_4MQNode_3QNone_Int_2_argbuf_r) && (! lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_buf <= lizzieLet10_1_4MQNode_3QNone_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet10_1_4MQNode_3QVal_Int,Go) > [(lizzieLet10_1_4MQNode_3QVal_Int_1,Go),
                                                       (lizzieLet10_1_4MQNode_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet10_1_4MQNode_3QVal_Int_emitted;
  logic [1:0] lizzieLet10_1_4MQNode_3QVal_Int_done;
  assign lizzieLet10_1_4MQNode_3QVal_Int_1_d = (lizzieLet10_1_4MQNode_3QVal_Int_d[0] && (! lizzieLet10_1_4MQNode_3QVal_Int_emitted[0]));
  assign lizzieLet10_1_4MQNode_3QVal_Int_2_d = (lizzieLet10_1_4MQNode_3QVal_Int_d[0] && (! lizzieLet10_1_4MQNode_3QVal_Int_emitted[1]));
  assign lizzieLet10_1_4MQNode_3QVal_Int_done = (lizzieLet10_1_4MQNode_3QVal_Int_emitted | ({lizzieLet10_1_4MQNode_3QVal_Int_2_d[0],
                                                                                             lizzieLet10_1_4MQNode_3QVal_Int_1_d[0]} & {lizzieLet10_1_4MQNode_3QVal_Int_2_r,
                                                                                                                                        lizzieLet10_1_4MQNode_3QVal_Int_1_r}));
  assign lizzieLet10_1_4MQNode_3QVal_Int_r = (& lizzieLet10_1_4MQNode_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet10_1_4MQNode_3QVal_Int_emitted <= (lizzieLet10_1_4MQNode_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet10_1_4MQNode_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet10_1_4MQNode_3QVal_Int_1,Go)] > (lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet10_1_4MQNode_3QVal_Int_1_d[0]}), lizzieLet10_1_4MQNode_3QVal_Int_1_d);
  assign {lizzieLet10_1_4MQNode_3QVal_Int_1_r} = {1 {(lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_r && lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet14_2_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_r = ((! lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_r)
        lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet14_2_1_argbuf_d = (lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf :
                                     lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet14_2_1_argbuf_r && lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet14_2_1_argbuf_r) && (! lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet10_1_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet10_1_4MQNode_3QVal_Int_2,Go) > (lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d;
  logic lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_r;
  assign lizzieLet10_1_4MQNode_3QVal_Int_2_r = ((! lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d[0]) || lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet10_1_4MQNode_3QVal_Int_2_r)
        lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d <= lizzieLet10_1_4MQNode_3QVal_Int_2_d;
  Go_t lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf;
  assign lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_r = (! lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_d = (lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf[0] ? lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf :
                                                       lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_r && lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet10_1_4MQNode_3QVal_Int_2_argbuf_r) && (! lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_buf <= lizzieLet10_1_4MQNode_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_4MQNode_4,QTree_Int) (lizzieLet10_1_6MQNode,Pointer_CTmain_mask_Int) > [(lizzieLet10_1_4MQNode_4QNone_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet10_1_4MQNode_4QVal_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet10_1_4MQNode_4QNode_Int,Pointer_CTmain_mask_Int),
                                                                                                                            (lizzieLet10_1_4MQNode_4QError_Int,Pointer_CTmain_mask_Int)] */
  logic [3:0] lizzieLet10_1_6MQNode_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_4_d[0] && lizzieLet10_1_6MQNode_d[0]))
      unique case (lizzieLet10_1_4MQNode_4_d[2:1])
        2'd0: lizzieLet10_1_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet10_1_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet10_1_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet10_1_6MQNode_onehotd = 4'd8;
        default: lizzieLet10_1_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet10_1_6MQNode_onehotd = 4'd0;
  assign lizzieLet10_1_4MQNode_4QNone_Int_d = {lizzieLet10_1_6MQNode_d[16:1],
                                               lizzieLet10_1_6MQNode_onehotd[0]};
  assign lizzieLet10_1_4MQNode_4QVal_Int_d = {lizzieLet10_1_6MQNode_d[16:1],
                                              lizzieLet10_1_6MQNode_onehotd[1]};
  assign lizzieLet10_1_4MQNode_4QNode_Int_d = {lizzieLet10_1_6MQNode_d[16:1],
                                               lizzieLet10_1_6MQNode_onehotd[2]};
  assign lizzieLet10_1_4MQNode_4QError_Int_d = {lizzieLet10_1_6MQNode_d[16:1],
                                                lizzieLet10_1_6MQNode_onehotd[3]};
  assign lizzieLet10_1_6MQNode_r = (| (lizzieLet10_1_6MQNode_onehotd & {lizzieLet10_1_4MQNode_4QError_Int_r,
                                                                        lizzieLet10_1_4MQNode_4QNode_Int_r,
                                                                        lizzieLet10_1_4MQNode_4QVal_Int_r,
                                                                        lizzieLet10_1_4MQNode_4QNone_Int_r}));
  assign lizzieLet10_1_4MQNode_4_r = lizzieLet10_1_6MQNode_r;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_4MQNode_4QError_Int,Pointer_CTmain_mask_Int) > (lizzieLet10_1_4MQNode_4QError_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QError_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_4QError_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_4QError_Int_r = ((! lizzieLet10_1_4MQNode_4QError_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_4MQNode_4QError_Int_r)
        lizzieLet10_1_4MQNode_4QError_Int_bufchan_d <= lizzieLet10_1_4MQNode_4QError_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_4QError_Int_bufchan_r = (! lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_d = (lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf :
                                                         lizzieLet10_1_4MQNode_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_r && lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_4MQNode_4QError_Int_1_argbuf_r) && (! lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_4QError_Int_bufchan_buf <= lizzieLet10_1_4MQNode_4QError_Int_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int3) : [(lizzieLet10_1_4MQNode_4QNode_Int,Pointer_CTmain_mask_Int),
                                    (t1acr_destruct,Pointer_QTree_Int),
                                    (lizzieLet10_1_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                    (t2acs_destruct,Pointer_QTree_Int),
                                    (lizzieLet10_1_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                    (t3act_destruct,Pointer_QTree_Int),
                                    (lizzieLet10_1_4MQNode_7QNode_Int,Pointer_MaskQTree)] > (lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3,CTmain_mask_Int) */
  assign lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d = Lcall_main_mask_Int3_dc((& {lizzieLet10_1_4MQNode_4QNode_Int_d[0],
                                                                                                                                                                                                                           t1acr_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet10_1_4MQNode_5QNode_Int_d[0],
                                                                                                                                                                                                                           t2acs_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet10_1_4MQNode_6QNode_Int_d[0],
                                                                                                                                                                                                                           t3act_destruct_d[0],
                                                                                                                                                                                                                           lizzieLet10_1_4MQNode_7QNode_Int_d[0]}), lizzieLet10_1_4MQNode_4QNode_Int_d, t1acr_destruct_d, lizzieLet10_1_4MQNode_5QNode_Int_d, t2acs_destruct_d, lizzieLet10_1_4MQNode_6QNode_Int_d, t3act_destruct_d, lizzieLet10_1_4MQNode_7QNode_Int_d);
  assign {lizzieLet10_1_4MQNode_4QNode_Int_r,
          t1acr_destruct_r,
          lizzieLet10_1_4MQNode_5QNode_Int_r,
          t2acs_destruct_r,
          lizzieLet10_1_4MQNode_6QNode_Int_r,
          t3act_destruct_r,
          lizzieLet10_1_4MQNode_7QNode_Int_r} = {7 {(lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r && lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3,CTmain_mask_Int) > (lizzieLet15_1_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d;
  logic lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r;
  assign lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r = ((! lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d[0]) || lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d <= {115'd0,
                                                                                                                                                                                                      1'd0};
    else
      if (lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_r)
        lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d <= lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_d;
  CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf;
  assign lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_r = (! lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0] ? lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf :
                                     lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                        1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                          1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_buf <= lizzieLet10_1_4MQNode_4QNode_Int_1t1acr_1lizzieLet10_1_4MQNode_5QNode_Int_1t2acs_1lizzieLet10_1_4MQNode_6QNode_Int_1t3act_1lizzieLet10_1_4MQNode_7QNode_Int_1Lcall_main_mask_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_4MQNode_4QNone_Int,Pointer_CTmain_mask_Int) > (lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_4QNone_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_4QNone_Int_r = ((! lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_4MQNode_4QNone_Int_r)
        lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d <= lizzieLet10_1_4MQNode_4QNone_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_4QNone_Int_bufchan_r = (! lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_d = (lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf :
                                                        lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_r && lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_4MQNode_4QNone_Int_1_argbuf_r) && (! lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_4QNone_Int_bufchan_buf <= lizzieLet10_1_4MQNode_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_4MQNode_4QVal_Int,Pointer_CTmain_mask_Int) > (lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_4QVal_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_4QVal_Int_r = ((! lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_4MQNode_4QVal_Int_r)
        lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d <= lizzieLet10_1_4MQNode_4QVal_Int_d;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_4QVal_Int_bufchan_r = (! lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_d = (lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf :
                                                       lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_r && lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_4MQNode_4QVal_Int_1_argbuf_r) && (! lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_4QVal_Int_bufchan_buf <= lizzieLet10_1_4MQNode_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet10_1_4MQNode_5,QTree_Int) (q1acm_destruct,Pointer_MaskQTree) > [(_40,Pointer_MaskQTree),
                                                                                                         (_39,Pointer_MaskQTree),
                                                                                                         (lizzieLet10_1_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                                                                                         (_38,Pointer_MaskQTree)] */
  logic [3:0] q1acm_destruct_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_5_d[0] && q1acm_destruct_d[0]))
      unique case (lizzieLet10_1_4MQNode_5_d[2:1])
        2'd0: q1acm_destruct_onehotd = 4'd1;
        2'd1: q1acm_destruct_onehotd = 4'd2;
        2'd2: q1acm_destruct_onehotd = 4'd4;
        2'd3: q1acm_destruct_onehotd = 4'd8;
        default: q1acm_destruct_onehotd = 4'd0;
      endcase
    else q1acm_destruct_onehotd = 4'd0;
  assign _40_d = {q1acm_destruct_d[16:1], q1acm_destruct_onehotd[0]};
  assign _39_d = {q1acm_destruct_d[16:1], q1acm_destruct_onehotd[1]};
  assign lizzieLet10_1_4MQNode_5QNode_Int_d = {q1acm_destruct_d[16:1],
                                               q1acm_destruct_onehotd[2]};
  assign _38_d = {q1acm_destruct_d[16:1], q1acm_destruct_onehotd[3]};
  assign q1acm_destruct_r = (| (q1acm_destruct_onehotd & {_38_r,
                                                          lizzieLet10_1_4MQNode_5QNode_Int_r,
                                                          _39_r,
                                                          _40_r}));
  assign lizzieLet10_1_4MQNode_5_r = q1acm_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet10_1_4MQNode_6,QTree_Int) (q2acn_destruct,Pointer_MaskQTree) > [(_37,Pointer_MaskQTree),
                                                                                                         (_36,Pointer_MaskQTree),
                                                                                                         (lizzieLet10_1_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                                                                                         (_35,Pointer_MaskQTree)] */
  logic [3:0] q2acn_destruct_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_6_d[0] && q2acn_destruct_d[0]))
      unique case (lizzieLet10_1_4MQNode_6_d[2:1])
        2'd0: q2acn_destruct_onehotd = 4'd1;
        2'd1: q2acn_destruct_onehotd = 4'd2;
        2'd2: q2acn_destruct_onehotd = 4'd4;
        2'd3: q2acn_destruct_onehotd = 4'd8;
        default: q2acn_destruct_onehotd = 4'd0;
      endcase
    else q2acn_destruct_onehotd = 4'd0;
  assign _37_d = {q2acn_destruct_d[16:1], q2acn_destruct_onehotd[0]};
  assign _36_d = {q2acn_destruct_d[16:1], q2acn_destruct_onehotd[1]};
  assign lizzieLet10_1_4MQNode_6QNode_Int_d = {q2acn_destruct_d[16:1],
                                               q2acn_destruct_onehotd[2]};
  assign _35_d = {q2acn_destruct_d[16:1], q2acn_destruct_onehotd[3]};
  assign q2acn_destruct_r = (| (q2acn_destruct_onehotd & {_35_r,
                                                          lizzieLet10_1_4MQNode_6QNode_Int_r,
                                                          _36_r,
                                                          _37_r}));
  assign lizzieLet10_1_4MQNode_6_r = q2acn_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet10_1_4MQNode_7,QTree_Int) (q3aco_destruct,Pointer_MaskQTree) > [(_34,Pointer_MaskQTree),
                                                                                                         (_33,Pointer_MaskQTree),
                                                                                                         (lizzieLet10_1_4MQNode_7QNode_Int,Pointer_MaskQTree),
                                                                                                         (_32,Pointer_MaskQTree)] */
  logic [3:0] q3aco_destruct_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_7_d[0] && q3aco_destruct_d[0]))
      unique case (lizzieLet10_1_4MQNode_7_d[2:1])
        2'd0: q3aco_destruct_onehotd = 4'd1;
        2'd1: q3aco_destruct_onehotd = 4'd2;
        2'd2: q3aco_destruct_onehotd = 4'd4;
        2'd3: q3aco_destruct_onehotd = 4'd8;
        default: q3aco_destruct_onehotd = 4'd0;
      endcase
    else q3aco_destruct_onehotd = 4'd0;
  assign _34_d = {q3aco_destruct_d[16:1], q3aco_destruct_onehotd[0]};
  assign _33_d = {q3aco_destruct_d[16:1], q3aco_destruct_onehotd[1]};
  assign lizzieLet10_1_4MQNode_7QNode_Int_d = {q3aco_destruct_d[16:1],
                                               q3aco_destruct_onehotd[2]};
  assign _32_d = {q3aco_destruct_d[16:1], q3aco_destruct_onehotd[3]};
  assign q3aco_destruct_r = (| (q3aco_destruct_onehotd & {_32_r,
                                                          lizzieLet10_1_4MQNode_7QNode_Int_r,
                                                          _33_r,
                                                          _34_r}));
  assign lizzieLet10_1_4MQNode_7_r = q3aco_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet10_1_4MQNode_8,QTree_Int) (q4acp_destruct,Pointer_MaskQTree) > [(_31,Pointer_MaskQTree),
                                                                                                         (_30,Pointer_MaskQTree),
                                                                                                         (lizzieLet10_1_4MQNode_8QNode_Int,Pointer_MaskQTree),
                                                                                                         (_29,Pointer_MaskQTree)] */
  logic [3:0] q4acp_destruct_onehotd;
  always_comb
    if ((lizzieLet10_1_4MQNode_8_d[0] && q4acp_destruct_d[0]))
      unique case (lizzieLet10_1_4MQNode_8_d[2:1])
        2'd0: q4acp_destruct_onehotd = 4'd1;
        2'd1: q4acp_destruct_onehotd = 4'd2;
        2'd2: q4acp_destruct_onehotd = 4'd4;
        2'd3: q4acp_destruct_onehotd = 4'd8;
        default: q4acp_destruct_onehotd = 4'd0;
      endcase
    else q4acp_destruct_onehotd = 4'd0;
  assign _31_d = {q4acp_destruct_d[16:1], q4acp_destruct_onehotd[0]};
  assign _30_d = {q4acp_destruct_d[16:1], q4acp_destruct_onehotd[1]};
  assign lizzieLet10_1_4MQNode_8QNode_Int_d = {q4acp_destruct_d[16:1],
                                               q4acp_destruct_onehotd[2]};
  assign _29_d = {q4acp_destruct_d[16:1], q4acp_destruct_onehotd[3]};
  assign q4acp_destruct_r = (| (q4acp_destruct_onehotd & {_29_r,
                                                          lizzieLet10_1_4MQNode_8QNode_Int_r,
                                                          _30_r,
                                                          _31_r}));
  assign lizzieLet10_1_4MQNode_8_r = q4acp_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet10_1_4MQNode_8QNode_Int,Pointer_MaskQTree) > (lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d;
  logic lizzieLet10_1_4MQNode_8QNode_Int_bufchan_r;
  assign lizzieLet10_1_4MQNode_8QNode_Int_r = ((! lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d[0]) || lizzieLet10_1_4MQNode_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_4MQNode_8QNode_Int_r)
        lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d <= lizzieLet10_1_4MQNode_8QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf;
  assign lizzieLet10_1_4MQNode_8QNode_Int_bufchan_r = (! lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_d = (lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf[0] ? lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf :
                                                        lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_r && lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf[0]))
        lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_4MQNode_8QNode_Int_1_argbuf_r) && (! lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf[0])))
        lizzieLet10_1_4MQNode_8QNode_Int_bufchan_buf <= lizzieLet10_1_4MQNode_8QNode_Int_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Int) : (lizzieLet10_1_5,MaskQTree) (mack_2,Pointer_QTree_Int) > [(_28,Pointer_QTree_Int),
                                                                                         (lizzieLet10_1_5MQVal,Pointer_QTree_Int),
                                                                                         (_27,Pointer_QTree_Int)] */
  logic [2:0] mack_2_onehotd;
  always_comb
    if ((lizzieLet10_1_5_d[0] && mack_2_d[0]))
      unique case (lizzieLet10_1_5_d[2:1])
        2'd0: mack_2_onehotd = 3'd1;
        2'd1: mack_2_onehotd = 3'd2;
        2'd2: mack_2_onehotd = 3'd4;
        default: mack_2_onehotd = 3'd0;
      endcase
    else mack_2_onehotd = 3'd0;
  assign _28_d = {mack_2_d[16:1], mack_2_onehotd[0]};
  assign lizzieLet10_1_5MQVal_d = {mack_2_d[16:1],
                                   mack_2_onehotd[1]};
  assign _27_d = {mack_2_d[16:1], mack_2_onehotd[2]};
  assign mack_2_r = (| (mack_2_onehotd & {_27_r,
                                          lizzieLet10_1_5MQVal_r,
                                          _28_r}));
  assign lizzieLet10_1_5_r = mack_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet10_1_5MQVal,Pointer_QTree_Int) > (lizzieLet10_1_5MQVal_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet10_1_5MQVal_bufchan_d;
  logic lizzieLet10_1_5MQVal_bufchan_r;
  assign lizzieLet10_1_5MQVal_r = ((! lizzieLet10_1_5MQVal_bufchan_d[0]) || lizzieLet10_1_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_5MQVal_r)
        lizzieLet10_1_5MQVal_bufchan_d <= lizzieLet10_1_5MQVal_d;
  Pointer_QTree_Int_t lizzieLet10_1_5MQVal_bufchan_buf;
  assign lizzieLet10_1_5MQVal_bufchan_r = (! lizzieLet10_1_5MQVal_bufchan_buf[0]);
  assign lizzieLet10_1_5MQVal_1_argbuf_d = (lizzieLet10_1_5MQVal_bufchan_buf[0] ? lizzieLet10_1_5MQVal_bufchan_buf :
                                            lizzieLet10_1_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_5MQVal_1_argbuf_r && lizzieLet10_1_5MQVal_bufchan_buf[0]))
        lizzieLet10_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_5MQVal_1_argbuf_r) && (! lizzieLet10_1_5MQVal_bufchan_buf[0])))
        lizzieLet10_1_5MQVal_bufchan_buf <= lizzieLet10_1_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_6,MaskQTree) (sc_0_2_goMux_mux,Pointer_CTmain_mask_Int) > [(lizzieLet10_1_6MQNone,Pointer_CTmain_mask_Int),
                                                                                                               (lizzieLet10_1_6MQVal,Pointer_CTmain_mask_Int),
                                                                                                               (lizzieLet10_1_6MQNode,Pointer_CTmain_mask_Int)] */
  logic [2:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet10_1_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet10_1_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 3'd4;
        default: sc_0_2_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 3'd0;
  assign lizzieLet10_1_6MQNone_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet10_1_6MQVal_d = {sc_0_2_goMux_mux_d[16:1],
                                   sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet10_1_6MQNode_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[2]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet10_1_6MQNode_r,
                                                              lizzieLet10_1_6MQVal_r,
                                                              lizzieLet10_1_6MQNone_r}));
  assign lizzieLet10_1_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_6MQNone,Pointer_CTmain_mask_Int) > (lizzieLet10_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQNone_bufchan_d;
  logic lizzieLet10_1_6MQNone_bufchan_r;
  assign lizzieLet10_1_6MQNone_r = ((! lizzieLet10_1_6MQNone_bufchan_d[0]) || lizzieLet10_1_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_6MQNone_r)
        lizzieLet10_1_6MQNone_bufchan_d <= lizzieLet10_1_6MQNone_d;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQNone_bufchan_buf;
  assign lizzieLet10_1_6MQNone_bufchan_r = (! lizzieLet10_1_6MQNone_bufchan_buf[0]);
  assign lizzieLet10_1_6MQNone_1_argbuf_d = (lizzieLet10_1_6MQNone_bufchan_buf[0] ? lizzieLet10_1_6MQNone_bufchan_buf :
                                             lizzieLet10_1_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_6MQNone_1_argbuf_r && lizzieLet10_1_6MQNone_bufchan_buf[0]))
        lizzieLet10_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_6MQNone_1_argbuf_r) && (! lizzieLet10_1_6MQNone_bufchan_buf[0])))
        lizzieLet10_1_6MQNone_bufchan_buf <= lizzieLet10_1_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (lizzieLet10_1_6MQVal,Pointer_CTmain_mask_Int) > (lizzieLet10_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQVal_bufchan_d;
  logic lizzieLet10_1_6MQVal_bufchan_r;
  assign lizzieLet10_1_6MQVal_r = ((! lizzieLet10_1_6MQVal_bufchan_d[0]) || lizzieLet10_1_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet10_1_6MQVal_r)
        lizzieLet10_1_6MQVal_bufchan_d <= lizzieLet10_1_6MQVal_d;
  Pointer_CTmain_mask_Int_t lizzieLet10_1_6MQVal_bufchan_buf;
  assign lizzieLet10_1_6MQVal_bufchan_r = (! lizzieLet10_1_6MQVal_bufchan_buf[0]);
  assign lizzieLet10_1_6MQVal_1_argbuf_d = (lizzieLet10_1_6MQVal_bufchan_buf[0] ? lizzieLet10_1_6MQVal_bufchan_buf :
                                            lizzieLet10_1_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet10_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_6MQVal_1_argbuf_r && lizzieLet10_1_6MQVal_bufchan_buf[0]))
        lizzieLet10_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_6MQVal_1_argbuf_r) && (! lizzieLet10_1_6MQVal_bufchan_buf[0])))
        lizzieLet10_1_6MQVal_bufchan_buf <= lizzieLet10_1_6MQVal_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_1QNode_Int,QTree_Int) > [(q1acH_destruct,Pointer_QTree_Int),
                                                                  (q2acI_destruct,Pointer_QTree_Int),
                                                                  (q3acJ_destruct,Pointer_QTree_Int),
                                                                  (q4acK_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_1QNode_Int_done;
  assign q1acH_destruct_d = {lizzieLet17_1QNode_Int_d[18:3],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[0]))};
  assign q2acI_destruct_d = {lizzieLet17_1QNode_Int_d[34:19],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[1]))};
  assign q3acJ_destruct_d = {lizzieLet17_1QNode_Int_d[50:35],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[2]))};
  assign q4acK_destruct_d = {lizzieLet17_1QNode_Int_d[66:51],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[3]))};
  assign lizzieLet17_1QNode_Int_done = (lizzieLet17_1QNode_Int_emitted | ({q4acK_destruct_d[0],
                                                                           q3acJ_destruct_d[0],
                                                                           q2acI_destruct_d[0],
                                                                           q1acH_destruct_d[0]} & {q4acK_destruct_r,
                                                                                                   q3acJ_destruct_r,
                                                                                                   q2acI_destruct_r,
                                                                                                   q1acH_destruct_r}));
  assign lizzieLet17_1QNode_Int_r = (& lizzieLet17_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_1QNode_Int_emitted <= (lizzieLet17_1QNode_Int_r ? 4'd0 :
                                         lizzieLet17_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_1QVal_Int,QTree_Int) > [(vacG_destruct,Int)] */
  assign vacG_destruct_d = {lizzieLet17_1QVal_Int_d[34:3],
                            lizzieLet17_1QVal_Int_d[0]};
  assign lizzieLet17_1QVal_Int_r = vacG_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_2,QTree_Int) (lizzieLet17_1,QTree_Int) > [(_26,QTree_Int),
                                                                              (lizzieLet17_1QVal_Int,QTree_Int),
                                                                              (lizzieLet17_1QNode_Int,QTree_Int),
                                                                              (_25,QTree_Int)] */
  logic [3:0] lizzieLet17_1_onehotd;
  always_comb
    if ((lizzieLet17_2_d[0] && lizzieLet17_1_d[0]))
      unique case (lizzieLet17_2_d[2:1])
        2'd0: lizzieLet17_1_onehotd = 4'd1;
        2'd1: lizzieLet17_1_onehotd = 4'd2;
        2'd2: lizzieLet17_1_onehotd = 4'd4;
        2'd3: lizzieLet17_1_onehotd = 4'd8;
        default: lizzieLet17_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_1_onehotd = 4'd0;
  assign _26_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[0]};
  assign lizzieLet17_1QVal_Int_d = {lizzieLet17_1_d[66:1],
                                    lizzieLet17_1_onehotd[1]};
  assign lizzieLet17_1QNode_Int_d = {lizzieLet17_1_d[66:1],
                                     lizzieLet17_1_onehotd[2]};
  assign _25_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[3]};
  assign lizzieLet17_1_r = (| (lizzieLet17_1_onehotd & {_25_r,
                                                        lizzieLet17_1QNode_Int_r,
                                                        lizzieLet17_1QVal_Int_r,
                                                        _26_r}));
  assign lizzieLet17_2_r = lizzieLet17_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet17_3,QTree_Int) (gacD_goMux_mux,MyDTInt_Int_Int) > [(_24,MyDTInt_Int_Int),
                                                                                           (lizzieLet17_3QVal_Int,MyDTInt_Int_Int),
                                                                                           (lizzieLet17_3QNode_Int,MyDTInt_Int_Int),
                                                                                           (_23,MyDTInt_Int_Int)] */
  logic [3:0] gacD_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_3_d[0] && gacD_goMux_mux_d[0]))
      unique case (lizzieLet17_3_d[2:1])
        2'd0: gacD_goMux_mux_onehotd = 4'd1;
        2'd1: gacD_goMux_mux_onehotd = 4'd2;
        2'd2: gacD_goMux_mux_onehotd = 4'd4;
        2'd3: gacD_goMux_mux_onehotd = 4'd8;
        default: gacD_goMux_mux_onehotd = 4'd0;
      endcase
    else gacD_goMux_mux_onehotd = 4'd0;
  assign _24_d = gacD_goMux_mux_onehotd[0];
  assign lizzieLet17_3QVal_Int_d = gacD_goMux_mux_onehotd[1];
  assign lizzieLet17_3QNode_Int_d = gacD_goMux_mux_onehotd[2];
  assign _23_d = gacD_goMux_mux_onehotd[3];
  assign gacD_goMux_mux_r = (| (gacD_goMux_mux_onehotd & {_23_r,
                                                          lizzieLet17_3QNode_Int_r,
                                                          lizzieLet17_3QVal_Int_r,
                                                          _24_r}));
  assign lizzieLet17_3_r = gacD_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet17_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet17_3QNode_Int_1,MyDTInt_Int_Int),
                                                                        (lizzieLet17_3QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet17_3QNode_Int_emitted;
  logic [1:0] lizzieLet17_3QNode_Int_done;
  assign lizzieLet17_3QNode_Int_1_d = (lizzieLet17_3QNode_Int_d[0] && (! lizzieLet17_3QNode_Int_emitted[0]));
  assign lizzieLet17_3QNode_Int_2_d = (lizzieLet17_3QNode_Int_d[0] && (! lizzieLet17_3QNode_Int_emitted[1]));
  assign lizzieLet17_3QNode_Int_done = (lizzieLet17_3QNode_Int_emitted | ({lizzieLet17_3QNode_Int_2_d[0],
                                                                           lizzieLet17_3QNode_Int_1_d[0]} & {lizzieLet17_3QNode_Int_2_r,
                                                                                                             lizzieLet17_3QNode_Int_1_r}));
  assign lizzieLet17_3QNode_Int_r = (& lizzieLet17_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_3QNode_Int_emitted <= (lizzieLet17_3QNode_Int_r ? 2'd0 :
                                         lizzieLet17_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_3QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet17_3QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_2_bufchan_d;
  logic lizzieLet17_3QNode_Int_2_bufchan_r;
  assign lizzieLet17_3QNode_Int_2_r = ((! lizzieLet17_3QNode_Int_2_bufchan_d[0]) || lizzieLet17_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_3QNode_Int_2_r)
        lizzieLet17_3QNode_Int_2_bufchan_d <= lizzieLet17_3QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet17_3QNode_Int_2_bufchan_buf;
  assign lizzieLet17_3QNode_Int_2_bufchan_r = (! lizzieLet17_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_3QNode_Int_2_argbuf_d = (lizzieLet17_3QNode_Int_2_bufchan_buf[0] ? lizzieLet17_3QNode_Int_2_bufchan_buf :
                                              lizzieLet17_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_3QNode_Int_2_argbuf_r && lizzieLet17_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_3QNode_Int_2_argbuf_r) && (! lizzieLet17_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_3QNode_Int_2_bufchan_buf <= lizzieLet17_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet17_3QVal_Int,MyDTInt_Int_Int) > (lizzieLet17_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet17_3QVal_Int_bufchan_d;
  logic lizzieLet17_3QVal_Int_bufchan_r;
  assign lizzieLet17_3QVal_Int_r = ((! lizzieLet17_3QVal_Int_bufchan_d[0]) || lizzieLet17_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_3QVal_Int_r)
        lizzieLet17_3QVal_Int_bufchan_d <= lizzieLet17_3QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet17_3QVal_Int_bufchan_buf;
  assign lizzieLet17_3QVal_Int_bufchan_r = (! lizzieLet17_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_3QVal_Int_1_argbuf_d = (lizzieLet17_3QVal_Int_bufchan_buf[0] ? lizzieLet17_3QVal_Int_bufchan_buf :
                                             lizzieLet17_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_3QVal_Int_1_argbuf_r && lizzieLet17_3QVal_Int_bufchan_buf[0]))
        lizzieLet17_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_3QVal_Int_1_argbuf_r) && (! lizzieLet17_3QVal_Int_bufchan_buf[0])))
        lizzieLet17_3QVal_Int_bufchan_buf <= lizzieLet17_3QVal_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet17_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet17_7QVal_Int_1_argbuf,Int),
                                              (vacG_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet17_3QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet17_7QVal_Int_1_argbuf_d[0],
                                                                                                        vacG_1_argbuf_d[0]}), lizzieLet17_3QVal_Int_1_argbuf_d, lizzieLet17_7QVal_Int_1_argbuf_d, vacG_1_argbuf_d);
  assign {lizzieLet17_3QVal_Int_1_argbuf_r,
          lizzieLet17_7QVal_Int_1_argbuf_r,
          vacG_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_4,QTree_Int) (go_11_goMux_data,Go) > [(lizzieLet17_4QNone_Int,Go),
                                                                   (lizzieLet17_4QVal_Int,Go),
                                                                   (lizzieLet17_4QNode_Int,Go),
                                                                   (lizzieLet17_4QError_Int,Go)] */
  logic [3:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet17_4_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet17_4_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 4'd1;
        2'd1: go_11_goMux_data_onehotd = 4'd2;
        2'd2: go_11_goMux_data_onehotd = 4'd4;
        2'd3: go_11_goMux_data_onehotd = 4'd8;
        default: go_11_goMux_data_onehotd = 4'd0;
      endcase
    else go_11_goMux_data_onehotd = 4'd0;
  assign lizzieLet17_4QNone_Int_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet17_4QVal_Int_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet17_4QNode_Int_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet17_4QError_Int_d = go_11_goMux_data_onehotd[3];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet17_4QError_Int_r,
                                                              lizzieLet17_4QNode_Int_r,
                                                              lizzieLet17_4QVal_Int_r,
                                                              lizzieLet17_4QNone_Int_r}));
  assign lizzieLet17_4_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet17_4QError_Int,Go) > [(lizzieLet17_4QError_Int_1,Go),
                                               (lizzieLet17_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_4QError_Int_emitted;
  logic [1:0] lizzieLet17_4QError_Int_done;
  assign lizzieLet17_4QError_Int_1_d = (lizzieLet17_4QError_Int_d[0] && (! lizzieLet17_4QError_Int_emitted[0]));
  assign lizzieLet17_4QError_Int_2_d = (lizzieLet17_4QError_Int_d[0] && (! lizzieLet17_4QError_Int_emitted[1]));
  assign lizzieLet17_4QError_Int_done = (lizzieLet17_4QError_Int_emitted | ({lizzieLet17_4QError_Int_2_d[0],
                                                                             lizzieLet17_4QError_Int_1_d[0]} & {lizzieLet17_4QError_Int_2_r,
                                                                                                                lizzieLet17_4QError_Int_1_r}));
  assign lizzieLet17_4QError_Int_r = (& lizzieLet17_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_4QError_Int_emitted <= (lizzieLet17_4QError_Int_r ? 2'd0 :
                                          lizzieLet17_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet17_4QError_Int_1,Go)] > (lizzieLet17_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet17_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet17_4QError_Int_1_d[0]}), lizzieLet17_4QError_Int_1_d);
  assign {lizzieLet17_4QError_Int_1_r} = {1 {(lizzieLet17_4QError_Int_1QError_Int_r && lizzieLet17_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet22_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet17_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet17_4QError_Int_1QError_Int_r = ((! lizzieLet17_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet17_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_4QError_Int_1QError_Int_r)
        lizzieLet17_4QError_Int_1QError_Int_bufchan_d <= lizzieLet17_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet17_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet17_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet17_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet17_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet17_4QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet17_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet17_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet17_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet17_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet17_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet17_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QError_Int_2,Go) > (lizzieLet17_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_4QError_Int_2_bufchan_d;
  logic lizzieLet17_4QError_Int_2_bufchan_r;
  assign lizzieLet17_4QError_Int_2_r = ((! lizzieLet17_4QError_Int_2_bufchan_d[0]) || lizzieLet17_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QError_Int_2_r)
        lizzieLet17_4QError_Int_2_bufchan_d <= lizzieLet17_4QError_Int_2_d;
  Go_t lizzieLet17_4QError_Int_2_bufchan_buf;
  assign lizzieLet17_4QError_Int_2_bufchan_r = (! lizzieLet17_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_4QError_Int_2_argbuf_d = (lizzieLet17_4QError_Int_2_bufchan_buf[0] ? lizzieLet17_4QError_Int_2_bufchan_buf :
                                               lizzieLet17_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QError_Int_2_argbuf_r && lizzieLet17_4QError_Int_2_bufchan_buf[0]))
        lizzieLet17_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QError_Int_2_argbuf_r) && (! lizzieLet17_4QError_Int_2_bufchan_buf[0])))
        lizzieLet17_4QError_Int_2_bufchan_buf <= lizzieLet17_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QNode_Int,Go) > (lizzieLet17_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet17_4QNode_Int_bufchan_d;
  logic lizzieLet17_4QNode_Int_bufchan_r;
  assign lizzieLet17_4QNode_Int_r = ((! lizzieLet17_4QNode_Int_bufchan_d[0]) || lizzieLet17_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QNode_Int_r)
        lizzieLet17_4QNode_Int_bufchan_d <= lizzieLet17_4QNode_Int_d;
  Go_t lizzieLet17_4QNode_Int_bufchan_buf;
  assign lizzieLet17_4QNode_Int_bufchan_r = (! lizzieLet17_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_4QNode_Int_1_argbuf_d = (lizzieLet17_4QNode_Int_bufchan_buf[0] ? lizzieLet17_4QNode_Int_bufchan_buf :
                                              lizzieLet17_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QNode_Int_1_argbuf_r && lizzieLet17_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QNode_Int_1_argbuf_r) && (! lizzieLet17_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_4QNode_Int_bufchan_buf <= lizzieLet17_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_4QNone_Int,Go) > [(lizzieLet17_4QNone_Int_1,Go),
                                              (lizzieLet17_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet17_4QNone_Int_emitted;
  logic [1:0] lizzieLet17_4QNone_Int_done;
  assign lizzieLet17_4QNone_Int_1_d = (lizzieLet17_4QNone_Int_d[0] && (! lizzieLet17_4QNone_Int_emitted[0]));
  assign lizzieLet17_4QNone_Int_2_d = (lizzieLet17_4QNone_Int_d[0] && (! lizzieLet17_4QNone_Int_emitted[1]));
  assign lizzieLet17_4QNone_Int_done = (lizzieLet17_4QNone_Int_emitted | ({lizzieLet17_4QNone_Int_2_d[0],
                                                                           lizzieLet17_4QNone_Int_1_d[0]} & {lizzieLet17_4QNone_Int_2_r,
                                                                                                             lizzieLet17_4QNone_Int_1_r}));
  assign lizzieLet17_4QNone_Int_r = (& lizzieLet17_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet17_4QNone_Int_emitted <= (lizzieLet17_4QNone_Int_r ? 2'd0 :
                                         lizzieLet17_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet17_4QNone_Int_1,Go)] > (lizzieLet17_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet17_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet17_4QNone_Int_1_d[0]}), lizzieLet17_4QNone_Int_1_d);
  assign {lizzieLet17_4QNone_Int_1_r} = {1 {(lizzieLet17_4QNone_Int_1QNone_Int_r && lizzieLet17_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet17_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet18_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet17_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet17_4QNone_Int_1QNone_Int_r = ((! lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet17_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_4QNone_Int_1QNone_Int_r)
        lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet17_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet17_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf :
                                   lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet17_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet17_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QNone_Int_2,Go) > (lizzieLet17_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet17_4QNone_Int_2_bufchan_d;
  logic lizzieLet17_4QNone_Int_2_bufchan_r;
  assign lizzieLet17_4QNone_Int_2_r = ((! lizzieLet17_4QNone_Int_2_bufchan_d[0]) || lizzieLet17_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QNone_Int_2_r)
        lizzieLet17_4QNone_Int_2_bufchan_d <= lizzieLet17_4QNone_Int_2_d;
  Go_t lizzieLet17_4QNone_Int_2_bufchan_buf;
  assign lizzieLet17_4QNone_Int_2_bufchan_r = (! lizzieLet17_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet17_4QNone_Int_2_argbuf_d = (lizzieLet17_4QNone_Int_2_bufchan_buf[0] ? lizzieLet17_4QNone_Int_2_bufchan_buf :
                                              lizzieLet17_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QNone_Int_2_argbuf_r && lizzieLet17_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet17_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QNone_Int_2_argbuf_r) && (! lizzieLet17_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet17_4QNone_Int_2_bufchan_buf <= lizzieLet17_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet17_4QNone_Int_2_argbuf,Go),
                           (lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf,Go),
                           (es_0_2_1MyFalse_1_argbuf,Go),
                           (es_0_2_1MyTrue_2_argbuf,Go),
                           (lizzieLet17_4QError_Int_2_argbuf,Go)] > (go_18_goMux_choice,C5) (go_18_goMux_data,Go) */
  logic [4:0] lizzieLet17_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet17_4QNone_Int_2_argbuf_select_d = ((| lizzieLet17_4QNone_Int_2_argbuf_select_q) ? lizzieLet17_4QNone_Int_2_argbuf_select_q :
                                                     (lizzieLet17_4QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                      (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d [0] ? 5'd2 :
                                                       (es_0_2_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                        (es_0_2_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                         (lizzieLet17_4QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] lizzieLet17_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet17_4QNone_Int_2_argbuf_select_q <= (lizzieLet17_4QNone_Int_2_argbuf_done ? 5'd0 :
                                                   lizzieLet17_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet17_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet17_4QNone_Int_2_argbuf_emit_q <= (lizzieLet17_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                 lizzieLet17_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet17_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet17_4QNone_Int_2_argbuf_emit_d = (lizzieLet17_4QNone_Int_2_argbuf_emit_q | ({go_18_goMux_choice_d[0],
                                                                                              go_18_goMux_data_d[0]} & {go_18_goMux_choice_r,
                                                                                                                        go_18_goMux_data_r}));
  logic lizzieLet17_4QNone_Int_2_argbuf_done;
  assign lizzieLet17_4QNone_Int_2_argbuf_done = (& lizzieLet17_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet17_4QError_Int_2_argbuf_r,
          es_0_2_1MyTrue_2_argbuf_r,
          es_0_2_1MyFalse_1_argbuf_r,
          \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ,
          lizzieLet17_4QNone_Int_2_argbuf_r} = (lizzieLet17_4QNone_Int_2_argbuf_done ? lizzieLet17_4QNone_Int_2_argbuf_select_d :
                                                5'd0);
  assign go_18_goMux_data_d = ((lizzieLet17_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_4QNone_Int_2_argbuf_d :
                               ((lizzieLet17_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d  :
                                ((lizzieLet17_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_2_1MyFalse_1_argbuf_d :
                                 ((lizzieLet17_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_2_1MyTrue_2_argbuf_d :
                                  ((lizzieLet17_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_4QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_18_goMux_choice_d = ((lizzieLet17_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet17_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet17_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet17_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet17_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet17_4QVal_Int,Go) > [(lizzieLet17_4QVal_Int_1,Go),
                                             (lizzieLet17_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet17_4QVal_Int_emitted;
  logic [1:0] lizzieLet17_4QVal_Int_done;
  assign lizzieLet17_4QVal_Int_1_d = (lizzieLet17_4QVal_Int_d[0] && (! lizzieLet17_4QVal_Int_emitted[0]));
  assign lizzieLet17_4QVal_Int_2_d = (lizzieLet17_4QVal_Int_d[0] && (! lizzieLet17_4QVal_Int_emitted[1]));
  assign lizzieLet17_4QVal_Int_done = (lizzieLet17_4QVal_Int_emitted | ({lizzieLet17_4QVal_Int_2_d[0],
                                                                         lizzieLet17_4QVal_Int_1_d[0]} & {lizzieLet17_4QVal_Int_2_r,
                                                                                                          lizzieLet17_4QVal_Int_1_r}));
  assign lizzieLet17_4QVal_Int_r = (& lizzieLet17_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet17_4QVal_Int_emitted <= (lizzieLet17_4QVal_Int_r ? 2'd0 :
                                        lizzieLet17_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_4QVal_Int_1,Go) > (lizzieLet17_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet17_4QVal_Int_1_bufchan_d;
  logic lizzieLet17_4QVal_Int_1_bufchan_r;
  assign lizzieLet17_4QVal_Int_1_r = ((! lizzieLet17_4QVal_Int_1_bufchan_d[0]) || lizzieLet17_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QVal_Int_1_r)
        lizzieLet17_4QVal_Int_1_bufchan_d <= lizzieLet17_4QVal_Int_1_d;
  Go_t lizzieLet17_4QVal_Int_1_bufchan_buf;
  assign lizzieLet17_4QVal_Int_1_bufchan_r = (! lizzieLet17_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_4QVal_Int_1_argbuf_d = (lizzieLet17_4QVal_Int_1_bufchan_buf[0] ? lizzieLet17_4QVal_Int_1_bufchan_buf :
                                             lizzieLet17_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QVal_Int_1_argbuf_r && lizzieLet17_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QVal_Int_1_argbuf_r) && (! lizzieLet17_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_4QVal_Int_1_bufchan_buf <= lizzieLet17_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet17_4QVal_Int_1_argbuf,Go),
                                          (lizzieLet17_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (xac0_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet17_4QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet17_5QVal_Int_1_argbuf_d[0],
                                                                                             xac0_1_argbuf_d[0]}), lizzieLet17_4QVal_Int_1_argbuf_d, lizzieLet17_5QVal_Int_1_argbuf_d, xac0_1_argbuf_d);
  assign {lizzieLet17_4QVal_Int_1_argbuf_r,
          lizzieLet17_5QVal_Int_1_argbuf_r,
          xac0_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_5,QTree_Int) (isZacC_goMux_mux,MyDTInt_Bool) > [(_22,MyDTInt_Bool),
                                                                                       (lizzieLet17_5QVal_Int,MyDTInt_Bool),
                                                                                       (lizzieLet17_5QNode_Int,MyDTInt_Bool),
                                                                                       (_21,MyDTInt_Bool)] */
  logic [3:0] isZacC_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_5_d[0] && isZacC_goMux_mux_d[0]))
      unique case (lizzieLet17_5_d[2:1])
        2'd0: isZacC_goMux_mux_onehotd = 4'd1;
        2'd1: isZacC_goMux_mux_onehotd = 4'd2;
        2'd2: isZacC_goMux_mux_onehotd = 4'd4;
        2'd3: isZacC_goMux_mux_onehotd = 4'd8;
        default: isZacC_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacC_goMux_mux_onehotd = 4'd0;
  assign _22_d = isZacC_goMux_mux_onehotd[0];
  assign lizzieLet17_5QVal_Int_d = isZacC_goMux_mux_onehotd[1];
  assign lizzieLet17_5QNode_Int_d = isZacC_goMux_mux_onehotd[2];
  assign _21_d = isZacC_goMux_mux_onehotd[3];
  assign isZacC_goMux_mux_r = (| (isZacC_goMux_mux_onehotd & {_21_r,
                                                              lizzieLet17_5QNode_Int_r,
                                                              lizzieLet17_5QVal_Int_r,
                                                              _22_r}));
  assign lizzieLet17_5_r = isZacC_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int,MyDTInt_Bool) > [(lizzieLet17_5QNode_Int_1,MyDTInt_Bool),
                                                                  (lizzieLet17_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet17_5QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_done;
  assign lizzieLet17_5QNode_Int_1_d = (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_2_d = (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_done = (lizzieLet17_5QNode_Int_emitted | ({lizzieLet17_5QNode_Int_2_d[0],
                                                                           lizzieLet17_5QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_2_r,
                                                                                                             lizzieLet17_5QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_r = (& lizzieLet17_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_emitted <= (lizzieLet17_5QNode_Int_r ? 2'd0 :
                                         lizzieLet17_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet17_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_2_r)
        lizzieLet17_5QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_5QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_2_bufchan_buf :
                                              lizzieLet17_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_5QVal_Int,MyDTInt_Bool) > (lizzieLet17_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_r = ((! lizzieLet17_5QVal_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_r)
        lizzieLet17_5QVal_Int_bufchan_d <= lizzieLet17_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet17_5QVal_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_bufchan_r = (! lizzieLet17_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_bufchan_buf :
                                             lizzieLet17_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_bufchan_buf <= lizzieLet17_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet17_6,QTree_Int) (sc_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) > [(lizzieLet17_6QNone_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                 (lizzieLet17_6QVal_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                 (lizzieLet17_6QNode_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                                 (lizzieLet17_6QError_Int,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [3:0] sc_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_6_d[0] && sc_0_3_goMux_mux_d[0]))
      unique case (lizzieLet17_6_d[2:1])
        2'd0: sc_0_3_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_3_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_3_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_3_goMux_mux_onehotd = 4'd8;
        default: sc_0_3_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_3_goMux_mux_onehotd = 4'd0;
  assign lizzieLet17_6QNone_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                     sc_0_3_goMux_mux_onehotd[0]};
  assign lizzieLet17_6QVal_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                    sc_0_3_goMux_mux_onehotd[1]};
  assign lizzieLet17_6QNode_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                     sc_0_3_goMux_mux_onehotd[2]};
  assign lizzieLet17_6QError_Int_d = {sc_0_3_goMux_mux_d[16:1],
                                      sc_0_3_goMux_mux_onehotd[3]};
  assign sc_0_3_goMux_mux_r = (| (sc_0_3_goMux_mux_onehotd & {lizzieLet17_6QError_Int_r,
                                                              lizzieLet17_6QNode_Int_r,
                                                              lizzieLet17_6QVal_Int_r,
                                                              lizzieLet17_6QNone_Int_r}));
  assign lizzieLet17_6_r = sc_0_3_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet17_6QError_Int,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet17_6QError_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QError_Int_bufchan_d;
  logic lizzieLet17_6QError_Int_bufchan_r;
  assign lizzieLet17_6QError_Int_r = ((! lizzieLet17_6QError_Int_bufchan_d[0]) || lizzieLet17_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_6QError_Int_r)
        lizzieLet17_6QError_Int_bufchan_d <= lizzieLet17_6QError_Int_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QError_Int_bufchan_buf;
  assign lizzieLet17_6QError_Int_bufchan_r = (! lizzieLet17_6QError_Int_bufchan_buf[0]);
  assign lizzieLet17_6QError_Int_1_argbuf_d = (lizzieLet17_6QError_Int_bufchan_buf[0] ? lizzieLet17_6QError_Int_bufchan_buf :
                                               lizzieLet17_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_6QError_Int_1_argbuf_r && lizzieLet17_6QError_Int_bufchan_buf[0]))
        lizzieLet17_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_6QError_Int_1_argbuf_r) && (! lizzieLet17_6QError_Int_bufchan_buf[0])))
        lizzieLet17_6QError_Int_bufchan_buf <= lizzieLet17_6QError_Int_bufchan_d;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int3) : [(lizzieLet17_6QNode_Int,Pointer_CTmap''_map''_Int_Int_Int),
                                              (lizzieLet17_5QNode_Int_1,MyDTInt_Bool),
                                              (lizzieLet17_3QNode_Int_1,MyDTInt_Int_Int),
                                              (lizzieLet17_7QNode_Int_1,Int),
                                              (q1acH_destruct,Pointer_QTree_Int),
                                              (q2acI_destruct,Pointer_QTree_Int),
                                              (q3acJ_destruct,Pointer_QTree_Int)] > (lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_d  = \Lcall_map''_map''_Int_Int_Int3_dc ((& {lizzieLet17_6QNode_Int_d[0],
                                                                                                                                                                                                           lizzieLet17_5QNode_Int_1_d[0],
                                                                                                                                                                                                           lizzieLet17_3QNode_Int_1_d[0],
                                                                                                                                                                                                           lizzieLet17_7QNode_Int_1_d[0],
                                                                                                                                                                                                           q1acH_destruct_d[0],
                                                                                                                                                                                                           q2acI_destruct_d[0],
                                                                                                                                                                                                           q3acJ_destruct_d[0]}), lizzieLet17_6QNode_Int_d, lizzieLet17_5QNode_Int_1_d, lizzieLet17_3QNode_Int_1_d, lizzieLet17_7QNode_Int_1_d, q1acH_destruct_d, q2acI_destruct_d, q3acJ_destruct_d);
  assign {lizzieLet17_6QNode_Int_r,
          lizzieLet17_5QNode_Int_1_r,
          lizzieLet17_3QNode_Int_1_r,
          lizzieLet17_7QNode_Int_1_r,
          q1acH_destruct_r,
          q2acI_destruct_r,
          q3acJ_destruct_r} = {7 {(\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_r  && \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) > (lizzieLet21_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_r  = ((! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d [0]) || \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= {99'd0,
                                                                                                                                                                          1'd0};
    else
      if (\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_r )
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_r  = (! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]);
  assign lizzieLet21_1_argbuf_d = (\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  :
                                   \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                            1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                              1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1lizzieLet17_7QNode_Int_1q1acH_1q2acI_1q3acJ_1Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (lizzieLet17_6QNone_Int,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet17_6QNone_Int_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QNone_Int_bufchan_d;
  logic lizzieLet17_6QNone_Int_bufchan_r;
  assign lizzieLet17_6QNone_Int_r = ((! lizzieLet17_6QNone_Int_bufchan_d[0]) || lizzieLet17_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_6QNone_Int_r)
        lizzieLet17_6QNone_Int_bufchan_d <= lizzieLet17_6QNone_Int_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  lizzieLet17_6QNone_Int_bufchan_buf;
  assign lizzieLet17_6QNone_Int_bufchan_r = (! lizzieLet17_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_6QNone_Int_1_argbuf_d = (lizzieLet17_6QNone_Int_bufchan_buf[0] ? lizzieLet17_6QNone_Int_bufchan_buf :
                                              lizzieLet17_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_6QNone_Int_1_argbuf_r && lizzieLet17_6QNone_Int_bufchan_buf[0]))
        lizzieLet17_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_6QNone_Int_1_argbuf_r) && (! lizzieLet17_6QNone_Int_bufchan_buf[0])))
        lizzieLet17_6QNone_Int_bufchan_buf <= lizzieLet17_6QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet17_7,QTree_Int) (v'acE_goMux_mux,Int) > [(_20,Int),
                                                                    (lizzieLet17_7QVal_Int,Int),
                                                                    (lizzieLet17_7QNode_Int,Int),
                                                                    (_19,Int)] */
  logic [3:0] \v'acE_goMux_mux_onehotd ;
  always_comb
    if ((lizzieLet17_7_d[0] && \v'acE_goMux_mux_d [0]))
      unique case (lizzieLet17_7_d[2:1])
        2'd0: \v'acE_goMux_mux_onehotd  = 4'd1;
        2'd1: \v'acE_goMux_mux_onehotd  = 4'd2;
        2'd2: \v'acE_goMux_mux_onehotd  = 4'd4;
        2'd3: \v'acE_goMux_mux_onehotd  = 4'd8;
        default: \v'acE_goMux_mux_onehotd  = 4'd0;
      endcase
    else \v'acE_goMux_mux_onehotd  = 4'd0;
  assign _20_d = {\v'acE_goMux_mux_d [32:1],
                  \v'acE_goMux_mux_onehotd [0]};
  assign lizzieLet17_7QVal_Int_d = {\v'acE_goMux_mux_d [32:1],
                                    \v'acE_goMux_mux_onehotd [1]};
  assign lizzieLet17_7QNode_Int_d = {\v'acE_goMux_mux_d [32:1],
                                     \v'acE_goMux_mux_onehotd [2]};
  assign _19_d = {\v'acE_goMux_mux_d [32:1],
                  \v'acE_goMux_mux_onehotd [3]};
  assign \v'acE_goMux_mux_r  = (| (\v'acE_goMux_mux_onehotd  & {_19_r,
                                                                lizzieLet17_7QNode_Int_r,
                                                                lizzieLet17_7QVal_Int_r,
                                                                _20_r}));
  assign lizzieLet17_7_r = \v'acE_goMux_mux_r ;
  
  /* fork (Ty Int) : (lizzieLet17_7QNode_Int,Int) > [(lizzieLet17_7QNode_Int_1,Int),
                                                (lizzieLet17_7QNode_Int_2,Int)] */
  logic [1:0] lizzieLet17_7QNode_Int_emitted;
  logic [1:0] lizzieLet17_7QNode_Int_done;
  assign lizzieLet17_7QNode_Int_1_d = {lizzieLet17_7QNode_Int_d[32:1],
                                       (lizzieLet17_7QNode_Int_d[0] && (! lizzieLet17_7QNode_Int_emitted[0]))};
  assign lizzieLet17_7QNode_Int_2_d = {lizzieLet17_7QNode_Int_d[32:1],
                                       (lizzieLet17_7QNode_Int_d[0] && (! lizzieLet17_7QNode_Int_emitted[1]))};
  assign lizzieLet17_7QNode_Int_done = (lizzieLet17_7QNode_Int_emitted | ({lizzieLet17_7QNode_Int_2_d[0],
                                                                           lizzieLet17_7QNode_Int_1_d[0]} & {lizzieLet17_7QNode_Int_2_r,
                                                                                                             lizzieLet17_7QNode_Int_1_r}));
  assign lizzieLet17_7QNode_Int_r = (& lizzieLet17_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_7QNode_Int_emitted <= (lizzieLet17_7QNode_Int_r ? 2'd0 :
                                         lizzieLet17_7QNode_Int_done);
  
  /* buf (Ty Int) : (lizzieLet17_7QNode_Int_2,Int) > (lizzieLet17_7QNode_Int_2_argbuf,Int) */
  Int_t lizzieLet17_7QNode_Int_2_bufchan_d;
  logic lizzieLet17_7QNode_Int_2_bufchan_r;
  assign lizzieLet17_7QNode_Int_2_r = ((! lizzieLet17_7QNode_Int_2_bufchan_d[0]) || lizzieLet17_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_7QNode_Int_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet17_7QNode_Int_2_r)
        lizzieLet17_7QNode_Int_2_bufchan_d <= lizzieLet17_7QNode_Int_2_d;
  Int_t lizzieLet17_7QNode_Int_2_bufchan_buf;
  assign lizzieLet17_7QNode_Int_2_bufchan_r = (! lizzieLet17_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_7QNode_Int_2_argbuf_d = (lizzieLet17_7QNode_Int_2_bufchan_buf[0] ? lizzieLet17_7QNode_Int_2_bufchan_buf :
                                              lizzieLet17_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_7QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet17_7QNode_Int_2_argbuf_r && lizzieLet17_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_7QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet17_7QNode_Int_2_argbuf_r) && (! lizzieLet17_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_7QNode_Int_2_bufchan_buf <= lizzieLet17_7QNode_Int_2_bufchan_d;
  
  /* buf (Ty Int) : (lizzieLet17_7QVal_Int,Int) > (lizzieLet17_7QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet17_7QVal_Int_bufchan_d;
  logic lizzieLet17_7QVal_Int_bufchan_r;
  assign lizzieLet17_7QVal_Int_r = ((! lizzieLet17_7QVal_Int_bufchan_d[0]) || lizzieLet17_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_7QVal_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet17_7QVal_Int_r)
        lizzieLet17_7QVal_Int_bufchan_d <= lizzieLet17_7QVal_Int_d;
  Int_t lizzieLet17_7QVal_Int_bufchan_buf;
  assign lizzieLet17_7QVal_Int_bufchan_r = (! lizzieLet17_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_7QVal_Int_1_argbuf_d = (lizzieLet17_7QVal_Int_bufchan_buf[0] ? lizzieLet17_7QVal_Int_bufchan_buf :
                                             lizzieLet17_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet17_7QVal_Int_1_argbuf_r && lizzieLet17_7QVal_Int_bufchan_buf[0]))
        lizzieLet17_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet17_7QVal_Int_1_argbuf_r) && (! lizzieLet17_7QVal_Int_bufchan_buf[0])))
        lizzieLet17_7QVal_Int_bufchan_buf <= lizzieLet17_7QVal_Int_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1X1j_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1X1j_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1X1j_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1X1j_1_Eq_r = ((! lizzieLet1_1wild1X1j_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1X1j_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X1j_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1X1j_1_Eq_r)
        lizzieLet1_1wild1X1j_1_Eq_bufchan_d <= lizzieLet1_1wild1X1j_1_Eq_d;
  Bool_t lizzieLet1_1wild1X1j_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1X1j_1_Eq_bufchan_r = (! lizzieLet1_1wild1X1j_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1X1j_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1X1j_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1X1j_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X1j_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1X1j_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1X1j_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1X1j_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1X1j_1_Eq_bufchan_buf <= lizzieLet1_1wild1X1j_1_Eq_bufchan_d;
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int0) : (lizzieLet26_1Lcall_$wnnz_Int0,CT$wnnz_Int) > [(wwsxo_4_destruct,Int#),
                                                                                  (ww1XyC_2_destruct,Int#),
                                                                                  (ww2XyF_1_destruct,Int#),
                                                                                  (sc_0_7_destruct,Pointer_CT$wnnz_Int)] */
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int0_emitted;
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int0_done;
  assign wwsxo_4_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int0_d[35:4],
                               (lizzieLet26_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int0_emitted[0]))};
  assign ww1XyC_2_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int0_d[67:36],
                                (lizzieLet26_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int0_emitted[1]))};
  assign ww2XyF_1_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int0_d[99:68],
                                (lizzieLet26_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int0_emitted[2]))};
  assign sc_0_7_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int0_d[115:100],
                              (lizzieLet26_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int0_emitted[3]))};
  assign lizzieLet26_1Lcall_$wnnz_Int0_done = (lizzieLet26_1Lcall_$wnnz_Int0_emitted | ({sc_0_7_destruct_d[0],
                                                                                         ww2XyF_1_destruct_d[0],
                                                                                         ww1XyC_2_destruct_d[0],
                                                                                         wwsxo_4_destruct_d[0]} & {sc_0_7_destruct_r,
                                                                                                                   ww2XyF_1_destruct_r,
                                                                                                                   ww1XyC_2_destruct_r,
                                                                                                                   wwsxo_4_destruct_r}));
  assign lizzieLet26_1Lcall_$wnnz_Int0_r = (& lizzieLet26_1Lcall_$wnnz_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet26_1Lcall_$wnnz_Int0_emitted <= 4'd0;
    else
      lizzieLet26_1Lcall_$wnnz_Int0_emitted <= (lizzieLet26_1Lcall_$wnnz_Int0_r ? 4'd0 :
                                                lizzieLet26_1Lcall_$wnnz_Int0_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int1) : (lizzieLet26_1Lcall_$wnnz_Int1,CT$wnnz_Int) > [(wwsxo_3_destruct,Int#),
                                                                                  (ww1XyC_1_destruct,Int#),
                                                                                  (sc_0_6_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4acY_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int1_emitted;
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int1_done;
  assign wwsxo_3_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int1_d[35:4],
                               (lizzieLet26_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int1_emitted[0]))};
  assign ww1XyC_1_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int1_d[67:36],
                                (lizzieLet26_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int1_emitted[1]))};
  assign sc_0_6_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int1_d[83:68],
                              (lizzieLet26_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int1_emitted[2]))};
  assign q4acY_3_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int1_d[99:84],
                               (lizzieLet26_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int1_emitted[3]))};
  assign lizzieLet26_1Lcall_$wnnz_Int1_done = (lizzieLet26_1Lcall_$wnnz_Int1_emitted | ({q4acY_3_destruct_d[0],
                                                                                         sc_0_6_destruct_d[0],
                                                                                         ww1XyC_1_destruct_d[0],
                                                                                         wwsxo_3_destruct_d[0]} & {q4acY_3_destruct_r,
                                                                                                                   sc_0_6_destruct_r,
                                                                                                                   ww1XyC_1_destruct_r,
                                                                                                                   wwsxo_3_destruct_r}));
  assign lizzieLet26_1Lcall_$wnnz_Int1_r = (& lizzieLet26_1Lcall_$wnnz_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet26_1Lcall_$wnnz_Int1_emitted <= 4'd0;
    else
      lizzieLet26_1Lcall_$wnnz_Int1_emitted <= (lizzieLet26_1Lcall_$wnnz_Int1_r ? 4'd0 :
                                                lizzieLet26_1Lcall_$wnnz_Int1_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int2) : (lizzieLet26_1Lcall_$wnnz_Int2,CT$wnnz_Int) > [(wwsxo_2_destruct,Int#),
                                                                                  (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4acY_2_destruct,Pointer_QTree_Int),
                                                                                  (q3acX_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int2_emitted;
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int2_done;
  assign wwsxo_2_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int2_d[35:4],
                               (lizzieLet26_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int2_emitted[0]))};
  assign sc_0_5_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int2_d[51:36],
                              (lizzieLet26_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int2_emitted[1]))};
  assign q4acY_2_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int2_d[67:52],
                               (lizzieLet26_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int2_emitted[2]))};
  assign q3acX_2_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int2_d[83:68],
                               (lizzieLet26_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int2_emitted[3]))};
  assign lizzieLet26_1Lcall_$wnnz_Int2_done = (lizzieLet26_1Lcall_$wnnz_Int2_emitted | ({q3acX_2_destruct_d[0],
                                                                                         q4acY_2_destruct_d[0],
                                                                                         sc_0_5_destruct_d[0],
                                                                                         wwsxo_2_destruct_d[0]} & {q3acX_2_destruct_r,
                                                                                                                   q4acY_2_destruct_r,
                                                                                                                   sc_0_5_destruct_r,
                                                                                                                   wwsxo_2_destruct_r}));
  assign lizzieLet26_1Lcall_$wnnz_Int2_r = (& lizzieLet26_1Lcall_$wnnz_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet26_1Lcall_$wnnz_Int2_emitted <= 4'd0;
    else
      lizzieLet26_1Lcall_$wnnz_Int2_emitted <= (lizzieLet26_1Lcall_$wnnz_Int2_r ? 4'd0 :
                                                lizzieLet26_1Lcall_$wnnz_Int2_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int3) : (lizzieLet26_1Lcall_$wnnz_Int3,CT$wnnz_Int) > [(sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4acY_1_destruct,Pointer_QTree_Int),
                                                                                  (q3acX_1_destruct,Pointer_QTree_Int),
                                                                                  (q2acW_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int3_emitted;
  logic [3:0] lizzieLet26_1Lcall_$wnnz_Int3_done;
  assign sc_0_4_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int3_d[19:4],
                              (lizzieLet26_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int3_emitted[0]))};
  assign q4acY_1_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int3_d[35:20],
                               (lizzieLet26_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int3_emitted[1]))};
  assign q3acX_1_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int3_d[51:36],
                               (lizzieLet26_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int3_emitted[2]))};
  assign q2acW_1_destruct_d = {lizzieLet26_1Lcall_$wnnz_Int3_d[67:52],
                               (lizzieLet26_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet26_1Lcall_$wnnz_Int3_emitted[3]))};
  assign lizzieLet26_1Lcall_$wnnz_Int3_done = (lizzieLet26_1Lcall_$wnnz_Int3_emitted | ({q2acW_1_destruct_d[0],
                                                                                         q3acX_1_destruct_d[0],
                                                                                         q4acY_1_destruct_d[0],
                                                                                         sc_0_4_destruct_d[0]} & {q2acW_1_destruct_r,
                                                                                                                  q3acX_1_destruct_r,
                                                                                                                  q4acY_1_destruct_r,
                                                                                                                  sc_0_4_destruct_r}));
  assign lizzieLet26_1Lcall_$wnnz_Int3_r = (& lizzieLet26_1Lcall_$wnnz_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet26_1Lcall_$wnnz_Int3_emitted <= 4'd0;
    else
      lizzieLet26_1Lcall_$wnnz_Int3_emitted <= (lizzieLet26_1Lcall_$wnnz_Int3_r ? 4'd0 :
                                                lizzieLet26_1Lcall_$wnnz_Int3_done);
  
  /* demux (Ty CT$wnnz_Int,
       Ty CT$wnnz_Int) : (lizzieLet26_2,CT$wnnz_Int) (lizzieLet26_1,CT$wnnz_Int) > [(_18,CT$wnnz_Int),
                                                                                    (lizzieLet26_1Lcall_$wnnz_Int3,CT$wnnz_Int),
                                                                                    (lizzieLet26_1Lcall_$wnnz_Int2,CT$wnnz_Int),
                                                                                    (lizzieLet26_1Lcall_$wnnz_Int1,CT$wnnz_Int),
                                                                                    (lizzieLet26_1Lcall_$wnnz_Int0,CT$wnnz_Int)] */
  logic [4:0] lizzieLet26_1_onehotd;
  always_comb
    if ((lizzieLet26_2_d[0] && lizzieLet26_1_d[0]))
      unique case (lizzieLet26_2_d[3:1])
        3'd0: lizzieLet26_1_onehotd = 5'd1;
        3'd1: lizzieLet26_1_onehotd = 5'd2;
        3'd2: lizzieLet26_1_onehotd = 5'd4;
        3'd3: lizzieLet26_1_onehotd = 5'd8;
        3'd4: lizzieLet26_1_onehotd = 5'd16;
        default: lizzieLet26_1_onehotd = 5'd0;
      endcase
    else lizzieLet26_1_onehotd = 5'd0;
  assign _18_d = {lizzieLet26_1_d[115:1], lizzieLet26_1_onehotd[0]};
  assign lizzieLet26_1Lcall_$wnnz_Int3_d = {lizzieLet26_1_d[115:1],
                                            lizzieLet26_1_onehotd[1]};
  assign lizzieLet26_1Lcall_$wnnz_Int2_d = {lizzieLet26_1_d[115:1],
                                            lizzieLet26_1_onehotd[2]};
  assign lizzieLet26_1Lcall_$wnnz_Int1_d = {lizzieLet26_1_d[115:1],
                                            lizzieLet26_1_onehotd[3]};
  assign lizzieLet26_1Lcall_$wnnz_Int0_d = {lizzieLet26_1_d[115:1],
                                            lizzieLet26_1_onehotd[4]};
  assign lizzieLet26_1_r = (| (lizzieLet26_1_onehotd & {lizzieLet26_1Lcall_$wnnz_Int0_r,
                                                        lizzieLet26_1Lcall_$wnnz_Int1_r,
                                                        lizzieLet26_1Lcall_$wnnz_Int2_r,
                                                        lizzieLet26_1Lcall_$wnnz_Int3_r,
                                                        _18_r}));
  assign lizzieLet26_2_r = lizzieLet26_1_r;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Go) : (lizzieLet26_3,CT$wnnz_Int) (go_15_goMux_data,Go) > [(_17,Go),
                                                                     (lizzieLet26_3Lcall_$wnnz_Int3,Go),
                                                                     (lizzieLet26_3Lcall_$wnnz_Int2,Go),
                                                                     (lizzieLet26_3Lcall_$wnnz_Int1,Go),
                                                                     (lizzieLet26_3Lcall_$wnnz_Int0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet26_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet26_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _17_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet26_3Lcall_$wnnz_Int3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet26_3Lcall_$wnnz_Int2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet26_3Lcall_$wnnz_Int1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet26_3Lcall_$wnnz_Int0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet26_3Lcall_$wnnz_Int0_r,
                                                              lizzieLet26_3Lcall_$wnnz_Int1_r,
                                                              lizzieLet26_3Lcall_$wnnz_Int2_r,
                                                              lizzieLet26_3Lcall_$wnnz_Int3_r,
                                                              _17_r}));
  assign lizzieLet26_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet26_3Lcall_$wnnz_Int0,Go) > (lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf,Go) */
  Go_t lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d;
  logic lizzieLet26_3Lcall_$wnnz_Int0_bufchan_r;
  assign lizzieLet26_3Lcall_$wnnz_Int0_r = ((! lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d[0]) || lizzieLet26_3Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet26_3Lcall_$wnnz_Int0_r)
        lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d <= lizzieLet26_3Lcall_$wnnz_Int0_d;
  Go_t lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf;
  assign lizzieLet26_3Lcall_$wnnz_Int0_bufchan_r = (! lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_d = (lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf[0] ? lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf :
                                                     lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_r && lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf[0]))
        lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_r) && (! lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf[0])))
        lizzieLet26_3Lcall_$wnnz_Int0_bufchan_buf <= lizzieLet26_3Lcall_$wnnz_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet26_3Lcall_$wnnz_Int1,Go) > (lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf,Go) */
  Go_t lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d;
  logic lizzieLet26_3Lcall_$wnnz_Int1_bufchan_r;
  assign lizzieLet26_3Lcall_$wnnz_Int1_r = ((! lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d[0]) || lizzieLet26_3Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet26_3Lcall_$wnnz_Int1_r)
        lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d <= lizzieLet26_3Lcall_$wnnz_Int1_d;
  Go_t lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf;
  assign lizzieLet26_3Lcall_$wnnz_Int1_bufchan_r = (! lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_d = (lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf[0] ? lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf :
                                                     lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_r && lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf[0]))
        lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet26_3Lcall_$wnnz_Int1_1_argbuf_r) && (! lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf[0])))
        lizzieLet26_3Lcall_$wnnz_Int1_bufchan_buf <= lizzieLet26_3Lcall_$wnnz_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet26_3Lcall_$wnnz_Int2,Go) > (lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf,Go) */
  Go_t lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet26_3Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet26_3Lcall_$wnnz_Int2_r = ((! lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet26_3Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet26_3Lcall_$wnnz_Int2_r)
        lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d <= lizzieLet26_3Lcall_$wnnz_Int2_d;
  Go_t lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet26_3Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_d = (lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf :
                                                     lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_r && lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet26_3Lcall_$wnnz_Int2_1_argbuf_r) && (! lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet26_3Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet26_3Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet26_3Lcall_$wnnz_Int3,Go) > (lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf,Go) */
  Go_t lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet26_3Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet26_3Lcall_$wnnz_Int3_r = ((! lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet26_3Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet26_3Lcall_$wnnz_Int3_r)
        lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d <= lizzieLet26_3Lcall_$wnnz_Int3_d;
  Go_t lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet26_3Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_d = (lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf :
                                                     lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_r && lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet26_3Lcall_$wnnz_Int3_1_argbuf_r) && (! lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet26_3Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet26_3Lcall_$wnnz_Int3_bufchan_d;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Int#) : (lizzieLet26_4,CT$wnnz_Int) (srtarg_0_goMux_mux,Int#) > [(lizzieLet26_4L$wnnz_Intsbos,Int#),
                                                                           (lizzieLet26_4Lcall_$wnnz_Int3,Int#),
                                                                           (lizzieLet26_4Lcall_$wnnz_Int2,Int#),
                                                                           (lizzieLet26_4Lcall_$wnnz_Int1,Int#),
                                                                           (lizzieLet26_4Lcall_$wnnz_Int0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet26_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet26_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet26_4L$wnnz_Intsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                          srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet26_4Lcall_$wnnz_Int3_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet26_4Lcall_$wnnz_Int2_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet26_4Lcall_$wnnz_Int1_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet26_4Lcall_$wnnz_Int0_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet26_4Lcall_$wnnz_Int0_r,
                                                                  lizzieLet26_4Lcall_$wnnz_Int1_r,
                                                                  lizzieLet26_4Lcall_$wnnz_Int2_r,
                                                                  lizzieLet26_4Lcall_$wnnz_Int3_r,
                                                                  lizzieLet26_4L$wnnz_Intsbos_r}));
  assign lizzieLet26_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet26_4L$wnnz_Intsbos,Int#) > [(lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#),
                                                       (lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet26_4L$wnnz_Intsbos_emitted;
  logic [1:0] lizzieLet26_4L$wnnz_Intsbos_done;
  assign lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_d = {lizzieLet26_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet26_4L$wnnz_Intsbos_d[0] && (! lizzieLet26_4L$wnnz_Intsbos_emitted[0]))};
  assign lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_d = {lizzieLet26_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet26_4L$wnnz_Intsbos_d[0] && (! lizzieLet26_4L$wnnz_Intsbos_emitted[1]))};
  assign lizzieLet26_4L$wnnz_Intsbos_done = (lizzieLet26_4L$wnnz_Intsbos_emitted | ({lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                     lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet26_4L$wnnz_Intsbos_r = (& lizzieLet26_4L$wnnz_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet26_4L$wnnz_Intsbos_emitted <= 2'd0;
    else
      lizzieLet26_4L$wnnz_Intsbos_emitted <= (lizzieLet26_4L$wnnz_Intsbos_r ? 2'd0 :
                                              lizzieLet26_4L$wnnz_Intsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_Int_goConst,Go) */
  assign call_$wnnz_Int_goConst_d = lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_1_r = call_$wnnz_Int_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#) > ($wnnz_Int_resbuf,Int#) */
  \Int#_t  lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                     1'd0};
    else
      if (lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_Int_resbuf_d  = (lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                       1'd0};
    else
      if ((\$wnnz_Int_resbuf_r  && lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                         1'd0};
      else if (((! \$wnnz_Int_resbuf_r ) && (! lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet26_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int2) : [(lizzieLet26_4Lcall_$wnnz_Int3,Int#),
                                (sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                (q4acY_1_destruct,Pointer_QTree_Int),
                                (q3acX_1_destruct,Pointer_QTree_Int)] > (lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) */
  assign lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_d = Lcall_$wnnz_Int2_dc((& {lizzieLet26_4Lcall_$wnnz_Int3_d[0],
                                                                                                               sc_0_4_destruct_d[0],
                                                                                                               q4acY_1_destruct_d[0],
                                                                                                               q3acX_1_destruct_d[0]}), lizzieLet26_4Lcall_$wnnz_Int3_d, sc_0_4_destruct_d, q4acY_1_destruct_d, q3acX_1_destruct_d);
  assign {lizzieLet26_4Lcall_$wnnz_Int3_r,
          sc_0_4_destruct_r,
          q4acY_1_destruct_r,
          q3acX_1_destruct_r} = {4 {(lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_r && lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) > (lizzieLet27_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_r = ((! lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_r)
        lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d <= lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_d;
  CT$wnnz_Int_t lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf :
                                   lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet26_4Lcall_$wnnz_Int3_1sc_0_4_1q4acY_1_1q3acX_1_1Lcall_$wnnz_Int2_bufchan_d;
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int0) : (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) > [(es_1_1_destruct,Pointer_QTree_Int),
                                                                                                                      (es_2_1_destruct,Pointer_QTree_Int),
                                                                                                                      (es_3_3_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_11_destruct,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [3:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted;
  logic [3:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_done;
  assign es_1_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[19:4],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted[0]))};
  assign es_2_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[35:20],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted[1]))};
  assign es_3_3_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[51:36],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted[2]))};
  assign sc_0_11_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[67:52],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted[3]))};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_done = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted | ({sc_0_11_destruct_d[0],
                                                                                                                 es_3_3_destruct_d[0],
                                                                                                                 es_2_1_destruct_d[0],
                                                                                                                 es_1_1_destruct_d[0]} & {sc_0_11_destruct_r,
                                                                                                                                          es_3_3_destruct_r,
                                                                                                                                          es_2_1_destruct_r,
                                                                                                                                          es_1_1_destruct_r}));
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_r = (& lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted <= 4'd0;
    else
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_emitted <= (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_r ? 4'd0 :
                                                            lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int1) : (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) > [(es_2_destruct,Pointer_QTree_Int),
                                                                                                                      (es_3_2_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_10_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZacL_4_destruct,MyDTInt_Bool),
                                                                                                                      (gacM_4_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1acQ_3_destruct,Pointer_QTree_Int),
                                                                                                                      (m2acO_4_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted;
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_done;
  assign es_2_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[19:4],
                            (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[35:20],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[1]))};
  assign sc_0_10_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[51:36],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[2]))};
  assign isZacL_4_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[3]));
  assign gacM_4_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[4]));
  assign q1acQ_3_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[67:52],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[5]))};
  assign m2acO_4_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[83:68],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted[6]))};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_done = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted | ({m2acO_4_destruct_d[0],
                                                                                                                 q1acQ_3_destruct_d[0],
                                                                                                                 gacM_4_destruct_d[0],
                                                                                                                 isZacL_4_destruct_d[0],
                                                                                                                 sc_0_10_destruct_d[0],
                                                                                                                 es_3_2_destruct_d[0],
                                                                                                                 es_2_destruct_d[0]} & {m2acO_4_destruct_r,
                                                                                                                                        q1acQ_3_destruct_r,
                                                                                                                                        gacM_4_destruct_r,
                                                                                                                                        isZacL_4_destruct_r,
                                                                                                                                        sc_0_10_destruct_r,
                                                                                                                                        es_3_2_destruct_r,
                                                                                                                                        es_2_destruct_r}));
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_r = (& lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted <= 7'd0;
    else
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_emitted <= (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_r ? 7'd0 :
                                                            lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int2) : (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) > [(es_3_1_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_9_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZacL_3_destruct,MyDTInt_Bool),
                                                                                                                      (gacM_3_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1acQ_2_destruct,Pointer_QTree_Int),
                                                                                                                      (m2acO_3_destruct,Pointer_QTree_Int),
                                                                                                                      (q2acR_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted;
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_done;
  assign es_3_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[19:4],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[0]))};
  assign sc_0_9_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[35:20],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[1]))};
  assign isZacL_3_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[2]));
  assign gacM_3_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[3]));
  assign q1acQ_2_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[51:36],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[4]))};
  assign m2acO_3_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[67:52],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[5]))};
  assign q2acR_2_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[83:68],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted[6]))};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_done = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted | ({q2acR_2_destruct_d[0],
                                                                                                                 m2acO_3_destruct_d[0],
                                                                                                                 q1acQ_2_destruct_d[0],
                                                                                                                 gacM_3_destruct_d[0],
                                                                                                                 isZacL_3_destruct_d[0],
                                                                                                                 sc_0_9_destruct_d[0],
                                                                                                                 es_3_1_destruct_d[0]} & {q2acR_2_destruct_r,
                                                                                                                                          m2acO_3_destruct_r,
                                                                                                                                          q1acQ_2_destruct_r,
                                                                                                                                          gacM_3_destruct_r,
                                                                                                                                          isZacL_3_destruct_r,
                                                                                                                                          sc_0_9_destruct_r,
                                                                                                                                          es_3_1_destruct_r}));
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_r = (& lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted <= 7'd0;
    else
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_emitted <= (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_r ? 7'd0 :
                                                            lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_done);
  
  /* destruct (Ty CTkron_kron_Int_Int_Int,
          Dcon Lcall_kron_kron_Int_Int_Int3) : (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) > [(sc_0_8_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                      (isZacL_2_destruct,MyDTInt_Bool),
                                                                                                                      (gacM_2_destruct,MyDTInt_Int_Int),
                                                                                                                      (q1acQ_1_destruct,Pointer_QTree_Int),
                                                                                                                      (m2acO_2_destruct,Pointer_QTree_Int),
                                                                                                                      (q2acR_1_destruct,Pointer_QTree_Int),
                                                                                                                      (q3acS_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted;
  logic [6:0] lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_done;
  assign sc_0_8_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[19:4],
                              (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[0]))};
  assign isZacL_2_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[1]));
  assign gacM_2_destruct_d = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[2]));
  assign q1acQ_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[35:20],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[3]))};
  assign m2acO_2_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[51:36],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[4]))};
  assign q2acR_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[67:52],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[5]))};
  assign q3acS_1_destruct_d = {lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[83:68],
                               (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d[0] && (! lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted[6]))};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_done = (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted | ({q3acS_1_destruct_d[0],
                                                                                                                 q2acR_1_destruct_d[0],
                                                                                                                 m2acO_2_destruct_d[0],
                                                                                                                 q1acQ_1_destruct_d[0],
                                                                                                                 gacM_2_destruct_d[0],
                                                                                                                 isZacL_2_destruct_d[0],
                                                                                                                 sc_0_8_destruct_d[0]} & {q3acS_1_destruct_r,
                                                                                                                                          q2acR_1_destruct_r,
                                                                                                                                          m2acO_2_destruct_r,
                                                                                                                                          q1acQ_1_destruct_r,
                                                                                                                                          gacM_2_destruct_r,
                                                                                                                                          isZacL_2_destruct_r,
                                                                                                                                          sc_0_8_destruct_r}));
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_r = (& lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted <= 7'd0;
    else
      lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_emitted <= (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_r ? 7'd0 :
                                                            lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_done);
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty CTkron_kron_Int_Int_Int) : (lizzieLet30_2,CTkron_kron_Int_Int_Int) (lizzieLet30_1,CTkron_kron_Int_Int_Int) > [(_16,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet30_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet30_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet30_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int),
                                                                                                                        (lizzieLet30_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int)] */
  logic [4:0] lizzieLet30_1_onehotd;
  always_comb
    if ((lizzieLet30_2_d[0] && lizzieLet30_1_d[0]))
      unique case (lizzieLet30_2_d[3:1])
        3'd0: lizzieLet30_1_onehotd = 5'd1;
        3'd1: lizzieLet30_1_onehotd = 5'd2;
        3'd2: lizzieLet30_1_onehotd = 5'd4;
        3'd3: lizzieLet30_1_onehotd = 5'd8;
        3'd4: lizzieLet30_1_onehotd = 5'd16;
        default: lizzieLet30_1_onehotd = 5'd0;
      endcase
    else lizzieLet30_1_onehotd = 5'd0;
  assign _16_d = {lizzieLet30_1_d[83:1], lizzieLet30_1_onehotd[0]};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_d = {lizzieLet30_1_d[83:1],
                                                        lizzieLet30_1_onehotd[1]};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_d = {lizzieLet30_1_d[83:1],
                                                        lizzieLet30_1_onehotd[2]};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_d = {lizzieLet30_1_d[83:1],
                                                        lizzieLet30_1_onehotd[3]};
  assign lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_d = {lizzieLet30_1_d[83:1],
                                                        lizzieLet30_1_onehotd[4]};
  assign lizzieLet30_1_r = (| (lizzieLet30_1_onehotd & {lizzieLet30_1Lcall_kron_kron_Int_Int_Int0_r,
                                                        lizzieLet30_1Lcall_kron_kron_Int_Int_Int1_r,
                                                        lizzieLet30_1Lcall_kron_kron_Int_Int_Int2_r,
                                                        lizzieLet30_1Lcall_kron_kron_Int_Int_Int3_r,
                                                        _16_r}));
  assign lizzieLet30_2_r = lizzieLet30_1_r;
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty Go) : (lizzieLet30_3,CTkron_kron_Int_Int_Int) (go_16_goMux_data,Go) > [(_15,Go),
                                                                                 (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3,Go),
                                                                                 (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2,Go),
                                                                                 (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1,Go),
                                                                                 (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0,Go)] */
  logic [4:0] go_16_goMux_data_onehotd;
  always_comb
    if ((lizzieLet30_3_d[0] && go_16_goMux_data_d[0]))
      unique case (lizzieLet30_3_d[3:1])
        3'd0: go_16_goMux_data_onehotd = 5'd1;
        3'd1: go_16_goMux_data_onehotd = 5'd2;
        3'd2: go_16_goMux_data_onehotd = 5'd4;
        3'd3: go_16_goMux_data_onehotd = 5'd8;
        3'd4: go_16_goMux_data_onehotd = 5'd16;
        default: go_16_goMux_data_onehotd = 5'd0;
      endcase
    else go_16_goMux_data_onehotd = 5'd0;
  assign _15_d = go_16_goMux_data_onehotd[0];
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_d = go_16_goMux_data_onehotd[1];
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_d = go_16_goMux_data_onehotd[2];
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_d = go_16_goMux_data_onehotd[3];
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_d = go_16_goMux_data_onehotd[4];
  assign go_16_goMux_data_r = (| (go_16_goMux_data_onehotd & {lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_r,
                                                              lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_r,
                                                              lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_r,
                                                              lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_r,
                                                              _15_r}));
  assign lizzieLet30_3_r = go_16_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0,Go) > (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf,Go) */
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_r;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_r = ((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d[0]) || lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_r)
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_d;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_r = (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d = (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0] ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf :
                                                                 lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r && lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r) && (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1,Go) > (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf,Go) */
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_r;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_r = ((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d[0]) || lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_r)
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_d;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_r = (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_d = (lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0] ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf :
                                                                 lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r && lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_1_argbuf_r) && (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2,Go) > (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf,Go) */
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_r;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_r = ((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d[0]) || lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_r)
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_d;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_r = (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_d = (lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0] ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf :
                                                                 lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r && lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_1_argbuf_r) && (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3,Go) > (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf,Go) */
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  logic lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_r;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_r = ((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d[0]) || lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_r)
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_d;
  Go_t lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf;
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_r = (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_d = (lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0] ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf :
                                                                 lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r && lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_1_argbuf_r) && (! lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= lizzieLet30_3Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  
  /* demux (Ty CTkron_kron_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet30_4,CTkron_kron_Int_Int_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet30_4Lkron_kron_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                   (lizzieLet30_4Lcall_kron_kron_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                   (lizzieLet30_4Lcall_kron_kron_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                   (lizzieLet30_4Lcall_kron_kron_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                   (lizzieLet30_4Lcall_kron_kron_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet30_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet30_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                      srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_r,
                                                                      lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_r,
                                                                      lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_r,
                                                                      lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_r,
                                                                      lizzieLet30_4Lkron_kron_Int_Int_Intsbos_r}));
  assign lizzieLet30_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet30_4Lcall_kron_kron_Int_Int_Int0,Pointer_QTree_Int),
                         (es_1_1_destruct,Pointer_QTree_Int),
                         (es_2_1_destruct,Pointer_QTree_Int),
                         (es_3_3_destruct,Pointer_QTree_Int)] > (lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int,QTree_Int) */
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_d = QNode_Int_dc((& {lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_d[0],
                                                                                                           es_1_1_destruct_d[0],
                                                                                                           es_2_1_destruct_d[0],
                                                                                                           es_3_3_destruct_d[0]}), lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_d, es_1_1_destruct_d, es_2_1_destruct_d, es_3_3_destruct_d);
  assign {lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_r,
          es_1_1_destruct_r,
          es_2_1_destruct_r,
          es_3_3_destruct_r} = {4 {(lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int,QTree_Int) > (lizzieLet34_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_r;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_r = ((! lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d[0]) || lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d <= {66'd0,
                                                                                                 1'd0};
    else
      if (lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_r)
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_d;
  QTree_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_r = (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf[0] ? lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf :
                                   lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf[0]))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf[0])))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_buf <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int0_1es_1_1_1es_2_1_1es_3_3_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int0) : [(lizzieLet30_4Lcall_kron_kron_Int_Int_Int1,Pointer_QTree_Int),
                                            (es_2_destruct,Pointer_QTree_Int),
                                            (es_3_2_destruct,Pointer_QTree_Int),
                                            (sc_0_10_destruct,Pointer_CTkron_kron_Int_Int_Int)] > (lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) */
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d = Lcall_kron_kron_Int_Int_Int0_dc((& {lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_d[0],
                                                                                                                                                es_2_destruct_d[0],
                                                                                                                                                es_3_2_destruct_d[0],
                                                                                                                                                sc_0_10_destruct_d[0]}), lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_d, es_2_destruct_d, es_3_2_destruct_d, sc_0_10_destruct_d);
  assign {lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_r,
          es_2_destruct_r,
          es_3_2_destruct_r,
          sc_0_10_destruct_r} = {4 {(lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0,CTkron_kron_Int_Int_Int) > (lizzieLet33_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r = ((! lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d[0]) || lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d <= {83'd0,
                                                                                                                   1'd0};
    else
      if (lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_r)
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_d;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_r = (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0] ? lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf :
                                   lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                     1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                       1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_buf <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int1_1es_2_1es_3_2_1sc_0_10_1Lcall_kron_kron_Int_Int_Int0_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int1) : [(lizzieLet30_4Lcall_kron_kron_Int_Int_Int2,Pointer_QTree_Int),
                                            (es_3_1_destruct,Pointer_QTree_Int),
                                            (sc_0_9_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                            (isZacL_3_1,MyDTInt_Bool),
                                            (gacM_3_1,MyDTInt_Int_Int),
                                            (q1acQ_2_destruct,Pointer_QTree_Int),
                                            (m2acO_3_1,Pointer_QTree_Int)] > (lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) */
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_d = Lcall_kron_kron_Int_Int_Int1_dc((& {lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_d[0],
                                                                                                                                                                             es_3_1_destruct_d[0],
                                                                                                                                                                             sc_0_9_destruct_d[0],
                                                                                                                                                                             isZacL_3_1_d[0],
                                                                                                                                                                             gacM_3_1_d[0],
                                                                                                                                                                             q1acQ_2_destruct_d[0],
                                                                                                                                                                             m2acO_3_1_d[0]}), lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_d, es_3_1_destruct_d, sc_0_9_destruct_d, isZacL_3_1_d, gacM_3_1_d, q1acQ_2_destruct_d, m2acO_3_1_d);
  assign {lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_r,
          es_3_1_destruct_r,
          sc_0_9_destruct_r,
          isZacL_3_1_r,
          gacM_3_1_r,
          q1acQ_2_destruct_r,
          m2acO_3_1_r} = {7 {(lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1,CTkron_kron_Int_Int_Int) > (lizzieLet32_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_r = ((! lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d[0]) || lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d <= {83'd0,
                                                                                                                                                1'd0};
    else
      if (lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_r)
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_d;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_r = (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0] ? lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf :
                                   lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                  1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                    1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_buf <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int2_1es_3_1_1sc_0_9_1isZacL_3_1gacM_3_1q1acQ_2_1m2acO_3_1Lcall_kron_kron_Int_Int_Int1_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int2) : [(lizzieLet30_4Lcall_kron_kron_Int_Int_Int3,Pointer_QTree_Int),
                                            (sc_0_8_destruct,Pointer_CTkron_kron_Int_Int_Int),
                                            (isZacL_2_1,MyDTInt_Bool),
                                            (gacM_2_1,MyDTInt_Int_Int),
                                            (q1acQ_1_destruct,Pointer_QTree_Int),
                                            (m2acO_2_1,Pointer_QTree_Int),
                                            (q2acR_1_destruct,Pointer_QTree_Int)] > (lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) */
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_d = Lcall_kron_kron_Int_Int_Int2_dc((& {lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_d[0],
                                                                                                                                                                              sc_0_8_destruct_d[0],
                                                                                                                                                                              isZacL_2_1_d[0],
                                                                                                                                                                              gacM_2_1_d[0],
                                                                                                                                                                              q1acQ_1_destruct_d[0],
                                                                                                                                                                              m2acO_2_1_d[0],
                                                                                                                                                                              q2acR_1_destruct_d[0]}), lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_d, sc_0_8_destruct_d, isZacL_2_1_d, gacM_2_1_d, q1acQ_1_destruct_d, m2acO_2_1_d, q2acR_1_destruct_d);
  assign {lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_r,
          sc_0_8_destruct_r,
          isZacL_2_1_r,
          gacM_2_1_r,
          q1acQ_1_destruct_r,
          m2acO_2_1_r,
          q2acR_1_destruct_r} = {7 {(lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2,CTkron_kron_Int_Int_Int) > (lizzieLet31_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  logic lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_r = ((! lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d[0]) || lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d <= {83'd0,
                                                                                                                                                 1'd0};
    else
      if (lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_r)
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_d;
  CTkron_kron_Int_Int_Int_t lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf;
  assign lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_r = (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0] ? lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf :
                                   lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                   1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                     1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_buf <= lizzieLet30_4Lcall_kron_kron_Int_Int_Int3_1sc_0_8_1isZacL_2_1gacM_2_1q1acQ_1_1m2acO_2_1q2acR_1_1Lcall_kron_kron_Int_Int_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet30_4Lkron_kron_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                             (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted;
  logic [1:0] lizzieLet30_4Lkron_kron_Int_Int_Intsbos_done;
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d = {lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d[16:1],
                                                                           (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d[0] && (! lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted[0]))};
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d = {lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d[16:1],
                                                                           (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_d[0] && (! lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted[1]))};
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_done = (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted | ({lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                                             lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                                                   lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_r = (& lizzieLet30_4Lkron_kron_Int_Int_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted <= 2'd0;
    else
      lizzieLet30_4Lkron_kron_Int_Int_Intsbos_emitted <= (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_r ? 2'd0 :
                                                          lizzieLet30_4Lkron_kron_Int_Int_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_kron_kron_Int_Int_Int_goConst,Go) */
  assign call_kron_kron_Int_Int_Int_goConst_d = lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_1_r = call_kron_kron_Int_Int_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (kron_kron_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                                 1'd0};
    else
      if (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign kron_kron_Int_Int_Int_resbuf_d = (lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                           lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                   1'd0};
    else
      if ((kron_kron_Int_Int_Int_resbuf_r && lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                     1'd0};
      else if (((! kron_kron_Int_Int_Int_resbuf_r) && (! lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet30_4Lkron_kron_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int0) : (lizzieLet35_1Lcall_main_mask_Int0,CTmain_mask_Int) > [(es_1_2_destruct,Pointer_QTree_Int),
                                                                                              (es_2_3_destruct,Pointer_QTree_Int),
                                                                                              (es_3_6_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_15_destruct,Pointer_CTmain_mask_Int)] */
  logic [3:0] lizzieLet35_1Lcall_main_mask_Int0_emitted;
  logic [3:0] lizzieLet35_1Lcall_main_mask_Int0_done;
  assign es_1_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int0_d[19:4],
                              (lizzieLet35_1Lcall_main_mask_Int0_d[0] && (! lizzieLet35_1Lcall_main_mask_Int0_emitted[0]))};
  assign es_2_3_destruct_d = {lizzieLet35_1Lcall_main_mask_Int0_d[35:20],
                              (lizzieLet35_1Lcall_main_mask_Int0_d[0] && (! lizzieLet35_1Lcall_main_mask_Int0_emitted[1]))};
  assign es_3_6_destruct_d = {lizzieLet35_1Lcall_main_mask_Int0_d[51:36],
                              (lizzieLet35_1Lcall_main_mask_Int0_d[0] && (! lizzieLet35_1Lcall_main_mask_Int0_emitted[2]))};
  assign sc_0_15_destruct_d = {lizzieLet35_1Lcall_main_mask_Int0_d[67:52],
                               (lizzieLet35_1Lcall_main_mask_Int0_d[0] && (! lizzieLet35_1Lcall_main_mask_Int0_emitted[3]))};
  assign lizzieLet35_1Lcall_main_mask_Int0_done = (lizzieLet35_1Lcall_main_mask_Int0_emitted | ({sc_0_15_destruct_d[0],
                                                                                                 es_3_6_destruct_d[0],
                                                                                                 es_2_3_destruct_d[0],
                                                                                                 es_1_2_destruct_d[0]} & {sc_0_15_destruct_r,
                                                                                                                          es_3_6_destruct_r,
                                                                                                                          es_2_3_destruct_r,
                                                                                                                          es_1_2_destruct_r}));
  assign lizzieLet35_1Lcall_main_mask_Int0_r = (& lizzieLet35_1Lcall_main_mask_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_1Lcall_main_mask_Int0_emitted <= 4'd0;
    else
      lizzieLet35_1Lcall_main_mask_Int0_emitted <= (lizzieLet35_1Lcall_main_mask_Int0_r ? 4'd0 :
                                                    lizzieLet35_1Lcall_main_mask_Int0_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int1) : (lizzieLet35_1Lcall_main_mask_Int1,CTmain_mask_Int) > [(es_2_2_destruct,Pointer_QTree_Int),
                                                                                              (es_3_5_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_14_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1acr_3_destruct,Pointer_QTree_Int),
                                                                                              (q1acm_3_destruct,Pointer_MaskQTree)] */
  logic [4:0] lizzieLet35_1Lcall_main_mask_Int1_emitted;
  logic [4:0] lizzieLet35_1Lcall_main_mask_Int1_done;
  assign es_2_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int1_d[19:4],
                              (lizzieLet35_1Lcall_main_mask_Int1_d[0] && (! lizzieLet35_1Lcall_main_mask_Int1_emitted[0]))};
  assign es_3_5_destruct_d = {lizzieLet35_1Lcall_main_mask_Int1_d[35:20],
                              (lizzieLet35_1Lcall_main_mask_Int1_d[0] && (! lizzieLet35_1Lcall_main_mask_Int1_emitted[1]))};
  assign sc_0_14_destruct_d = {lizzieLet35_1Lcall_main_mask_Int1_d[51:36],
                               (lizzieLet35_1Lcall_main_mask_Int1_d[0] && (! lizzieLet35_1Lcall_main_mask_Int1_emitted[2]))};
  assign t1acr_3_destruct_d = {lizzieLet35_1Lcall_main_mask_Int1_d[67:52],
                               (lizzieLet35_1Lcall_main_mask_Int1_d[0] && (! lizzieLet35_1Lcall_main_mask_Int1_emitted[3]))};
  assign q1acm_3_destruct_d = {lizzieLet35_1Lcall_main_mask_Int1_d[83:68],
                               (lizzieLet35_1Lcall_main_mask_Int1_d[0] && (! lizzieLet35_1Lcall_main_mask_Int1_emitted[4]))};
  assign lizzieLet35_1Lcall_main_mask_Int1_done = (lizzieLet35_1Lcall_main_mask_Int1_emitted | ({q1acm_3_destruct_d[0],
                                                                                                 t1acr_3_destruct_d[0],
                                                                                                 sc_0_14_destruct_d[0],
                                                                                                 es_3_5_destruct_d[0],
                                                                                                 es_2_2_destruct_d[0]} & {q1acm_3_destruct_r,
                                                                                                                          t1acr_3_destruct_r,
                                                                                                                          sc_0_14_destruct_r,
                                                                                                                          es_3_5_destruct_r,
                                                                                                                          es_2_2_destruct_r}));
  assign lizzieLet35_1Lcall_main_mask_Int1_r = (& lizzieLet35_1Lcall_main_mask_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_1Lcall_main_mask_Int1_emitted <= 5'd0;
    else
      lizzieLet35_1Lcall_main_mask_Int1_emitted <= (lizzieLet35_1Lcall_main_mask_Int1_r ? 5'd0 :
                                                    lizzieLet35_1Lcall_main_mask_Int1_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int2) : (lizzieLet35_1Lcall_main_mask_Int2,CTmain_mask_Int) > [(es_3_4_destruct,Pointer_QTree_Int),
                                                                                              (sc_0_13_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1acr_2_destruct,Pointer_QTree_Int),
                                                                                              (q1acm_2_destruct,Pointer_MaskQTree),
                                                                                              (t2acs_2_destruct,Pointer_QTree_Int),
                                                                                              (q2acn_2_destruct,Pointer_MaskQTree)] */
  logic [5:0] lizzieLet35_1Lcall_main_mask_Int2_emitted;
  logic [5:0] lizzieLet35_1Lcall_main_mask_Int2_done;
  assign es_3_4_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[19:4],
                              (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[0]))};
  assign sc_0_13_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[35:20],
                               (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[1]))};
  assign t1acr_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[51:36],
                               (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[2]))};
  assign q1acm_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[67:52],
                               (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[3]))};
  assign t2acs_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[83:68],
                               (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[4]))};
  assign q2acn_2_destruct_d = {lizzieLet35_1Lcall_main_mask_Int2_d[99:84],
                               (lizzieLet35_1Lcall_main_mask_Int2_d[0] && (! lizzieLet35_1Lcall_main_mask_Int2_emitted[5]))};
  assign lizzieLet35_1Lcall_main_mask_Int2_done = (lizzieLet35_1Lcall_main_mask_Int2_emitted | ({q2acn_2_destruct_d[0],
                                                                                                 t2acs_2_destruct_d[0],
                                                                                                 q1acm_2_destruct_d[0],
                                                                                                 t1acr_2_destruct_d[0],
                                                                                                 sc_0_13_destruct_d[0],
                                                                                                 es_3_4_destruct_d[0]} & {q2acn_2_destruct_r,
                                                                                                                          t2acs_2_destruct_r,
                                                                                                                          q1acm_2_destruct_r,
                                                                                                                          t1acr_2_destruct_r,
                                                                                                                          sc_0_13_destruct_r,
                                                                                                                          es_3_4_destruct_r}));
  assign lizzieLet35_1Lcall_main_mask_Int2_r = (& lizzieLet35_1Lcall_main_mask_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_1Lcall_main_mask_Int2_emitted <= 6'd0;
    else
      lizzieLet35_1Lcall_main_mask_Int2_emitted <= (lizzieLet35_1Lcall_main_mask_Int2_r ? 6'd0 :
                                                    lizzieLet35_1Lcall_main_mask_Int2_done);
  
  /* destruct (Ty CTmain_mask_Int,
          Dcon Lcall_main_mask_Int3) : (lizzieLet35_1Lcall_main_mask_Int3,CTmain_mask_Int) > [(sc_0_12_destruct,Pointer_CTmain_mask_Int),
                                                                                              (t1acr_1_destruct,Pointer_QTree_Int),
                                                                                              (q1acm_1_destruct,Pointer_MaskQTree),
                                                                                              (t2acs_1_destruct,Pointer_QTree_Int),
                                                                                              (q2acn_1_destruct,Pointer_MaskQTree),
                                                                                              (t3act_1_destruct,Pointer_QTree_Int),
                                                                                              (q3aco_1_destruct,Pointer_MaskQTree)] */
  logic [6:0] lizzieLet35_1Lcall_main_mask_Int3_emitted;
  logic [6:0] lizzieLet35_1Lcall_main_mask_Int3_done;
  assign sc_0_12_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[19:4],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[0]))};
  assign t1acr_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[35:20],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[1]))};
  assign q1acm_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[51:36],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[2]))};
  assign t2acs_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[67:52],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[3]))};
  assign q2acn_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[83:68],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[4]))};
  assign t3act_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[99:84],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[5]))};
  assign q3aco_1_destruct_d = {lizzieLet35_1Lcall_main_mask_Int3_d[115:100],
                               (lizzieLet35_1Lcall_main_mask_Int3_d[0] && (! lizzieLet35_1Lcall_main_mask_Int3_emitted[6]))};
  assign lizzieLet35_1Lcall_main_mask_Int3_done = (lizzieLet35_1Lcall_main_mask_Int3_emitted | ({q3aco_1_destruct_d[0],
                                                                                                 t3act_1_destruct_d[0],
                                                                                                 q2acn_1_destruct_d[0],
                                                                                                 t2acs_1_destruct_d[0],
                                                                                                 q1acm_1_destruct_d[0],
                                                                                                 t1acr_1_destruct_d[0],
                                                                                                 sc_0_12_destruct_d[0]} & {q3aco_1_destruct_r,
                                                                                                                           t3act_1_destruct_r,
                                                                                                                           q2acn_1_destruct_r,
                                                                                                                           t2acs_1_destruct_r,
                                                                                                                           q1acm_1_destruct_r,
                                                                                                                           t1acr_1_destruct_r,
                                                                                                                           sc_0_12_destruct_r}));
  assign lizzieLet35_1Lcall_main_mask_Int3_r = (& lizzieLet35_1Lcall_main_mask_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_1Lcall_main_mask_Int3_emitted <= 7'd0;
    else
      lizzieLet35_1Lcall_main_mask_Int3_emitted <= (lizzieLet35_1Lcall_main_mask_Int3_r ? 7'd0 :
                                                    lizzieLet35_1Lcall_main_mask_Int3_done);
  
  /* demux (Ty CTmain_mask_Int,
       Ty CTmain_mask_Int) : (lizzieLet35_2,CTmain_mask_Int) (lizzieLet35_1,CTmain_mask_Int) > [(_14,CTmain_mask_Int),
                                                                                                (lizzieLet35_1Lcall_main_mask_Int3,CTmain_mask_Int),
                                                                                                (lizzieLet35_1Lcall_main_mask_Int2,CTmain_mask_Int),
                                                                                                (lizzieLet35_1Lcall_main_mask_Int1,CTmain_mask_Int),
                                                                                                (lizzieLet35_1Lcall_main_mask_Int0,CTmain_mask_Int)] */
  logic [4:0] lizzieLet35_1_onehotd;
  always_comb
    if ((lizzieLet35_2_d[0] && lizzieLet35_1_d[0]))
      unique case (lizzieLet35_2_d[3:1])
        3'd0: lizzieLet35_1_onehotd = 5'd1;
        3'd1: lizzieLet35_1_onehotd = 5'd2;
        3'd2: lizzieLet35_1_onehotd = 5'd4;
        3'd3: lizzieLet35_1_onehotd = 5'd8;
        3'd4: lizzieLet35_1_onehotd = 5'd16;
        default: lizzieLet35_1_onehotd = 5'd0;
      endcase
    else lizzieLet35_1_onehotd = 5'd0;
  assign _14_d = {lizzieLet35_1_d[115:1], lizzieLet35_1_onehotd[0]};
  assign lizzieLet35_1Lcall_main_mask_Int3_d = {lizzieLet35_1_d[115:1],
                                                lizzieLet35_1_onehotd[1]};
  assign lizzieLet35_1Lcall_main_mask_Int2_d = {lizzieLet35_1_d[115:1],
                                                lizzieLet35_1_onehotd[2]};
  assign lizzieLet35_1Lcall_main_mask_Int1_d = {lizzieLet35_1_d[115:1],
                                                lizzieLet35_1_onehotd[3]};
  assign lizzieLet35_1Lcall_main_mask_Int0_d = {lizzieLet35_1_d[115:1],
                                                lizzieLet35_1_onehotd[4]};
  assign lizzieLet35_1_r = (| (lizzieLet35_1_onehotd & {lizzieLet35_1Lcall_main_mask_Int0_r,
                                                        lizzieLet35_1Lcall_main_mask_Int1_r,
                                                        lizzieLet35_1Lcall_main_mask_Int2_r,
                                                        lizzieLet35_1Lcall_main_mask_Int3_r,
                                                        _14_r}));
  assign lizzieLet35_2_r = lizzieLet35_1_r;
  
  /* demux (Ty CTmain_mask_Int,
       Ty Go) : (lizzieLet35_3,CTmain_mask_Int) (go_17_goMux_data,Go) > [(_13,Go),
                                                                         (lizzieLet35_3Lcall_main_mask_Int3,Go),
                                                                         (lizzieLet35_3Lcall_main_mask_Int2,Go),
                                                                         (lizzieLet35_3Lcall_main_mask_Int1,Go),
                                                                         (lizzieLet35_3Lcall_main_mask_Int0,Go)] */
  logic [4:0] go_17_goMux_data_onehotd;
  always_comb
    if ((lizzieLet35_3_d[0] && go_17_goMux_data_d[0]))
      unique case (lizzieLet35_3_d[3:1])
        3'd0: go_17_goMux_data_onehotd = 5'd1;
        3'd1: go_17_goMux_data_onehotd = 5'd2;
        3'd2: go_17_goMux_data_onehotd = 5'd4;
        3'd3: go_17_goMux_data_onehotd = 5'd8;
        3'd4: go_17_goMux_data_onehotd = 5'd16;
        default: go_17_goMux_data_onehotd = 5'd0;
      endcase
    else go_17_goMux_data_onehotd = 5'd0;
  assign _13_d = go_17_goMux_data_onehotd[0];
  assign lizzieLet35_3Lcall_main_mask_Int3_d = go_17_goMux_data_onehotd[1];
  assign lizzieLet35_3Lcall_main_mask_Int2_d = go_17_goMux_data_onehotd[2];
  assign lizzieLet35_3Lcall_main_mask_Int1_d = go_17_goMux_data_onehotd[3];
  assign lizzieLet35_3Lcall_main_mask_Int0_d = go_17_goMux_data_onehotd[4];
  assign go_17_goMux_data_r = (| (go_17_goMux_data_onehotd & {lizzieLet35_3Lcall_main_mask_Int0_r,
                                                              lizzieLet35_3Lcall_main_mask_Int1_r,
                                                              lizzieLet35_3Lcall_main_mask_Int2_r,
                                                              lizzieLet35_3Lcall_main_mask_Int3_r,
                                                              _13_r}));
  assign lizzieLet35_3_r = go_17_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_main_mask_Int0,Go) > (lizzieLet35_3Lcall_main_mask_Int0_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_main_mask_Int0_bufchan_d;
  logic lizzieLet35_3Lcall_main_mask_Int0_bufchan_r;
  assign lizzieLet35_3Lcall_main_mask_Int0_r = ((! lizzieLet35_3Lcall_main_mask_Int0_bufchan_d[0]) || lizzieLet35_3Lcall_main_mask_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_main_mask_Int0_r)
        lizzieLet35_3Lcall_main_mask_Int0_bufchan_d <= lizzieLet35_3Lcall_main_mask_Int0_d;
  Go_t lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf;
  assign lizzieLet35_3Lcall_main_mask_Int0_bufchan_r = (! lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_d = (lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf[0] ? lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf :
                                                         lizzieLet35_3Lcall_main_mask_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_r && lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf[0]))
        lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_main_mask_Int0_1_argbuf_r) && (! lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf[0])))
        lizzieLet35_3Lcall_main_mask_Int0_bufchan_buf <= lizzieLet35_3Lcall_main_mask_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_main_mask_Int1,Go) > (lizzieLet35_3Lcall_main_mask_Int1_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_main_mask_Int1_bufchan_d;
  logic lizzieLet35_3Lcall_main_mask_Int1_bufchan_r;
  assign lizzieLet35_3Lcall_main_mask_Int1_r = ((! lizzieLet35_3Lcall_main_mask_Int1_bufchan_d[0]) || lizzieLet35_3Lcall_main_mask_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_main_mask_Int1_r)
        lizzieLet35_3Lcall_main_mask_Int1_bufchan_d <= lizzieLet35_3Lcall_main_mask_Int1_d;
  Go_t lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf;
  assign lizzieLet35_3Lcall_main_mask_Int1_bufchan_r = (! lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_d = (lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf[0] ? lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf :
                                                         lizzieLet35_3Lcall_main_mask_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_r && lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf[0]))
        lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_main_mask_Int1_1_argbuf_r) && (! lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf[0])))
        lizzieLet35_3Lcall_main_mask_Int1_bufchan_buf <= lizzieLet35_3Lcall_main_mask_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_main_mask_Int2,Go) > (lizzieLet35_3Lcall_main_mask_Int2_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_main_mask_Int2_bufchan_d;
  logic lizzieLet35_3Lcall_main_mask_Int2_bufchan_r;
  assign lizzieLet35_3Lcall_main_mask_Int2_r = ((! lizzieLet35_3Lcall_main_mask_Int2_bufchan_d[0]) || lizzieLet35_3Lcall_main_mask_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_main_mask_Int2_r)
        lizzieLet35_3Lcall_main_mask_Int2_bufchan_d <= lizzieLet35_3Lcall_main_mask_Int2_d;
  Go_t lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf;
  assign lizzieLet35_3Lcall_main_mask_Int2_bufchan_r = (! lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_d = (lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf[0] ? lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf :
                                                         lizzieLet35_3Lcall_main_mask_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_r && lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf[0]))
        lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_main_mask_Int2_1_argbuf_r) && (! lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf[0])))
        lizzieLet35_3Lcall_main_mask_Int2_bufchan_buf <= lizzieLet35_3Lcall_main_mask_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet35_3Lcall_main_mask_Int3,Go) > (lizzieLet35_3Lcall_main_mask_Int3_1_argbuf,Go) */
  Go_t lizzieLet35_3Lcall_main_mask_Int3_bufchan_d;
  logic lizzieLet35_3Lcall_main_mask_Int3_bufchan_r;
  assign lizzieLet35_3Lcall_main_mask_Int3_r = ((! lizzieLet35_3Lcall_main_mask_Int3_bufchan_d[0]) || lizzieLet35_3Lcall_main_mask_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet35_3Lcall_main_mask_Int3_r)
        lizzieLet35_3Lcall_main_mask_Int3_bufchan_d <= lizzieLet35_3Lcall_main_mask_Int3_d;
  Go_t lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf;
  assign lizzieLet35_3Lcall_main_mask_Int3_bufchan_r = (! lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf[0]);
  assign lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_d = (lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf[0] ? lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf :
                                                         lizzieLet35_3Lcall_main_mask_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_r && lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf[0]))
        lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet35_3Lcall_main_mask_Int3_1_argbuf_r) && (! lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf[0])))
        lizzieLet35_3Lcall_main_mask_Int3_bufchan_buf <= lizzieLet35_3Lcall_main_mask_Int3_bufchan_d;
  
  /* demux (Ty CTmain_mask_Int,
       Ty Pointer_QTree_Int) : (lizzieLet35_4,CTmain_mask_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet35_4Lmain_mask_Intsbos,Pointer_QTree_Int),
                                                                                                           (lizzieLet35_4Lcall_main_mask_Int3,Pointer_QTree_Int),
                                                                                                           (lizzieLet35_4Lcall_main_mask_Int2,Pointer_QTree_Int),
                                                                                                           (lizzieLet35_4Lcall_main_mask_Int1,Pointer_QTree_Int),
                                                                                                           (lizzieLet35_4Lcall_main_mask_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet35_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet35_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet35_4Lmain_mask_Intsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet35_4Lcall_main_mask_Int3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet35_4Lcall_main_mask_Int2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet35_4Lcall_main_mask_Int1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet35_4Lcall_main_mask_Int0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet35_4Lcall_main_mask_Int0_r,
                                                                      lizzieLet35_4Lcall_main_mask_Int1_r,
                                                                      lizzieLet35_4Lcall_main_mask_Int2_r,
                                                                      lizzieLet35_4Lcall_main_mask_Int3_r,
                                                                      lizzieLet35_4Lmain_mask_Intsbos_r}));
  assign lizzieLet35_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet35_4Lcall_main_mask_Int0,Pointer_QTree_Int),
                         (es_1_2_destruct,Pointer_QTree_Int),
                         (es_2_3_destruct,Pointer_QTree_Int),
                         (es_3_6_destruct,Pointer_QTree_Int)] > (lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int,QTree_Int) */
  assign lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_d = QNode_Int_dc((& {lizzieLet35_4Lcall_main_mask_Int0_d[0],
                                                                                                   es_1_2_destruct_d[0],
                                                                                                   es_2_3_destruct_d[0],
                                                                                                   es_3_6_destruct_d[0]}), lizzieLet35_4Lcall_main_mask_Int0_d, es_1_2_destruct_d, es_2_3_destruct_d, es_3_6_destruct_d);
  assign {lizzieLet35_4Lcall_main_mask_Int0_r,
          es_1_2_destruct_r,
          es_2_3_destruct_r,
          es_3_6_destruct_r} = {4 {(lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_r && lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int,QTree_Int) > (lizzieLet39_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d;
  logic lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_r;
  assign lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_r = ((! lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d[0]) || lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d <= {66'd0,
                                                                                         1'd0};
    else
      if (lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_r)
        lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d <= lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_d;
  QTree_Int_t lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf;
  assign lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_r = (! lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf[0] ? lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf :
                                   lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                           1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf[0]))
        lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                             1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf[0])))
        lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_buf <= lizzieLet35_4Lcall_main_mask_Int0_1es_1_2_1es_2_3_1es_3_6_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int0) : [(lizzieLet35_4Lcall_main_mask_Int1,Pointer_QTree_Int),
                                    (es_2_2_destruct,Pointer_QTree_Int),
                                    (es_3_5_destruct,Pointer_QTree_Int),
                                    (sc_0_14_destruct,Pointer_CTmain_mask_Int)] > (lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0,CTmain_mask_Int) */
  assign lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_d = Lcall_main_mask_Int0_dc((& {lizzieLet35_4Lcall_main_mask_Int1_d[0],
                                                                                                                          es_2_2_destruct_d[0],
                                                                                                                          es_3_5_destruct_d[0],
                                                                                                                          sc_0_14_destruct_d[0]}), lizzieLet35_4Lcall_main_mask_Int1_d, es_2_2_destruct_d, es_3_5_destruct_d, sc_0_14_destruct_d);
  assign {lizzieLet35_4Lcall_main_mask_Int1_r,
          es_2_2_destruct_r,
          es_3_5_destruct_r,
          sc_0_14_destruct_r} = {4 {(lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_r && lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0,CTmain_mask_Int) > (lizzieLet38_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d;
  logic lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_r;
  assign lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_r = ((! lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d[0]) || lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d <= {115'd0,
                                                                                                     1'd0};
    else
      if (lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_r)
        lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d <= lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_d;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf;
  assign lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_r = (! lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf[0] ? lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf :
                                   lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf <= {115'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf[0]))
        lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf <= {115'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf[0])))
        lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_buf <= lizzieLet35_4Lcall_main_mask_Int1_1es_2_2_1es_3_5_1sc_0_14_1Lcall_main_mask_Int0_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int1) : [(lizzieLet35_4Lcall_main_mask_Int2,Pointer_QTree_Int),
                                    (es_3_4_destruct,Pointer_QTree_Int),
                                    (sc_0_13_destruct,Pointer_CTmain_mask_Int),
                                    (t1acr_2_destruct,Pointer_QTree_Int),
                                    (q1acm_2_destruct,Pointer_MaskQTree)] > (lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1,CTmain_mask_Int) */
  assign lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_d = Lcall_main_mask_Int1_dc((& {lizzieLet35_4Lcall_main_mask_Int2_d[0],
                                                                                                                                    es_3_4_destruct_d[0],
                                                                                                                                    sc_0_13_destruct_d[0],
                                                                                                                                    t1acr_2_destruct_d[0],
                                                                                                                                    q1acm_2_destruct_d[0]}), lizzieLet35_4Lcall_main_mask_Int2_d, es_3_4_destruct_d, sc_0_13_destruct_d, t1acr_2_destruct_d, q1acm_2_destruct_d);
  assign {lizzieLet35_4Lcall_main_mask_Int2_r,
          es_3_4_destruct_r,
          sc_0_13_destruct_r,
          t1acr_2_destruct_r,
          q1acm_2_destruct_r} = {5 {(lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_r && lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1,CTmain_mask_Int) > (lizzieLet37_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d;
  logic lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_r;
  assign lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_r = ((! lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d[0]) || lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d <= {115'd0,
                                                                                                               1'd0};
    else
      if (lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_r)
        lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d <= lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_d;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf;
  assign lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_r = (! lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf[0]);
  assign lizzieLet37_1_argbuf_d = (lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf[0] ? lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf :
                                   lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf <= {115'd0,
                                                                                                                 1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf[0]))
        lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf <= {115'd0,
                                                                                                                   1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf[0])))
        lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_buf <= lizzieLet35_4Lcall_main_mask_Int2_1es_3_4_1sc_0_13_1t1acr_2_1q1acm_2_1Lcall_main_mask_Int1_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Int,
      Dcon Lcall_main_mask_Int2) : [(lizzieLet35_4Lcall_main_mask_Int3,Pointer_QTree_Int),
                                    (sc_0_12_destruct,Pointer_CTmain_mask_Int),
                                    (t1acr_1_destruct,Pointer_QTree_Int),
                                    (q1acm_1_destruct,Pointer_MaskQTree),
                                    (t2acs_1_destruct,Pointer_QTree_Int),
                                    (q2acn_1_destruct,Pointer_MaskQTree)] > (lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2,CTmain_mask_Int) */
  assign lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_d = Lcall_main_mask_Int2_dc((& {lizzieLet35_4Lcall_main_mask_Int3_d[0],
                                                                                                                                              sc_0_12_destruct_d[0],
                                                                                                                                              t1acr_1_destruct_d[0],
                                                                                                                                              q1acm_1_destruct_d[0],
                                                                                                                                              t2acs_1_destruct_d[0],
                                                                                                                                              q2acn_1_destruct_d[0]}), lizzieLet35_4Lcall_main_mask_Int3_d, sc_0_12_destruct_d, t1acr_1_destruct_d, q1acm_1_destruct_d, t2acs_1_destruct_d, q2acn_1_destruct_d);
  assign {lizzieLet35_4Lcall_main_mask_Int3_r,
          sc_0_12_destruct_r,
          t1acr_1_destruct_r,
          q1acm_1_destruct_r,
          t2acs_1_destruct_r,
          q2acn_1_destruct_r} = {6 {(lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_r && lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_d[0])}};
  
  /* buf (Ty CTmain_mask_Int) : (lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2,CTmain_mask_Int) > (lizzieLet36_1_argbuf,CTmain_mask_Int) */
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d;
  logic lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_r;
  assign lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_r = ((! lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d[0]) || lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d <= {115'd0,
                                                                                                                         1'd0};
    else
      if (lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_r)
        lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d <= lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_d;
  CTmain_mask_Int_t lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf;
  assign lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_r = (! lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf[0] ? lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf :
                                   lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf <= {115'd0,
                                                                                                                           1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf[0]))
        lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf <= {115'd0,
                                                                                                                             1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf[0])))
        lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_buf <= lizzieLet35_4Lcall_main_mask_Int3_1sc_0_12_1t1acr_1_1q1acm_1_1t2acs_1_1q2acn_1_1Lcall_main_mask_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet35_4Lmain_mask_Intsbos,Pointer_QTree_Int) > [(lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                     (lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet35_4Lmain_mask_Intsbos_emitted;
  logic [1:0] lizzieLet35_4Lmain_mask_Intsbos_done;
  assign lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d = {lizzieLet35_4Lmain_mask_Intsbos_d[16:1],
                                                                   (lizzieLet35_4Lmain_mask_Intsbos_d[0] && (! lizzieLet35_4Lmain_mask_Intsbos_emitted[0]))};
  assign lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d = {lizzieLet35_4Lmain_mask_Intsbos_d[16:1],
                                                                   (lizzieLet35_4Lmain_mask_Intsbos_d[0] && (! lizzieLet35_4Lmain_mask_Intsbos_emitted[1]))};
  assign lizzieLet35_4Lmain_mask_Intsbos_done = (lizzieLet35_4Lmain_mask_Intsbos_emitted | ({lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                             lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                           lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet35_4Lmain_mask_Intsbos_r = (& lizzieLet35_4Lmain_mask_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lmain_mask_Intsbos_emitted <= 2'd0;
    else
      lizzieLet35_4Lmain_mask_Intsbos_emitted <= (lizzieLet35_4Lmain_mask_Intsbos_r ? 2'd0 :
                                                  lizzieLet35_4Lmain_mask_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_main_mask_Int_goConst,Go) */
  assign call_main_mask_Int_goConst_d = lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_1_r = call_main_mask_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (main_mask_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign main_mask_Int_resbuf_d = (lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                   lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((main_mask_Int_resbuf_r && lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! main_mask_Int_resbuf_r) && (! lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet35_4Lmain_mask_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_main1_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                     (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_main1_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_main1_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_main1_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_main1_3I#_3_onehotd [1];
  assign \arg0_1Dcon_main1_3I#_3_r  = (| (\arg0_1Dcon_main1_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                              lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_main1_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_r;
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = ((! lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d[0]) || lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d <= {1'd0,
                                                                                       1'd0};
    else
      if (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r)
        lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d <= lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf;
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_r = (! lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf[0] ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf :
                                       lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf <= {1'd0,
                                                                                         1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf[0]))
        lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf <= {1'd0,
                                                                                           1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf[0])))
        lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_buf <= lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int0) : (lizzieLet40_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) > [(es_2_4_destruct,Pointer_QTree_Int),
                                                                                                                            (es_3_8_destruct,Pointer_QTree_Int),
                                                                                                                            (es_4_4_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_19_destruct,Pointer_CTmap''_map''_Int_Int_Int)] */
  logic [3:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted ;
  logic [3:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_done ;
  assign es_2_4_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [19:4],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted [0]))};
  assign es_3_8_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [35:20],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted [1]))};
  assign es_4_4_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [51:36],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted [2]))};
  assign sc_0_19_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [67:52],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted [3]))};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_done  = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted  | ({sc_0_19_destruct_d[0],
                                                                                                                         es_4_4_destruct_d[0],
                                                                                                                         es_3_8_destruct_d[0],
                                                                                                                         es_2_4_destruct_d[0]} & {sc_0_19_destruct_r,
                                                                                                                                                  es_4_4_destruct_r,
                                                                                                                                                  es_3_8_destruct_r,
                                                                                                                                                  es_2_4_destruct_r}));
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_r  = (& \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted  <= 4'd0;
    else
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_emitted  <= (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_r  ? 4'd0 :
                                                                \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int1) : (lizzieLet40_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) > [(es_3_7_destruct,Pointer_QTree_Int),
                                                                                                                            (es_4_3_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_18_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacC_4_destruct,MyDTInt_Bool),
                                                                                                                            (gacD_4_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acE_4_destruct,Int),
                                                                                                                            (q1acH_3_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted ;
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_done ;
  assign es_3_7_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [19:4],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [0]))};
  assign es_4_3_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [35:20],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [1]))};
  assign sc_0_18_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [51:36],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [2]))};
  assign isZacC_4_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [3]));
  assign gacD_4_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [4]));
  assign \v'acE_4_destruct_d  = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [83:52],
                                 (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [5]))};
  assign q1acH_3_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [99:84],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted [6]))};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_done  = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted  | ({q1acH_3_destruct_d[0],
                                                                                                                         \v'acE_4_destruct_d [0],
                                                                                                                         gacD_4_destruct_d[0],
                                                                                                                         isZacC_4_destruct_d[0],
                                                                                                                         sc_0_18_destruct_d[0],
                                                                                                                         es_4_3_destruct_d[0],
                                                                                                                         es_3_7_destruct_d[0]} & {q1acH_3_destruct_r,
                                                                                                                                                  \v'acE_4_destruct_r ,
                                                                                                                                                  gacD_4_destruct_r,
                                                                                                                                                  isZacC_4_destruct_r,
                                                                                                                                                  sc_0_18_destruct_r,
                                                                                                                                                  es_4_3_destruct_r,
                                                                                                                                                  es_3_7_destruct_r}));
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_r  = (& \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted  <= 7'd0;
    else
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_emitted  <= (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_r  ? 7'd0 :
                                                                \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int2) : (lizzieLet40_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) > [(es_4_2_destruct,Pointer_QTree_Int),
                                                                                                                            (sc_0_17_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacC_3_destruct,MyDTInt_Bool),
                                                                                                                            (gacD_3_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acE_3_destruct,Int),
                                                                                                                            (q1acH_2_destruct,Pointer_QTree_Int),
                                                                                                                            (q2acI_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted ;
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_done ;
  assign es_4_2_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [19:4],
                              (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [0]))};
  assign sc_0_17_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [35:20],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [1]))};
  assign isZacC_3_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [2]));
  assign gacD_3_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [3]));
  assign \v'acE_3_destruct_d  = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [67:36],
                                 (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [4]))};
  assign q1acH_2_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [83:68],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [5]))};
  assign q2acI_2_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [99:84],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted [6]))};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_done  = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted  | ({q2acI_2_destruct_d[0],
                                                                                                                         q1acH_2_destruct_d[0],
                                                                                                                         \v'acE_3_destruct_d [0],
                                                                                                                         gacD_3_destruct_d[0],
                                                                                                                         isZacC_3_destruct_d[0],
                                                                                                                         sc_0_17_destruct_d[0],
                                                                                                                         es_4_2_destruct_d[0]} & {q2acI_2_destruct_r,
                                                                                                                                                  q1acH_2_destruct_r,
                                                                                                                                                  \v'acE_3_destruct_r ,
                                                                                                                                                  gacD_3_destruct_r,
                                                                                                                                                  isZacC_3_destruct_r,
                                                                                                                                                  sc_0_17_destruct_r,
                                                                                                                                                  es_4_2_destruct_r}));
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_r  = (& \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted  <= 7'd0;
    else
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_emitted  <= (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_r  ? 7'd0 :
                                                                \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_done );
  
  /* destruct (Ty CTmap''_map''_Int_Int_Int,
          Dcon Lcall_map''_map''_Int_Int_Int3) : (lizzieLet40_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int) > [(sc_0_16_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                                                                                                            (isZacC_2_destruct,MyDTInt_Bool),
                                                                                                                            (gacD_2_destruct,MyDTInt_Int_Int),
                                                                                                                            (v'acE_2_destruct,Int),
                                                                                                                            (q1acH_1_destruct,Pointer_QTree_Int),
                                                                                                                            (q2acI_1_destruct,Pointer_QTree_Int),
                                                                                                                            (q3acJ_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted ;
  logic [6:0] \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_done ;
  assign sc_0_16_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [19:4],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [0]))};
  assign isZacC_2_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [1]));
  assign gacD_2_destruct_d = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [2]));
  assign \v'acE_2_destruct_d  = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [51:20],
                                 (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [3]))};
  assign q1acH_1_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [67:52],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [4]))};
  assign q2acI_1_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [83:68],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [5]))};
  assign q3acJ_1_destruct_d = {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [99:84],
                               (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d [0] && (! \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted [6]))};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_done  = (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted  | ({q3acJ_1_destruct_d[0],
                                                                                                                         q2acI_1_destruct_d[0],
                                                                                                                         q1acH_1_destruct_d[0],
                                                                                                                         \v'acE_2_destruct_d [0],
                                                                                                                         gacD_2_destruct_d[0],
                                                                                                                         isZacC_2_destruct_d[0],
                                                                                                                         sc_0_16_destruct_d[0]} & {q3acJ_1_destruct_r,
                                                                                                                                                   q2acI_1_destruct_r,
                                                                                                                                                   q1acH_1_destruct_r,
                                                                                                                                                   \v'acE_2_destruct_r ,
                                                                                                                                                   gacD_2_destruct_r,
                                                                                                                                                   isZacC_2_destruct_r,
                                                                                                                                                   sc_0_16_destruct_r}));
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_r  = (& \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted  <= 7'd0;
    else
      \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_emitted  <= (\lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_r  ? 7'd0 :
                                                                \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_done );
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty CTmap''_map''_Int_Int_Int) : (lizzieLet40_2,CTmap''_map''_Int_Int_Int) (lizzieLet40_1,CTmap''_map''_Int_Int_Int) > [(_12,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet40_1Lcall_map''_map''_Int_Int_Int3,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet40_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet40_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int),
                                                                                                                              (lizzieLet40_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int)] */
  logic [4:0] lizzieLet40_1_onehotd;
  always_comb
    if ((lizzieLet40_2_d[0] && lizzieLet40_1_d[0]))
      unique case (lizzieLet40_2_d[3:1])
        3'd0: lizzieLet40_1_onehotd = 5'd1;
        3'd1: lizzieLet40_1_onehotd = 5'd2;
        3'd2: lizzieLet40_1_onehotd = 5'd4;
        3'd3: lizzieLet40_1_onehotd = 5'd8;
        3'd4: lizzieLet40_1_onehotd = 5'd16;
        default: lizzieLet40_1_onehotd = 5'd0;
      endcase
    else lizzieLet40_1_onehotd = 5'd0;
  assign _12_d = {lizzieLet40_1_d[99:1], lizzieLet40_1_onehotd[0]};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_d  = {lizzieLet40_1_d[99:1],
                                                            lizzieLet40_1_onehotd[1]};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_d  = {lizzieLet40_1_d[99:1],
                                                            lizzieLet40_1_onehotd[2]};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_d  = {lizzieLet40_1_d[99:1],
                                                            lizzieLet40_1_onehotd[3]};
  assign \lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_d  = {lizzieLet40_1_d[99:1],
                                                            lizzieLet40_1_onehotd[4]};
  assign lizzieLet40_1_r = (| (lizzieLet40_1_onehotd & {\lizzieLet40_1Lcall_map''_map''_Int_Int_Int0_r ,
                                                        \lizzieLet40_1Lcall_map''_map''_Int_Int_Int1_r ,
                                                        \lizzieLet40_1Lcall_map''_map''_Int_Int_Int2_r ,
                                                        \lizzieLet40_1Lcall_map''_map''_Int_Int_Int3_r ,
                                                        _12_r}));
  assign lizzieLet40_2_r = lizzieLet40_1_r;
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty Go) : (lizzieLet40_3,CTmap''_map''_Int_Int_Int) (go_18_goMux_data,Go) > [(_11,Go),
                                                                                   (lizzieLet40_3Lcall_map''_map''_Int_Int_Int3,Go),
                                                                                   (lizzieLet40_3Lcall_map''_map''_Int_Int_Int2,Go),
                                                                                   (lizzieLet40_3Lcall_map''_map''_Int_Int_Int1,Go),
                                                                                   (lizzieLet40_3Lcall_map''_map''_Int_Int_Int0,Go)] */
  logic [4:0] go_18_goMux_data_onehotd;
  always_comb
    if ((lizzieLet40_3_d[0] && go_18_goMux_data_d[0]))
      unique case (lizzieLet40_3_d[3:1])
        3'd0: go_18_goMux_data_onehotd = 5'd1;
        3'd1: go_18_goMux_data_onehotd = 5'd2;
        3'd2: go_18_goMux_data_onehotd = 5'd4;
        3'd3: go_18_goMux_data_onehotd = 5'd8;
        3'd4: go_18_goMux_data_onehotd = 5'd16;
        default: go_18_goMux_data_onehotd = 5'd0;
      endcase
    else go_18_goMux_data_onehotd = 5'd0;
  assign _11_d = go_18_goMux_data_onehotd[0];
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_d  = go_18_goMux_data_onehotd[1];
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_d  = go_18_goMux_data_onehotd[2];
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_d  = go_18_goMux_data_onehotd[3];
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_d  = go_18_goMux_data_onehotd[4];
  assign go_18_goMux_data_r = (| (go_18_goMux_data_onehotd & {\lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_r ,
                                                              \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_r ,
                                                              \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_r ,
                                                              \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_r ,
                                                              _11_r}));
  assign lizzieLet40_3_r = go_18_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet40_3Lcall_map''_map''_Int_Int_Int0,Go) > (lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf,Go) */
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_r  = ((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d [0]) || \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_r )
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_d ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_r  = (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]);
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_d  = (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  :
                                                                     \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r  && \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_1_argbuf_r ) && (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet40_3Lcall_map''_map''_Int_Int_Int1,Go) > (lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf,Go) */
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_r  = ((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d [0]) || \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_r )
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_d ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_r  = (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]);
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_d  = (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  :
                                                                     \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r  && \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_1_argbuf_r ) && (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet40_3Lcall_map''_map''_Int_Int_Int2,Go) > (lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf,Go) */
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_r  = ((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d [0]) || \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_r )
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_d ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_r  = (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]);
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_d  = (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  :
                                                                     \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r  && \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_1_argbuf_r ) && (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet40_3Lcall_map''_map''_Int_Int_Int3,Go) > (lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf,Go) */
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_r  = ((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d [0]) || \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_r )
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_d ;
  Go_t \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_r  = (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]);
  assign \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_d  = (\lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  :
                                                                     \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r  && \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_1_argbuf_r ) && (! \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_buf  <= \lizzieLet40_3Lcall_map''_map''_Int_Int_Int3_bufchan_d ;
  
  /* demux (Ty CTmap''_map''_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet40_4,CTmap''_map''_Int_Int_Int) (srtarg_0_3_goMux_mux,Pointer_QTree_Int) > [(lizzieLet40_4Lmap''_map''_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                     (lizzieLet40_4Lcall_map''_map''_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                     (lizzieLet40_4Lcall_map''_map''_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                     (lizzieLet40_4Lcall_map''_map''_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                     (lizzieLet40_4Lcall_map''_map''_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet40_4_d[0] && srtarg_0_3_goMux_mux_d[0]))
      unique case (lizzieLet40_4_d[3:1])
        3'd0: srtarg_0_3_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_3_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_3_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_3_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_3_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_3_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_3_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                          srtarg_0_3_goMux_mux_onehotd[0]};
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[1]};
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[2]};
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[3]};
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_d  = {srtarg_0_3_goMux_mux_d[16:1],
                                                            srtarg_0_3_goMux_mux_onehotd[4]};
  assign srtarg_0_3_goMux_mux_r = (| (srtarg_0_3_goMux_mux_onehotd & {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_r ,
                                                                      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_r ,
                                                                      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_r ,
                                                                      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_r ,
                                                                      \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_r }));
  assign lizzieLet40_4_r = srtarg_0_3_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet40_4Lcall_map''_map''_Int_Int_Int0,Pointer_QTree_Int),
                         (es_2_4_destruct,Pointer_QTree_Int),
                         (es_3_8_destruct,Pointer_QTree_Int),
                         (es_4_4_destruct,Pointer_QTree_Int)] > (lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int,QTree_Int) */
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_d [0],
                                                                                                               es_2_4_destruct_d[0],
                                                                                                               es_3_8_destruct_d[0],
                                                                                                               es_4_4_destruct_d[0]}), \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_d , es_2_4_destruct_d, es_3_8_destruct_d, es_4_4_destruct_d);
  assign {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_r ,
          es_2_4_destruct_r,
          es_3_8_destruct_r,
          es_4_4_destruct_r} = {4 {(\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_r  && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int,QTree_Int) > (lizzieLet44_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_r ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_r  = ((! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d [0]) || \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                     1'd0};
    else
      if (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_r )
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_d ;
  QTree_Int_t \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_r  = (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet44_1_argbuf_d = (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf [0] ? \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf  :
                                   \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet44_1_argbuf_r && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf [0]))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet44_1_argbuf_r) && (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf [0])))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_buf  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int0_1es_2_4_1es_3_8_1es_4_4_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int0) : [(lizzieLet40_4Lcall_map''_map''_Int_Int_Int1,Pointer_QTree_Int),
                                              (es_3_7_destruct,Pointer_QTree_Int),
                                              (es_4_3_destruct,Pointer_QTree_Int),
                                              (sc_0_18_destruct,Pointer_CTmap''_map''_Int_Int_Int)] > (lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d  = \Lcall_map''_map''_Int_Int_Int0_dc ((& {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_d [0],
                                                                                                                                                            es_3_7_destruct_d[0],
                                                                                                                                                            es_4_3_destruct_d[0],
                                                                                                                                                            sc_0_18_destruct_d[0]}), \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_d , es_3_7_destruct_d, es_4_3_destruct_d, sc_0_18_destruct_d);
  assign {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_r ,
          es_3_7_destruct_r,
          es_4_3_destruct_r,
          sc_0_18_destruct_r} = {4 {(\lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r  && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0,CTmap''_map''_Int_Int_Int) > (lizzieLet43_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r  = ((! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d [0]) || \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= {99'd0,
                                                                                                                           1'd0};
    else
      if (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_r )
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_r  = (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]);
  assign lizzieLet43_1_argbuf_d = (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  :
                                   \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                             1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                               1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_buf  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int1_1es_3_7_1es_4_3_1sc_0_18_1Lcall_map''_map''_Int_Int_Int0_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int1) : [(lizzieLet40_4Lcall_map''_map''_Int_Int_Int2,Pointer_QTree_Int),
                                              (es_4_2_destruct,Pointer_QTree_Int),
                                              (sc_0_17_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                              (isZacC_3_1,MyDTInt_Bool),
                                              (gacD_3_1,MyDTInt_Int_Int),
                                              (v'acE_3_1,Int),
                                              (q1acH_2_destruct,Pointer_QTree_Int)] > (lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_d  = \Lcall_map''_map''_Int_Int_Int1_dc ((& {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_d [0],
                                                                                                                                                                                        es_4_2_destruct_d[0],
                                                                                                                                                                                        sc_0_17_destruct_d[0],
                                                                                                                                                                                        isZacC_3_1_d[0],
                                                                                                                                                                                        gacD_3_1_d[0],
                                                                                                                                                                                        \v'acE_3_1_d [0],
                                                                                                                                                                                        q1acH_2_destruct_d[0]}), \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_d , es_4_2_destruct_d, sc_0_17_destruct_d, isZacC_3_1_d, gacD_3_1_d, \v'acE_3_1_d , q1acH_2_destruct_d);
  assign {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_r ,
          es_4_2_destruct_r,
          sc_0_17_destruct_r,
          isZacC_3_1_r,
          gacD_3_1_r,
          \v'acE_3_1_r ,
          q1acH_2_destruct_r} = {7 {(\lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_r  && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1,CTmap''_map''_Int_Int_Int) > (lizzieLet42_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_r  = ((! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d [0]) || \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= {99'd0,
                                                                                                                                                       1'd0};
    else
      if (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_r )
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_r  = (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]);
  assign lizzieLet42_1_argbuf_d = (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  :
                                   \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                         1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                           1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_buf  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int2_1es_4_2_1sc_0_17_1isZacC_3_1gacD_3_1v'acE_3_1q1acH_2_1Lcall_map''_map''_Int_Int_Int1_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Int_Int_Int,
      Dcon Lcall_map''_map''_Int_Int_Int2) : [(lizzieLet40_4Lcall_map''_map''_Int_Int_Int3,Pointer_QTree_Int),
                                              (sc_0_16_destruct,Pointer_CTmap''_map''_Int_Int_Int),
                                              (isZacC_2_1,MyDTInt_Bool),
                                              (gacD_2_1,MyDTInt_Int_Int),
                                              (v'acE_2_1,Int),
                                              (q1acH_1_destruct,Pointer_QTree_Int),
                                              (q2acI_1_destruct,Pointer_QTree_Int)] > (lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) */
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_d  = \Lcall_map''_map''_Int_Int_Int2_dc ((& {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_d [0],
                                                                                                                                                                                         sc_0_16_destruct_d[0],
                                                                                                                                                                                         isZacC_2_1_d[0],
                                                                                                                                                                                         gacD_2_1_d[0],
                                                                                                                                                                                         \v'acE_2_1_d [0],
                                                                                                                                                                                         q1acH_1_destruct_d[0],
                                                                                                                                                                                         q2acI_1_destruct_d[0]}), \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_d , sc_0_16_destruct_d, isZacC_2_1_d, gacD_2_1_d, \v'acE_2_1_d , q1acH_1_destruct_d, q2acI_1_destruct_d);
  assign {\lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_r ,
          sc_0_16_destruct_r,
          isZacC_2_1_r,
          gacD_2_1_r,
          \v'acE_2_1_r ,
          q1acH_1_destruct_r,
          q2acI_1_destruct_r} = {7 {(\lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_r  && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_d [0])}};
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2,CTmap''_map''_Int_Int_Int) > (lizzieLet41_1_argbuf,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_r  = ((! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d [0]) || \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= {99'd0,
                                                                                                                                                        1'd0};
    else
      if (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_r )
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_d ;
  \CTmap''_map''_Int_Int_Int_t  \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_r  = (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]);
  assign lizzieLet41_1_argbuf_d = (\lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  :
                                   \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                          1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                            1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_buf  <= \lizzieLet40_4Lcall_map''_map''_Int_Int_Int3_1sc_0_16_1isZacC_2_1gacD_2_1v'acE_2_1q1acH_1_1q2acI_1_1Lcall_map''_map''_Int_Int_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet40_4Lmap''_map''_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                               (lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted ;
  logic [1:0] \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_done ;
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d [16:1],
                                                                               (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d [0] && (! \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted [0]))};
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d [16:1],
                                                                               (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_d [0] && (! \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted [1]))};
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_done  = (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted  | ({\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                     \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                               \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_r  = (& \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_emitted  <= (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_r  ? 2'd0 :
                                                              \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_map''_map''_Int_Int_Int_goConst,Go) */
  assign \call_map''_map''_Int_Int_Int_goConst_d  = \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_1_r  = \call_map''_map''_Int_Int_Int_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (map''_map''_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                     1'd0};
    else
      if (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_r )
        \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Int_t \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \map''_map''_Int_Int_Int_resbuf_d  = (\lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  :
                                               \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
    else
      if ((\map''_map''_Int_Int_Int_resbuf_r  && \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                         1'd0};
      else if (((! \map''_map''_Int_Int_Int_resbuf_r ) && (! \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet40_4Lmap''_map''_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1acV_destruct,Pointer_QTree_Int),
                                                                 (q2acW_destruct,Pointer_QTree_Int),
                                                                 (q3acX_destruct,Pointer_QTree_Int),
                                                                 (q4acY_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1acV_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2acW_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3acX_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4acY_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4acY_destruct_d[0],
                                                                         q3acX_destruct_d[0],
                                                                         q2acW_destruct_d[0],
                                                                         q1acV_destruct_d[0]} & {q4acY_destruct_r,
                                                                                                 q3acX_destruct_r,
                                                                                                 q2acW_destruct_r,
                                                                                                 q1acV_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_10,QTree_Int),
                                                                            (_9,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_8,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _10_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _9_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _8_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_8_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _9_r,
                                                      _10_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_8_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                 (lizzieLet4_3QVal_Int,Go),
                                                                 (lizzieLet4_3QNode_Int,Go),
                                                                 (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_8_goMux_data_onehotd = 4'd1;
        2'd1: go_8_goMux_data_onehotd = 4'd2;
        2'd2: go_8_goMux_data_onehotd = 4'd4;
        2'd3: go_8_goMux_data_onehotd = 4'd8;
        default: go_8_goMux_data_onehotd = 4'd0;
      endcase
    else go_8_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_8_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_8_goMux_data_onehotd[3];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                            lizzieLet4_3QNode_Int_r,
                                                            lizzieLet4_3QVal_Int_r,
                                                            lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_8_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet14_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet14_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C4) (go_15_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                            go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                      go_15_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_15_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet26_3Lcall_$wnnz_Int0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_15_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet15_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz_Int) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                (q4acY_destruct,Pointer_QTree_Int),
                                (q3acX_destruct,Pointer_QTree_Int),
                                (q2acW_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3,CT$wnnz_Int) */
  assign lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_d = Lcall_$wnnz_Int3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                                  q4acY_destruct_d[0],
                                                                                                  q3acX_destruct_d[0],
                                                                                                  q2acW_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4acY_destruct_d, q3acX_destruct_d, q2acW_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4acY_destruct_r,
          q3acX_destruct_r,
          q2acW_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_r && lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3,CT$wnnz_Int) > (lizzieLet5_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_r = ((! lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d <= {115'd0,
                                                                                 1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_r)
        lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d <= lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_d;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                     1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4acY_1q3acX_1q2acW_1Lcall_$wnnz_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_1QNode_Int,QTree_Int) > [(q1acQ_destruct,Pointer_QTree_Int),
                                                                 (q2acR_destruct,Pointer_QTree_Int),
                                                                 (q3acS_destruct,Pointer_QTree_Int),
                                                                 (q4acT_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_1QNode_Int_done;
  assign q1acQ_destruct_d = {lizzieLet6_1QNode_Int_d[18:3],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[0]))};
  assign q2acR_destruct_d = {lizzieLet6_1QNode_Int_d[34:19],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[1]))};
  assign q3acS_destruct_d = {lizzieLet6_1QNode_Int_d[50:35],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[2]))};
  assign q4acT_destruct_d = {lizzieLet6_1QNode_Int_d[66:51],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[3]))};
  assign lizzieLet6_1QNode_Int_done = (lizzieLet6_1QNode_Int_emitted | ({q4acT_destruct_d[0],
                                                                         q3acS_destruct_d[0],
                                                                         q2acR_destruct_d[0],
                                                                         q1acQ_destruct_d[0]} & {q4acT_destruct_r,
                                                                                                 q3acS_destruct_r,
                                                                                                 q2acR_destruct_r,
                                                                                                 q1acQ_destruct_r}));
  assign lizzieLet6_1QNode_Int_r = (& lizzieLet6_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Int_emitted <= (lizzieLet6_1QNode_Int_r ? 4'd0 :
                                        lizzieLet6_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_1QVal_Int,QTree_Int) > [(vacP_destruct,Int)] */
  assign vacP_destruct_d = {lizzieLet6_1QVal_Int_d[34:3],
                            lizzieLet6_1QVal_Int_d[0]};
  assign lizzieLet6_1QVal_Int_r = vacP_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_2,QTree_Int) (lizzieLet6_1,QTree_Int) > [(_7,QTree_Int),
                                                                            (lizzieLet6_1QVal_Int,QTree_Int),
                                                                            (lizzieLet6_1QNode_Int,QTree_Int),
                                                                            (_6,QTree_Int)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _7_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Int_d = {lizzieLet6_1_d[66:1],
                                   lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Int_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[2]};
  assign _6_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_6_r,
                                                      lizzieLet6_1QNode_Int_r,
                                                      lizzieLet6_1QVal_Int_r,
                                                      _7_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_3,QTree_Int) (gacM_goMux_mux,MyDTInt_Int_Int) > [(_5,MyDTInt_Int_Int),
                                                                                          (lizzieLet6_3QVal_Int,MyDTInt_Int_Int),
                                                                                          (lizzieLet6_3QNode_Int,MyDTInt_Int_Int),
                                                                                          (_4,MyDTInt_Int_Int)] */
  logic [3:0] gacM_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && gacM_goMux_mux_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: gacM_goMux_mux_onehotd = 4'd1;
        2'd1: gacM_goMux_mux_onehotd = 4'd2;
        2'd2: gacM_goMux_mux_onehotd = 4'd4;
        2'd3: gacM_goMux_mux_onehotd = 4'd8;
        default: gacM_goMux_mux_onehotd = 4'd0;
      endcase
    else gacM_goMux_mux_onehotd = 4'd0;
  assign _5_d = gacM_goMux_mux_onehotd[0];
  assign lizzieLet6_3QVal_Int_d = gacM_goMux_mux_onehotd[1];
  assign lizzieLet6_3QNode_Int_d = gacM_goMux_mux_onehotd[2];
  assign _4_d = gacM_goMux_mux_onehotd[3];
  assign gacM_goMux_mux_r = (| (gacM_goMux_mux_onehotd & {_4_r,
                                                          lizzieLet6_3QNode_Int_r,
                                                          lizzieLet6_3QVal_Int_r,
                                                          _5_r}));
  assign lizzieLet6_3_r = gacM_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_3QNode_Int,MyDTInt_Int_Int) > [(lizzieLet6_3QNode_Int_1,MyDTInt_Int_Int),
                                                                       (lizzieLet6_3QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_3QNode_Int_emitted;
  logic [1:0] lizzieLet6_3QNode_Int_done;
  assign lizzieLet6_3QNode_Int_1_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[0]));
  assign lizzieLet6_3QNode_Int_2_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[1]));
  assign lizzieLet6_3QNode_Int_done = (lizzieLet6_3QNode_Int_emitted | ({lizzieLet6_3QNode_Int_2_d[0],
                                                                         lizzieLet6_3QNode_Int_1_d[0]} & {lizzieLet6_3QNode_Int_2_r,
                                                                                                          lizzieLet6_3QNode_Int_1_r}));
  assign lizzieLet6_3QNode_Int_r = (& lizzieLet6_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QNode_Int_emitted <= (lizzieLet6_3QNode_Int_r ? 2'd0 :
                                        lizzieLet6_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_3QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_bufchan_d;
  logic lizzieLet6_3QNode_Int_2_bufchan_r;
  assign lizzieLet6_3QNode_Int_2_r = ((! lizzieLet6_3QNode_Int_2_bufchan_d[0]) || lizzieLet6_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNode_Int_2_r)
        lizzieLet6_3QNode_Int_2_bufchan_d <= lizzieLet6_3QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet6_3QNode_Int_2_bufchan_buf;
  assign lizzieLet6_3QNode_Int_2_bufchan_r = (! lizzieLet6_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QNode_Int_2_argbuf_d = (lizzieLet6_3QNode_Int_2_bufchan_buf[0] ? lizzieLet6_3QNode_Int_2_bufchan_buf :
                                             lizzieLet6_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNode_Int_2_argbuf_r && lizzieLet6_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNode_Int_2_argbuf_r) && (! lizzieLet6_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= lizzieLet6_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_3QVal_Int,MyDTInt_Int_Int) > (lizzieLet6_3QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_bufchan_d;
  logic lizzieLet6_3QVal_Int_bufchan_r;
  assign lizzieLet6_3QVal_Int_r = ((! lizzieLet6_3QVal_Int_bufchan_d[0]) || lizzieLet6_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QVal_Int_r)
        lizzieLet6_3QVal_Int_bufchan_d <= lizzieLet6_3QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet6_3QVal_Int_bufchan_buf;
  assign lizzieLet6_3QVal_Int_bufchan_r = (! lizzieLet6_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_3QVal_Int_1_argbuf_d = (lizzieLet6_3QVal_Int_bufchan_buf[0] ? lizzieLet6_3QVal_Int_bufchan_buf :
                                            lizzieLet6_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QVal_Int_1_argbuf_r && lizzieLet6_3QVal_Int_bufchan_buf[0]))
        lizzieLet6_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QVal_Int_1_argbuf_r) && (! lizzieLet6_3QVal_Int_bufchan_buf[0])))
        lizzieLet6_3QVal_Int_bufchan_buf <= lizzieLet6_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_4,QTree_Int) (go_9_goMux_data,Go) > [(lizzieLet6_4QNone_Int,Go),
                                                                 (lizzieLet6_4QVal_Int,Go),
                                                                 (lizzieLet6_4QNode_Int,Go),
                                                                 (lizzieLet6_4QError_Int,Go)] */
  logic [3:0] go_9_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && go_9_goMux_data_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: go_9_goMux_data_onehotd = 4'd1;
        2'd1: go_9_goMux_data_onehotd = 4'd2;
        2'd2: go_9_goMux_data_onehotd = 4'd4;
        2'd3: go_9_goMux_data_onehotd = 4'd8;
        default: go_9_goMux_data_onehotd = 4'd0;
      endcase
    else go_9_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_4QNone_Int_d = go_9_goMux_data_onehotd[0];
  assign lizzieLet6_4QVal_Int_d = go_9_goMux_data_onehotd[1];
  assign lizzieLet6_4QNode_Int_d = go_9_goMux_data_onehotd[2];
  assign lizzieLet6_4QError_Int_d = go_9_goMux_data_onehotd[3];
  assign go_9_goMux_data_r = (| (go_9_goMux_data_onehotd & {lizzieLet6_4QError_Int_r,
                                                            lizzieLet6_4QNode_Int_r,
                                                            lizzieLet6_4QVal_Int_r,
                                                            lizzieLet6_4QNone_Int_r}));
  assign lizzieLet6_4_r = go_9_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_4QError_Int,Go) > [(lizzieLet6_4QError_Int_1,Go),
                                              (lizzieLet6_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QError_Int_emitted;
  logic [1:0] lizzieLet6_4QError_Int_done;
  assign lizzieLet6_4QError_Int_1_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[0]));
  assign lizzieLet6_4QError_Int_2_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[1]));
  assign lizzieLet6_4QError_Int_done = (lizzieLet6_4QError_Int_emitted | ({lizzieLet6_4QError_Int_2_d[0],
                                                                           lizzieLet6_4QError_Int_1_d[0]} & {lizzieLet6_4QError_Int_2_r,
                                                                                                             lizzieLet6_4QError_Int_1_r}));
  assign lizzieLet6_4QError_Int_r = (& lizzieLet6_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QError_Int_emitted <= (lizzieLet6_4QError_Int_r ? 2'd0 :
                                         lizzieLet6_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_4QError_Int_1,Go)] > (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_4QError_Int_1_d[0]}), lizzieLet6_4QError_Int_1_d);
  assign {lizzieLet6_4QError_Int_1_r} = {1 {(lizzieLet6_4QError_Int_1QError_Int_r && lizzieLet6_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_4QError_Int_1QError_Int_r = ((! lizzieLet6_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QError_Int_1QError_Int_r)
        lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= lizzieLet6_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_4QError_Int_1QError_Int_bufchan_buf :
                                  lizzieLet6_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QError_Int_2,Go) > (lizzieLet6_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QError_Int_2_bufchan_d;
  logic lizzieLet6_4QError_Int_2_bufchan_r;
  assign lizzieLet6_4QError_Int_2_r = ((! lizzieLet6_4QError_Int_2_bufchan_d[0]) || lizzieLet6_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QError_Int_2_r)
        lizzieLet6_4QError_Int_2_bufchan_d <= lizzieLet6_4QError_Int_2_d;
  Go_t lizzieLet6_4QError_Int_2_bufchan_buf;
  assign lizzieLet6_4QError_Int_2_bufchan_r = (! lizzieLet6_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QError_Int_2_argbuf_d = (lizzieLet6_4QError_Int_2_bufchan_buf[0] ? lizzieLet6_4QError_Int_2_bufchan_buf :
                                              lizzieLet6_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QError_Int_2_argbuf_r && lizzieLet6_4QError_Int_2_bufchan_buf[0]))
        lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QError_Int_2_argbuf_r) && (! lizzieLet6_4QError_Int_2_bufchan_buf[0])))
        lizzieLet6_4QError_Int_2_bufchan_buf <= lizzieLet6_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNode_Int,Go) > (lizzieLet6_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QNode_Int_bufchan_d;
  logic lizzieLet6_4QNode_Int_bufchan_r;
  assign lizzieLet6_4QNode_Int_r = ((! lizzieLet6_4QNode_Int_bufchan_d[0]) || lizzieLet6_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNode_Int_r)
        lizzieLet6_4QNode_Int_bufchan_d <= lizzieLet6_4QNode_Int_d;
  Go_t lizzieLet6_4QNode_Int_bufchan_buf;
  assign lizzieLet6_4QNode_Int_bufchan_r = (! lizzieLet6_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_4QNode_Int_1_argbuf_d = (lizzieLet6_4QNode_Int_bufchan_buf[0] ? lizzieLet6_4QNode_Int_bufchan_buf :
                                             lizzieLet6_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNode_Int_1_argbuf_r && lizzieLet6_4QNode_Int_bufchan_buf[0]))
        lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNode_Int_1_argbuf_r) && (! lizzieLet6_4QNode_Int_bufchan_buf[0])))
        lizzieLet6_4QNode_Int_bufchan_buf <= lizzieLet6_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4QNone_Int,Go) > [(lizzieLet6_4QNone_Int_1,Go),
                                             (lizzieLet6_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QNone_Int_emitted;
  logic [1:0] lizzieLet6_4QNone_Int_done;
  assign lizzieLet6_4QNone_Int_1_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[0]));
  assign lizzieLet6_4QNone_Int_2_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[1]));
  assign lizzieLet6_4QNone_Int_done = (lizzieLet6_4QNone_Int_emitted | ({lizzieLet6_4QNone_Int_2_d[0],
                                                                         lizzieLet6_4QNone_Int_1_d[0]} & {lizzieLet6_4QNone_Int_2_r,
                                                                                                          lizzieLet6_4QNone_Int_1_r}));
  assign lizzieLet6_4QNone_Int_r = (& lizzieLet6_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QNone_Int_emitted <= (lizzieLet6_4QNone_Int_r ? 2'd0 :
                                        lizzieLet6_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_4QNone_Int_1,Go)] > (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet6_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_4QNone_Int_1_d[0]}), lizzieLet6_4QNone_Int_1_d);
  assign {lizzieLet6_4QNone_Int_1_r} = {1 {(lizzieLet6_4QNone_Int_1QNone_Int_r && lizzieLet6_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet7_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet6_4QNone_Int_1QNone_Int_r = ((! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QNone_Int_1QNone_Int_r)
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet6_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf :
                                  lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNone_Int_2,Go) > (lizzieLet6_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QNone_Int_2_bufchan_d;
  logic lizzieLet6_4QNone_Int_2_bufchan_r;
  assign lizzieLet6_4QNone_Int_2_r = ((! lizzieLet6_4QNone_Int_2_bufchan_d[0]) || lizzieLet6_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNone_Int_2_r)
        lizzieLet6_4QNone_Int_2_bufchan_d <= lizzieLet6_4QNone_Int_2_d;
  Go_t lizzieLet6_4QNone_Int_2_bufchan_buf;
  assign lizzieLet6_4QNone_Int_2_bufchan_r = (! lizzieLet6_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QNone_Int_2_argbuf_d = (lizzieLet6_4QNone_Int_2_bufchan_buf[0] ? lizzieLet6_4QNone_Int_2_bufchan_buf :
                                             lizzieLet6_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNone_Int_2_argbuf_r && lizzieLet6_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNone_Int_2_argbuf_r) && (! lizzieLet6_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= lizzieLet6_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet6_4QNone_Int_2_argbuf,Go),
                           (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf,Go),
                           (lizzieLet6_4QVal_Int_2_argbuf,Go),
                           (lizzieLet6_4QError_Int_2_argbuf,Go)] > (go_16_goMux_choice,C4) (go_16_goMux_data,Go) */
  logic [3:0] lizzieLet6_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_select_d = ((| lizzieLet6_4QNone_Int_2_argbuf_select_q) ? lizzieLet6_4QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet6_4QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet6_4QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet6_4QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet6_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet6_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_emit_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_emit_d = (lizzieLet6_4QNone_Int_2_argbuf_emit_q | ({go_16_goMux_choice_d[0],
                                                                                            go_16_goMux_data_d[0]} & {go_16_goMux_choice_r,
                                                                                                                      go_16_goMux_data_r}));
  logic lizzieLet6_4QNone_Int_2_argbuf_done;
  assign lizzieLet6_4QNone_Int_2_argbuf_done = (& lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet6_4QError_Int_2_argbuf_r,
          lizzieLet6_4QVal_Int_2_argbuf_r,
          lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_r,
          lizzieLet6_4QNone_Int_2_argbuf_r} = (lizzieLet6_4QNone_Int_2_argbuf_done ? lizzieLet6_4QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_16_goMux_data_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QNone_Int_2_argbuf_d :
                               ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet30_3Lcall_kron_kron_Int_Int_Int0_1_argbuf_d :
                                ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QVal_Int_2_argbuf_d :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_16_goMux_choice_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet6_4QVal_Int,Go) > [(lizzieLet6_4QVal_Int_1,Go),
                                            (lizzieLet6_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QVal_Int_emitted;
  logic [1:0] lizzieLet6_4QVal_Int_done;
  assign lizzieLet6_4QVal_Int_1_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[0]));
  assign lizzieLet6_4QVal_Int_2_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[1]));
  assign lizzieLet6_4QVal_Int_done = (lizzieLet6_4QVal_Int_emitted | ({lizzieLet6_4QVal_Int_2_d[0],
                                                                       lizzieLet6_4QVal_Int_1_d[0]} & {lizzieLet6_4QVal_Int_2_r,
                                                                                                       lizzieLet6_4QVal_Int_1_r}));
  assign lizzieLet6_4QVal_Int_r = (& lizzieLet6_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QVal_Int_emitted <= (lizzieLet6_4QVal_Int_r ? 2'd0 :
                                       lizzieLet6_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Int_1,Go) > (lizzieLet6_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Int_1_bufchan_d;
  logic lizzieLet6_4QVal_Int_1_bufchan_r;
  assign lizzieLet6_4QVal_Int_1_r = ((! lizzieLet6_4QVal_Int_1_bufchan_d[0]) || lizzieLet6_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_1_r)
        lizzieLet6_4QVal_Int_1_bufchan_d <= lizzieLet6_4QVal_Int_1_d;
  Go_t lizzieLet6_4QVal_Int_1_bufchan_buf;
  assign lizzieLet6_4QVal_Int_1_bufchan_r = (! lizzieLet6_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_1_argbuf_d = (lizzieLet6_4QVal_Int_1_bufchan_buf[0] ? lizzieLet6_4QVal_Int_1_bufchan_buf :
                                            lizzieLet6_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_1_argbuf_r && lizzieLet6_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_1_argbuf_r) && (! lizzieLet6_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= lizzieLet6_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) : [(lizzieLet6_4QVal_Int_1_argbuf,Go),
                                                                                (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                                                                (lizzieLet6_3QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                                                                (vacP_1_argbuf,Int),
                                                                                (lizzieLet6_6QVal_Int_1_argbuf,Pointer_QTree_Int)] > (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) */
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d  = TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_dc((& {lizzieLet6_4QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_5QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_3QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                 vacP_1_argbuf_d[0],
                                                                                                                                                                                 lizzieLet6_6QVal_Int_1_argbuf_d[0]}), lizzieLet6_4QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_1_argbuf_d, lizzieLet6_3QVal_Int_1_argbuf_d, vacP_1_argbuf_d, lizzieLet6_6QVal_Int_1_argbuf_d);
  assign {lizzieLet6_4QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_1_argbuf_r,
          lizzieLet6_3QVal_Int_1_argbuf_r,
          vacP_1_argbuf_r,
          lizzieLet6_6QVal_Int_1_argbuf_r} = {5 {(\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Int_2,Go) > (lizzieLet6_4QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Int_2_bufchan_d;
  logic lizzieLet6_4QVal_Int_2_bufchan_r;
  assign lizzieLet6_4QVal_Int_2_r = ((! lizzieLet6_4QVal_Int_2_bufchan_d[0]) || lizzieLet6_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_2_r)
        lizzieLet6_4QVal_Int_2_bufchan_d <= lizzieLet6_4QVal_Int_2_d;
  Go_t lizzieLet6_4QVal_Int_2_bufchan_buf;
  assign lizzieLet6_4QVal_Int_2_bufchan_r = (! lizzieLet6_4QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_2_argbuf_d = (lizzieLet6_4QVal_Int_2_bufchan_buf[0] ? lizzieLet6_4QVal_Int_2_bufchan_buf :
                                            lizzieLet6_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_2_argbuf_r && lizzieLet6_4QVal_Int_2_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_2_argbuf_r) && (! lizzieLet6_4QVal_Int_2_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_2_bufchan_buf <= lizzieLet6_4QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_5,QTree_Int) (isZacL_goMux_mux,MyDTInt_Bool) > [(_3,MyDTInt_Bool),
                                                                                      (lizzieLet6_5QVal_Int,MyDTInt_Bool),
                                                                                      (lizzieLet6_5QNode_Int,MyDTInt_Bool),
                                                                                      (_2,MyDTInt_Bool)] */
  logic [3:0] isZacL_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && isZacL_goMux_mux_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: isZacL_goMux_mux_onehotd = 4'd1;
        2'd1: isZacL_goMux_mux_onehotd = 4'd2;
        2'd2: isZacL_goMux_mux_onehotd = 4'd4;
        2'd3: isZacL_goMux_mux_onehotd = 4'd8;
        default: isZacL_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacL_goMux_mux_onehotd = 4'd0;
  assign _3_d = isZacL_goMux_mux_onehotd[0];
  assign lizzieLet6_5QVal_Int_d = isZacL_goMux_mux_onehotd[1];
  assign lizzieLet6_5QNode_Int_d = isZacL_goMux_mux_onehotd[2];
  assign _2_d = isZacL_goMux_mux_onehotd[3];
  assign isZacL_goMux_mux_r = (| (isZacL_goMux_mux_onehotd & {_2_r,
                                                              lizzieLet6_5QNode_Int_r,
                                                              lizzieLet6_5QVal_Int_r,
                                                              _3_r}));
  assign lizzieLet6_5_r = isZacL_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int,MyDTInt_Bool) > [(lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                                                 (lizzieLet6_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_5QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_1_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_2_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_done = (lizzieLet6_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_2_d[0],
                                                                         lizzieLet6_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_2_r,
                                                                                                          lizzieLet6_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_r = (& lizzieLet6_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_r ? 2'd0 :
                                        lizzieLet6_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_2_r)
        lizzieLet6_5QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_2_bufchan_buf :
                                             lizzieLet6_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QVal_Int,MyDTInt_Bool) > (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_r = ((! lizzieLet6_5QVal_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_r)
        lizzieLet6_5QVal_Int_bufchan_d <= lizzieLet6_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_bufchan_r = (! lizzieLet6_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_bufchan_buf :
                                            lizzieLet6_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_bufchan_buf <= lizzieLet6_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet6_6,QTree_Int) (m2acO_goMux_mux,Pointer_QTree_Int) > [(_1,Pointer_QTree_Int),
                                                                                               (lizzieLet6_6QVal_Int,Pointer_QTree_Int),
                                                                                               (lizzieLet6_6QNode_Int,Pointer_QTree_Int),
                                                                                               (_0,Pointer_QTree_Int)] */
  logic [3:0] m2acO_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && m2acO_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: m2acO_goMux_mux_onehotd = 4'd1;
        2'd1: m2acO_goMux_mux_onehotd = 4'd2;
        2'd2: m2acO_goMux_mux_onehotd = 4'd4;
        2'd3: m2acO_goMux_mux_onehotd = 4'd8;
        default: m2acO_goMux_mux_onehotd = 4'd0;
      endcase
    else m2acO_goMux_mux_onehotd = 4'd0;
  assign _1_d = {m2acO_goMux_mux_d[16:1],
                 m2acO_goMux_mux_onehotd[0]};
  assign lizzieLet6_6QVal_Int_d = {m2acO_goMux_mux_d[16:1],
                                   m2acO_goMux_mux_onehotd[1]};
  assign lizzieLet6_6QNode_Int_d = {m2acO_goMux_mux_d[16:1],
                                    m2acO_goMux_mux_onehotd[2]};
  assign _0_d = {m2acO_goMux_mux_d[16:1],
                 m2acO_goMux_mux_onehotd[3]};
  assign m2acO_goMux_mux_r = (| (m2acO_goMux_mux_onehotd & {_0_r,
                                                            lizzieLet6_6QNode_Int_r,
                                                            lizzieLet6_6QVal_Int_r,
                                                            _1_r}));
  assign lizzieLet6_6_r = m2acO_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet6_6QNode_Int,Pointer_QTree_Int) > [(lizzieLet6_6QNode_Int_1,Pointer_QTree_Int),
                                                                           (lizzieLet6_6QNode_Int_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet6_6QNode_Int_emitted;
  logic [1:0] lizzieLet6_6QNode_Int_done;
  assign lizzieLet6_6QNode_Int_1_d = {lizzieLet6_6QNode_Int_d[16:1],
                                      (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[0]))};
  assign lizzieLet6_6QNode_Int_2_d = {lizzieLet6_6QNode_Int_d[16:1],
                                      (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[1]))};
  assign lizzieLet6_6QNode_Int_done = (lizzieLet6_6QNode_Int_emitted | ({lizzieLet6_6QNode_Int_2_d[0],
                                                                         lizzieLet6_6QNode_Int_1_d[0]} & {lizzieLet6_6QNode_Int_2_r,
                                                                                                          lizzieLet6_6QNode_Int_1_r}));
  assign lizzieLet6_6QNode_Int_r = (& lizzieLet6_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_6QNode_Int_emitted <= (lizzieLet6_6QNode_Int_r ? 2'd0 :
                                        lizzieLet6_6QNode_Int_done);
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_6QNode_Int_2,Pointer_QTree_Int) > (lizzieLet6_6QNode_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_bufchan_d;
  logic lizzieLet6_6QNode_Int_2_bufchan_r;
  assign lizzieLet6_6QNode_Int_2_r = ((! lizzieLet6_6QNode_Int_2_bufchan_d[0]) || lizzieLet6_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNode_Int_2_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QNode_Int_2_r)
        lizzieLet6_6QNode_Int_2_bufchan_d <= lizzieLet6_6QNode_Int_2_d;
  Pointer_QTree_Int_t lizzieLet6_6QNode_Int_2_bufchan_buf;
  assign lizzieLet6_6QNode_Int_2_bufchan_r = (! lizzieLet6_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_6QNode_Int_2_argbuf_d = (lizzieLet6_6QNode_Int_2_bufchan_buf[0] ? lizzieLet6_6QNode_Int_2_bufchan_buf :
                                             lizzieLet6_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QNode_Int_2_argbuf_r && lizzieLet6_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QNode_Int_2_argbuf_r) && (! lizzieLet6_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= lizzieLet6_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_6QVal_Int,Pointer_QTree_Int) > (lizzieLet6_6QVal_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_bufchan_d;
  logic lizzieLet6_6QVal_Int_bufchan_r;
  assign lizzieLet6_6QVal_Int_r = ((! lizzieLet6_6QVal_Int_bufchan_d[0]) || lizzieLet6_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QVal_Int_r)
        lizzieLet6_6QVal_Int_bufchan_d <= lizzieLet6_6QVal_Int_d;
  Pointer_QTree_Int_t lizzieLet6_6QVal_Int_bufchan_buf;
  assign lizzieLet6_6QVal_Int_bufchan_r = (! lizzieLet6_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_6QVal_Int_1_argbuf_d = (lizzieLet6_6QVal_Int_bufchan_buf[0] ? lizzieLet6_6QVal_Int_bufchan_buf :
                                            lizzieLet6_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QVal_Int_1_argbuf_r && lizzieLet6_6QVal_Int_bufchan_buf[0]))
        lizzieLet6_6QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QVal_Int_1_argbuf_r) && (! lizzieLet6_6QVal_Int_bufchan_buf[0])))
        lizzieLet6_6QVal_Int_bufchan_buf <= lizzieLet6_6QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) > [(lizzieLet6_7QNone_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QVal_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QNode_Int,Pointer_CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet6_7QError_Int,Pointer_CTkron_kron_Int_Int_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_7_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_7_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_7QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_7QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_7QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_7QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_7QError_Int_r,
                                                              lizzieLet6_7QNode_Int_r,
                                                              lizzieLet6_7QVal_Int_r,
                                                              lizzieLet6_7QNone_Int_r}));
  assign lizzieLet6_7_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QError_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QError_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_bufchan_d;
  logic lizzieLet6_7QError_Int_bufchan_r;
  assign lizzieLet6_7QError_Int_r = ((! lizzieLet6_7QError_Int_bufchan_d[0]) || lizzieLet6_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QError_Int_r)
        lizzieLet6_7QError_Int_bufchan_d <= lizzieLet6_7QError_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QError_Int_bufchan_buf;
  assign lizzieLet6_7QError_Int_bufchan_r = (! lizzieLet6_7QError_Int_bufchan_buf[0]);
  assign lizzieLet6_7QError_Int_1_argbuf_d = (lizzieLet6_7QError_Int_bufchan_buf[0] ? lizzieLet6_7QError_Int_bufchan_buf :
                                              lizzieLet6_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QError_Int_1_argbuf_r && lizzieLet6_7QError_Int_bufchan_buf[0]))
        lizzieLet6_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QError_Int_1_argbuf_r) && (! lizzieLet6_7QError_Int_bufchan_buf[0])))
        lizzieLet6_7QError_Int_bufchan_buf <= lizzieLet6_7QError_Int_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Int_Int_Int,
      Dcon Lcall_kron_kron_Int_Int_Int3) : [(lizzieLet6_7QNode_Int,Pointer_CTkron_kron_Int_Int_Int),
                                            (lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                            (lizzieLet6_3QNode_Int_1,MyDTInt_Int_Int),
                                            (q1acQ_destruct,Pointer_QTree_Int),
                                            (lizzieLet6_6QNode_Int_1,Pointer_QTree_Int),
                                            (q2acR_destruct,Pointer_QTree_Int),
                                            (q3acS_destruct,Pointer_QTree_Int)] > (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) */
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_d = Lcall_kron_kron_Int_Int_Int3_dc((& {lizzieLet6_7QNode_Int_d[0],
                                                                                                                                                                                               lizzieLet6_5QNode_Int_1_d[0],
                                                                                                                                                                                               lizzieLet6_3QNode_Int_1_d[0],
                                                                                                                                                                                               q1acQ_destruct_d[0],
                                                                                                                                                                                               lizzieLet6_6QNode_Int_1_d[0],
                                                                                                                                                                                               q2acR_destruct_d[0],
                                                                                                                                                                                               q3acS_destruct_d[0]}), lizzieLet6_7QNode_Int_d, lizzieLet6_5QNode_Int_1_d, lizzieLet6_3QNode_Int_1_d, q1acQ_destruct_d, lizzieLet6_6QNode_Int_1_d, q2acR_destruct_d, q3acS_destruct_d);
  assign {lizzieLet6_7QNode_Int_r,
          lizzieLet6_5QNode_Int_1_r,
          lizzieLet6_3QNode_Int_1_r,
          q1acQ_destruct_r,
          lizzieLet6_6QNode_Int_1_r,
          q2acR_destruct_r,
          q3acS_destruct_r} = {7 {(lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_r && lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_d[0])}};
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3,CTkron_kron_Int_Int_Int) > (lizzieLet8_1_argbuf,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  logic lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_r;
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_r = ((! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d[0]) || lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d <= {83'd0,
                                                                                                                                                                  1'd0};
    else
      if (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_r)
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d <= lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_d;
  CTkron_kron_Int_Int_Int_t lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf;
  assign lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_r = (! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0] ? lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf :
                                  lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                    1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                      1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_buf <= lizzieLet6_7QNode_Int_1lizzieLet6_5QNode_Int_1lizzieLet6_3QNode_Int_1q1acQ_1lizzieLet6_6QNode_Int_1q2acR_1q3acS_1Lcall_kron_kron_Int_Int_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QNone_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QNone_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_bufchan_d;
  logic lizzieLet6_7QNone_Int_bufchan_r;
  assign lizzieLet6_7QNone_Int_r = ((! lizzieLet6_7QNone_Int_bufchan_d[0]) || lizzieLet6_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QNone_Int_r)
        lizzieLet6_7QNone_Int_bufchan_d <= lizzieLet6_7QNone_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QNone_Int_bufchan_buf;
  assign lizzieLet6_7QNone_Int_bufchan_r = (! lizzieLet6_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_7QNone_Int_1_argbuf_d = (lizzieLet6_7QNone_Int_bufchan_buf[0] ? lizzieLet6_7QNone_Int_bufchan_buf :
                                             lizzieLet6_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QNone_Int_1_argbuf_r && lizzieLet6_7QNone_Int_bufchan_buf[0]))
        lizzieLet6_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QNone_Int_1_argbuf_r) && (! lizzieLet6_7QNone_Int_bufchan_buf[0])))
        lizzieLet6_7QNone_Int_bufchan_buf <= lizzieLet6_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (lizzieLet6_7QVal_Int,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet6_7QVal_Int_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_bufchan_d;
  logic lizzieLet6_7QVal_Int_bufchan_r;
  assign lizzieLet6_7QVal_Int_r = ((! lizzieLet6_7QVal_Int_bufchan_d[0]) || lizzieLet6_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_7QVal_Int_r)
        lizzieLet6_7QVal_Int_bufchan_d <= lizzieLet6_7QVal_Int_d;
  Pointer_CTkron_kron_Int_Int_Int_t lizzieLet6_7QVal_Int_bufchan_buf;
  assign lizzieLet6_7QVal_Int_bufchan_r = (! lizzieLet6_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_7QVal_Int_1_argbuf_d = (lizzieLet6_7QVal_Int_bufchan_buf[0] ? lizzieLet6_7QVal_Int_bufchan_buf :
                                            lizzieLet6_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_7QVal_Int_1_argbuf_r && lizzieLet6_7QVal_Int_bufchan_buf[0]))
        lizzieLet6_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_7QVal_Int_1_argbuf_r) && (! lizzieLet6_7QVal_Int_bufchan_buf[0])))
        lizzieLet6_7QVal_Int_bufchan_buf <= lizzieLet6_7QVal_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1acN_goMux_mux,Pointer_QTree_Int) > (m1acN_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1acN_goMux_mux_bufchan_d;
  logic m1acN_goMux_mux_bufchan_r;
  assign m1acN_goMux_mux_r = ((! m1acN_goMux_mux_bufchan_d[0]) || m1acN_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acN_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1acN_goMux_mux_r)
        m1acN_goMux_mux_bufchan_d <= m1acN_goMux_mux_d;
  Pointer_QTree_Int_t m1acN_goMux_mux_bufchan_buf;
  assign m1acN_goMux_mux_bufchan_r = (! m1acN_goMux_mux_bufchan_buf[0]);
  assign m1acN_1_argbuf_d = (m1acN_goMux_mux_bufchan_buf[0] ? m1acN_goMux_mux_bufchan_buf :
                             m1acN_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1acN_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1acN_1_argbuf_r && m1acN_goMux_mux_bufchan_buf[0]))
        m1acN_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1acN_1_argbuf_r) && (! m1acN_goMux_mux_bufchan_buf[0])))
        m1acN_goMux_mux_bufchan_buf <= m1acN_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2acO_2_2,Pointer_QTree_Int) > (m2acO_2_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2acO_2_2_bufchan_d;
  logic m2acO_2_2_bufchan_r;
  assign m2acO_2_2_r = ((! m2acO_2_2_bufchan_d[0]) || m2acO_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_2_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2acO_2_2_r) m2acO_2_2_bufchan_d <= m2acO_2_2_d;
  Pointer_QTree_Int_t m2acO_2_2_bufchan_buf;
  assign m2acO_2_2_bufchan_r = (! m2acO_2_2_bufchan_buf[0]);
  assign m2acO_2_2_argbuf_d = (m2acO_2_2_bufchan_buf[0] ? m2acO_2_2_bufchan_buf :
                               m2acO_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_2_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acO_2_2_argbuf_r && m2acO_2_2_bufchan_buf[0]))
        m2acO_2_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acO_2_2_argbuf_r) && (! m2acO_2_2_bufchan_buf[0])))
        m2acO_2_2_bufchan_buf <= m2acO_2_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2acO_2_destruct,Pointer_QTree_Int) > [(m2acO_2_1,Pointer_QTree_Int),
                                                                      (m2acO_2_2,Pointer_QTree_Int)] */
  logic [1:0] m2acO_2_destruct_emitted;
  logic [1:0] m2acO_2_destruct_done;
  assign m2acO_2_1_d = {m2acO_2_destruct_d[16:1],
                        (m2acO_2_destruct_d[0] && (! m2acO_2_destruct_emitted[0]))};
  assign m2acO_2_2_d = {m2acO_2_destruct_d[16:1],
                        (m2acO_2_destruct_d[0] && (! m2acO_2_destruct_emitted[1]))};
  assign m2acO_2_destruct_done = (m2acO_2_destruct_emitted | ({m2acO_2_2_d[0],
                                                               m2acO_2_1_d[0]} & {m2acO_2_2_r,
                                                                                  m2acO_2_1_r}));
  assign m2acO_2_destruct_r = (& m2acO_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_2_destruct_emitted <= 2'd0;
    else
      m2acO_2_destruct_emitted <= (m2acO_2_destruct_r ? 2'd0 :
                                   m2acO_2_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2acO_3_2,Pointer_QTree_Int) > (m2acO_3_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2acO_3_2_bufchan_d;
  logic m2acO_3_2_bufchan_r;
  assign m2acO_3_2_r = ((! m2acO_3_2_bufchan_d[0]) || m2acO_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_3_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2acO_3_2_r) m2acO_3_2_bufchan_d <= m2acO_3_2_d;
  Pointer_QTree_Int_t m2acO_3_2_bufchan_buf;
  assign m2acO_3_2_bufchan_r = (! m2acO_3_2_bufchan_buf[0]);
  assign m2acO_3_2_argbuf_d = (m2acO_3_2_bufchan_buf[0] ? m2acO_3_2_bufchan_buf :
                               m2acO_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_3_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acO_3_2_argbuf_r && m2acO_3_2_bufchan_buf[0]))
        m2acO_3_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acO_3_2_argbuf_r) && (! m2acO_3_2_bufchan_buf[0])))
        m2acO_3_2_bufchan_buf <= m2acO_3_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2acO_3_destruct,Pointer_QTree_Int) > [(m2acO_3_1,Pointer_QTree_Int),
                                                                      (m2acO_3_2,Pointer_QTree_Int)] */
  logic [1:0] m2acO_3_destruct_emitted;
  logic [1:0] m2acO_3_destruct_done;
  assign m2acO_3_1_d = {m2acO_3_destruct_d[16:1],
                        (m2acO_3_destruct_d[0] && (! m2acO_3_destruct_emitted[0]))};
  assign m2acO_3_2_d = {m2acO_3_destruct_d[16:1],
                        (m2acO_3_destruct_d[0] && (! m2acO_3_destruct_emitted[1]))};
  assign m2acO_3_destruct_done = (m2acO_3_destruct_emitted | ({m2acO_3_2_d[0],
                                                               m2acO_3_1_d[0]} & {m2acO_3_2_r,
                                                                                  m2acO_3_1_r}));
  assign m2acO_3_destruct_r = (& m2acO_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_3_destruct_emitted <= 2'd0;
    else
      m2acO_3_destruct_emitted <= (m2acO_3_destruct_r ? 2'd0 :
                                   m2acO_3_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2acO_4_destruct,Pointer_QTree_Int) > (m2acO_4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2acO_4_destruct_bufchan_d;
  logic m2acO_4_destruct_bufchan_r;
  assign m2acO_4_destruct_r = ((! m2acO_4_destruct_bufchan_d[0]) || m2acO_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2acO_4_destruct_r)
        m2acO_4_destruct_bufchan_d <= m2acO_4_destruct_d;
  Pointer_QTree_Int_t m2acO_4_destruct_bufchan_buf;
  assign m2acO_4_destruct_bufchan_r = (! m2acO_4_destruct_bufchan_buf[0]);
  assign m2acO_4_1_argbuf_d = (m2acO_4_destruct_bufchan_buf[0] ? m2acO_4_destruct_bufchan_buf :
                               m2acO_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2acO_4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2acO_4_1_argbuf_r && m2acO_4_destruct_bufchan_buf[0]))
        m2acO_4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2acO_4_1_argbuf_r) && (! m2acO_4_destruct_bufchan_buf[0])))
        m2acO_4_destruct_bufchan_buf <= m2acO_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (macF_goMux_mux,Pointer_QTree_Int) > (macF_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t macF_goMux_mux_bufchan_d;
  logic macF_goMux_mux_bufchan_r;
  assign macF_goMux_mux_r = ((! macF_goMux_mux_bufchan_d[0]) || macF_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macF_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (macF_goMux_mux_r) macF_goMux_mux_bufchan_d <= macF_goMux_mux_d;
  Pointer_QTree_Int_t macF_goMux_mux_bufchan_buf;
  assign macF_goMux_mux_bufchan_r = (! macF_goMux_mux_bufchan_buf[0]);
  assign macF_1_argbuf_d = (macF_goMux_mux_bufchan_buf[0] ? macF_goMux_mux_bufchan_buf :
                            macF_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macF_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((macF_1_argbuf_r && macF_goMux_mux_bufchan_buf[0]))
        macF_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! macF_1_argbuf_r) && (! macF_goMux_mux_bufchan_buf[0])))
        macF_goMux_mux_bufchan_buf <= macF_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (mack_1,Pointer_QTree_Int) > (mack_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t mack_1_bufchan_d;
  logic mack_1_bufchan_r;
  assign mack_1_r = ((! mack_1_bufchan_d[0]) || mack_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mack_1_bufchan_d <= {16'd0, 1'd0};
    else if (mack_1_r) mack_1_bufchan_d <= mack_1_d;
  Pointer_QTree_Int_t mack_1_bufchan_buf;
  assign mack_1_bufchan_r = (! mack_1_bufchan_buf[0]);
  assign mack_1_argbuf_d = (mack_1_bufchan_buf[0] ? mack_1_bufchan_buf :
                            mack_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mack_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mack_1_argbuf_r && mack_1_bufchan_buf[0]))
        mack_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mack_1_argbuf_r) && (! mack_1_bufchan_buf[0])))
        mack_1_bufchan_buf <= mack_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (mack_goMux_mux,Pointer_QTree_Int) > [(mack_1,Pointer_QTree_Int),
                                                                    (mack_2,Pointer_QTree_Int)] */
  logic [1:0] mack_goMux_mux_emitted;
  logic [1:0] mack_goMux_mux_done;
  assign mack_1_d = {mack_goMux_mux_d[16:1],
                     (mack_goMux_mux_d[0] && (! mack_goMux_mux_emitted[0]))};
  assign mack_2_d = {mack_goMux_mux_d[16:1],
                     (mack_goMux_mux_d[0] && (! mack_goMux_mux_emitted[1]))};
  assign mack_goMux_mux_done = (mack_goMux_mux_emitted | ({mack_2_d[0],
                                                           mack_1_d[0]} & {mack_2_r, mack_1_r}));
  assign mack_goMux_mux_r = (& mack_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mack_goMux_mux_emitted <= 2'd0;
    else
      mack_goMux_mux_emitted <= (mack_goMux_mux_r ? 2'd0 :
                                 mack_goMux_mux_done);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_MaskQTree,
          Dcon TupGo___Pointer_QTree_Int___Pointer_MaskQTree) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Int___Pointer_MaskQTree) > [(main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13,Go),
                                                                                                                                                                                (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1,Pointer_QTree_Int),
                                                                                                                                                                                (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1,Pointer_MaskQTree)] */
  logic [2:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted;
  logic [2:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[0]));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_d = {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[16:1],
                                                                               (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[1]))};
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_d = {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[32:17],
                                                                                 (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted[2]))};
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted | ({main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_d[0],
                                                                                                                                                       main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_d[0],
                                                                                                                                                       main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_d[0]} & {main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_r,
                                                                                                                                                                                                                                main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_r,
                                                                                                                                                                                                                                main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_r}));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r = (& main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted <= 3'd0;
    else
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_emitted <= (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_r ? 3'd0 :
                                                                               main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTree_1_done);
  
  /* fork (Ty Go) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13,Go) > [(go_13_1,Go),
                                                                                       (go_13_2,Go)] */
  logic [1:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted;
  logic [1:0] main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_done;
  assign go_13_1_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted[0]));
  assign go_13_2_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_d[0] && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted[1]));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_done = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted | ({go_13_2_d[0],
                                                                                                                                                             go_13_1_d[0]} & {go_13_2_r,
                                                                                                                                                                              go_13_1_r}));
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_r = (& main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted <= 2'd0;
    else
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_emitted <= (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_r ? 2'd0 :
                                                                                  main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreego_13_done);
  
  /* buf (Ty Pointer_QTree_Int) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1,Pointer_QTree_Int) > (mack_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_r;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_r = ((! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d[0]) || main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d <= {16'd0,
                                                                                     1'd0};
    else
      if (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_r)
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_d;
  Pointer_QTree_Int_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_r = (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf[0]);
  assign mack_1_1_argbuf_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf[0] ? main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf :
                              main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf <= {16'd0,
                                                                                       1'd0};
    else
      if ((mack_1_1_argbuf_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf[0]))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
      else if (((! mack_1_1_argbuf_r) && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf[0])))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_buf <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemack_1_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1,Pointer_MaskQTree) > (mskacl_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d;
  logic main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_r;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_r = ((! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d[0]) || main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d <= {16'd0,
                                                                                       1'd0};
    else
      if (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_r)
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_d;
  Pointer_MaskQTree_t main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf;
  assign main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_r = (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf[0]);
  assign mskacl_1_1_argbuf_d = (main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf[0] ? main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf :
                                main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
    else
      if ((mskacl_1_1_argbuf_r && main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf[0]))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
      else if (((! mskacl_1_1_argbuf_r) && (! main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf[0])))
        main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_buf <= main_mask_IntTupGo___Pointer_QTree_Int___Pointer_MaskQTreemskacl_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (main_mask_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t main_mask_Int_resbuf_bufchan_d;
  logic main_mask_Int_resbuf_bufchan_r;
  assign main_mask_Int_resbuf_r = ((! main_mask_Int_resbuf_bufchan_d[0]) || main_mask_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (main_mask_Int_resbuf_r)
        main_mask_Int_resbuf_bufchan_d <= main_mask_Int_resbuf_d;
  Pointer_QTree_Int_t main_mask_Int_resbuf_bufchan_buf;
  assign main_mask_Int_resbuf_bufchan_r = (! main_mask_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (main_mask_Int_resbuf_bufchan_buf[0] ? main_mask_Int_resbuf_bufchan_buf :
                            main_mask_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && main_mask_Int_resbuf_bufchan_buf[0]))
        main_mask_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! main_mask_Int_resbuf_bufchan_buf[0])))
        main_mask_Int_resbuf_bufchan_buf <= main_mask_Int_resbuf_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int) > [(map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14,Go),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1,Int),
                                                                                                                                                                                                                                                   (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1,Pointer_QTree_Int)] */
  logic [4:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted ;
  logic [4:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [0]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [1]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [2]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_d  = {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [32:1],
                                                                                                               (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [3]))};
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_d  = {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [48:33],
                                                                                                              (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted [4]))};
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  | ({\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_d [0],
                                                                                                                                                                                                                     \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_d [0]} & {\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_r ,
                                                                                                                                                                                                                                                                                                                             \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_r }));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  = (& \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  <= 5'd0;
    else
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_emitted  <= (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_r  ? 5'd0 :
                                                                                                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Int_1_done );
  
  /* buf (Ty MyDTInt_Int_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1,MyDTInt_Int_Int) > (gacD_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_d ;
  MyDTInt_Int_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf [0]);
  assign gacD_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf  :
                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf  <= 1'd0;
    else
      if ((gacD_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf  <= 1'd0;
      else if (((! gacD_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntgacD_1_bufchan_d ;
  
  /* fork (Ty Go) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14,Go) > [(go_14_1,Go),
                                                                                                                    (go_14_2,Go)] */
  logic [1:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted ;
  logic [1:0] \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_done ;
  assign go_14_1_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted [0]));
  assign go_14_2_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_d [0] && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted [1]));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_done  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted  | ({go_14_2_d[0],
                                                                                                                                                                                                                           go_14_1_d[0]} & {go_14_2_r,
                                                                                                                                                                                                                                            go_14_1_r}));
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_r  = (& \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted  <= 2'd0;
    else
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_emitted  <= (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_r  ? 2'd0 :
                                                                                                                 \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intgo_14_done );
  
  /* buf (Ty MyDTInt_Bool) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1,MyDTInt_Bool) > (isZacC_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_d ;
  MyDTInt_Bool_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf [0]);
  assign isZacC_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf  :
                                \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacC_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf  <= 1'd0;
      else if (((! isZacC_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntisZacC_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1,Pointer_QTree_Int) > (macF_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d  <= {16'd0,
                                                                                                                    1'd0};
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_d ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf [0]);
  assign macF_1_1_argbuf_d = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf  :
                              \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf  <= {16'd0,
                                                                                                                      1'd0};
    else
      if ((macF_1_1_argbuf_r && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf  <= {16'd0,
                                                                                                                        1'd0};
      else if (((! macF_1_1_argbuf_r) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_IntmacF_1_bufchan_d ;
  
  /* buf (Ty Int) : (map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1,Int) > (v'acE_1_1_argbuf,Int) */
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d ;
  logic \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_r ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_r  = ((! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d [0]) || \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d  <= {32'd0,
                                                                                                                     1'd0};
    else
      if (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_r )
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_d ;
  Int_t \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf ;
  assign \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_r  = (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf [0]);
  assign \v'acE_1_1_argbuf_d  = (\map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf [0] ? \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf  :
                                 \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf  <= {32'd0,
                                                                                                                       1'd0};
    else
      if ((\v'acE_1_1_argbuf_r  && \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf [0]))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf  <= {32'd0,
                                                                                                                         1'd0};
      else if (((! \v'acE_1_1_argbuf_r ) && (! \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf [0])))
        \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_buf  <= \map''_map''_Int_Int_IntTupGo___MyDTInt_Bool___MyDTInt_Int_Int___Int___Pointer_QTree_Intv'acE_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (map''_map''_Int_Int_Int_resbuf,Pointer_QTree_Int) > (lizzieLet11_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_bufchan_d ;
  logic \map''_map''_Int_Int_Int_resbuf_bufchan_r ;
  assign \map''_map''_Int_Int_Int_resbuf_r  = ((! \map''_map''_Int_Int_Int_resbuf_bufchan_d [0]) || \map''_map''_Int_Int_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\map''_map''_Int_Int_Int_resbuf_r )
        \map''_map''_Int_Int_Int_resbuf_bufchan_d  <= \map''_map''_Int_Int_Int_resbuf_d ;
  Pointer_QTree_Int_t \map''_map''_Int_Int_Int_resbuf_bufchan_buf ;
  assign \map''_map''_Int_Int_Int_resbuf_bufchan_r  = (! \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0]);
  assign lizzieLet11_1_argbuf_d = (\map''_map''_Int_Int_Int_resbuf_bufchan_buf [0] ? \map''_map''_Int_Int_Int_resbuf_bufchan_buf  :
                                   \map''_map''_Int_Int_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0]))
        \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! \map''_map''_Int_Int_Int_resbuf_bufchan_buf [0])))
        \map''_map''_Int_Int_Int_resbuf_bufchan_buf  <= \map''_map''_Int_Int_Int_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (mskacl_goMux_mux,Pointer_MaskQTree) > (mskacl_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t mskacl_goMux_mux_bufchan_d;
  logic mskacl_goMux_mux_bufchan_r;
  assign mskacl_goMux_mux_r = ((! mskacl_goMux_mux_bufchan_d[0]) || mskacl_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mskacl_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (mskacl_goMux_mux_r)
        mskacl_goMux_mux_bufchan_d <= mskacl_goMux_mux_d;
  Pointer_MaskQTree_t mskacl_goMux_mux_bufchan_buf;
  assign mskacl_goMux_mux_bufchan_r = (! mskacl_goMux_mux_bufchan_buf[0]);
  assign mskacl_1_argbuf_d = (mskacl_goMux_mux_bufchan_buf[0] ? mskacl_goMux_mux_bufchan_buf :
                              mskacl_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mskacl_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mskacl_1_argbuf_r && mskacl_goMux_mux_bufchan_buf[0]))
        mskacl_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mskacl_1_argbuf_r) && (! mskacl_goMux_mux_bufchan_buf[0])))
        mskacl_goMux_mux_bufchan_buf <= mskacl_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1acH_3_destruct,Pointer_QTree_Int) > (q1acH_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1acH_3_destruct_bufchan_d;
  logic q1acH_3_destruct_bufchan_r;
  assign q1acH_3_destruct_r = ((! q1acH_3_destruct_bufchan_d[0]) || q1acH_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acH_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acH_3_destruct_r)
        q1acH_3_destruct_bufchan_d <= q1acH_3_destruct_d;
  Pointer_QTree_Int_t q1acH_3_destruct_bufchan_buf;
  assign q1acH_3_destruct_bufchan_r = (! q1acH_3_destruct_bufchan_buf[0]);
  assign q1acH_3_1_argbuf_d = (q1acH_3_destruct_bufchan_buf[0] ? q1acH_3_destruct_bufchan_buf :
                               q1acH_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acH_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acH_3_1_argbuf_r && q1acH_3_destruct_bufchan_buf[0]))
        q1acH_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acH_3_1_argbuf_r) && (! q1acH_3_destruct_bufchan_buf[0])))
        q1acH_3_destruct_bufchan_buf <= q1acH_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1acQ_3_destruct,Pointer_QTree_Int) > (q1acQ_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1acQ_3_destruct_bufchan_d;
  logic q1acQ_3_destruct_bufchan_r;
  assign q1acQ_3_destruct_r = ((! q1acQ_3_destruct_bufchan_d[0]) || q1acQ_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acQ_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acQ_3_destruct_r)
        q1acQ_3_destruct_bufchan_d <= q1acQ_3_destruct_d;
  Pointer_QTree_Int_t q1acQ_3_destruct_bufchan_buf;
  assign q1acQ_3_destruct_bufchan_r = (! q1acQ_3_destruct_bufchan_buf[0]);
  assign q1acQ_3_1_argbuf_d = (q1acQ_3_destruct_bufchan_buf[0] ? q1acQ_3_destruct_bufchan_buf :
                               q1acQ_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acQ_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acQ_3_1_argbuf_r && q1acQ_3_destruct_bufchan_buf[0]))
        q1acQ_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acQ_3_1_argbuf_r) && (! q1acQ_3_destruct_bufchan_buf[0])))
        q1acQ_3_destruct_bufchan_buf <= q1acQ_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1acV_destruct,Pointer_QTree_Int) > (q1acV_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1acV_destruct_bufchan_d;
  logic q1acV_destruct_bufchan_r;
  assign q1acV_destruct_r = ((! q1acV_destruct_bufchan_d[0]) || q1acV_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acV_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acV_destruct_r) q1acV_destruct_bufchan_d <= q1acV_destruct_d;
  Pointer_QTree_Int_t q1acV_destruct_bufchan_buf;
  assign q1acV_destruct_bufchan_r = (! q1acV_destruct_bufchan_buf[0]);
  assign q1acV_1_argbuf_d = (q1acV_destruct_bufchan_buf[0] ? q1acV_destruct_bufchan_buf :
                             q1acV_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acV_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acV_1_argbuf_r && q1acV_destruct_bufchan_buf[0]))
        q1acV_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acV_1_argbuf_r) && (! q1acV_destruct_bufchan_buf[0])))
        q1acV_destruct_bufchan_buf <= q1acV_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1acm_3_destruct,Pointer_MaskQTree) > (q1acm_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1acm_3_destruct_bufchan_d;
  logic q1acm_3_destruct_bufchan_r;
  assign q1acm_3_destruct_r = ((! q1acm_3_destruct_bufchan_d[0]) || q1acm_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acm_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acm_3_destruct_r)
        q1acm_3_destruct_bufchan_d <= q1acm_3_destruct_d;
  Pointer_MaskQTree_t q1acm_3_destruct_bufchan_buf;
  assign q1acm_3_destruct_bufchan_r = (! q1acm_3_destruct_bufchan_buf[0]);
  assign q1acm_3_1_argbuf_d = (q1acm_3_destruct_bufchan_buf[0] ? q1acm_3_destruct_bufchan_buf :
                               q1acm_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acm_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acm_3_1_argbuf_r && q1acm_3_destruct_bufchan_buf[0]))
        q1acm_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acm_3_1_argbuf_r) && (! q1acm_3_destruct_bufchan_buf[0])))
        q1acm_3_destruct_bufchan_buf <= q1acm_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2acI_2_destruct,Pointer_QTree_Int) > (q2acI_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2acI_2_destruct_bufchan_d;
  logic q2acI_2_destruct_bufchan_r;
  assign q2acI_2_destruct_r = ((! q2acI_2_destruct_bufchan_d[0]) || q2acI_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acI_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acI_2_destruct_r)
        q2acI_2_destruct_bufchan_d <= q2acI_2_destruct_d;
  Pointer_QTree_Int_t q2acI_2_destruct_bufchan_buf;
  assign q2acI_2_destruct_bufchan_r = (! q2acI_2_destruct_bufchan_buf[0]);
  assign q2acI_2_1_argbuf_d = (q2acI_2_destruct_bufchan_buf[0] ? q2acI_2_destruct_bufchan_buf :
                               q2acI_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acI_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acI_2_1_argbuf_r && q2acI_2_destruct_bufchan_buf[0]))
        q2acI_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acI_2_1_argbuf_r) && (! q2acI_2_destruct_bufchan_buf[0])))
        q2acI_2_destruct_bufchan_buf <= q2acI_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2acR_2_destruct,Pointer_QTree_Int) > (q2acR_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2acR_2_destruct_bufchan_d;
  logic q2acR_2_destruct_bufchan_r;
  assign q2acR_2_destruct_r = ((! q2acR_2_destruct_bufchan_d[0]) || q2acR_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acR_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acR_2_destruct_r)
        q2acR_2_destruct_bufchan_d <= q2acR_2_destruct_d;
  Pointer_QTree_Int_t q2acR_2_destruct_bufchan_buf;
  assign q2acR_2_destruct_bufchan_r = (! q2acR_2_destruct_bufchan_buf[0]);
  assign q2acR_2_1_argbuf_d = (q2acR_2_destruct_bufchan_buf[0] ? q2acR_2_destruct_bufchan_buf :
                               q2acR_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acR_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acR_2_1_argbuf_r && q2acR_2_destruct_bufchan_buf[0]))
        q2acR_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acR_2_1_argbuf_r) && (! q2acR_2_destruct_bufchan_buf[0])))
        q2acR_2_destruct_bufchan_buf <= q2acR_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2acW_1_destruct,Pointer_QTree_Int) > (q2acW_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2acW_1_destruct_bufchan_d;
  logic q2acW_1_destruct_bufchan_r;
  assign q2acW_1_destruct_r = ((! q2acW_1_destruct_bufchan_d[0]) || q2acW_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acW_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acW_1_destruct_r)
        q2acW_1_destruct_bufchan_d <= q2acW_1_destruct_d;
  Pointer_QTree_Int_t q2acW_1_destruct_bufchan_buf;
  assign q2acW_1_destruct_bufchan_r = (! q2acW_1_destruct_bufchan_buf[0]);
  assign q2acW_1_1_argbuf_d = (q2acW_1_destruct_bufchan_buf[0] ? q2acW_1_destruct_bufchan_buf :
                               q2acW_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acW_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acW_1_1_argbuf_r && q2acW_1_destruct_bufchan_buf[0]))
        q2acW_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acW_1_1_argbuf_r) && (! q2acW_1_destruct_bufchan_buf[0])))
        q2acW_1_destruct_bufchan_buf <= q2acW_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2acn_2_destruct,Pointer_MaskQTree) > (q2acn_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2acn_2_destruct_bufchan_d;
  logic q2acn_2_destruct_bufchan_r;
  assign q2acn_2_destruct_r = ((! q2acn_2_destruct_bufchan_d[0]) || q2acn_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acn_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acn_2_destruct_r)
        q2acn_2_destruct_bufchan_d <= q2acn_2_destruct_d;
  Pointer_MaskQTree_t q2acn_2_destruct_bufchan_buf;
  assign q2acn_2_destruct_bufchan_r = (! q2acn_2_destruct_bufchan_buf[0]);
  assign q2acn_2_1_argbuf_d = (q2acn_2_destruct_bufchan_buf[0] ? q2acn_2_destruct_bufchan_buf :
                               q2acn_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acn_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acn_2_1_argbuf_r && q2acn_2_destruct_bufchan_buf[0]))
        q2acn_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acn_2_1_argbuf_r) && (! q2acn_2_destruct_bufchan_buf[0])))
        q2acn_2_destruct_bufchan_buf <= q2acn_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3acJ_1_destruct,Pointer_QTree_Int) > (q3acJ_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3acJ_1_destruct_bufchan_d;
  logic q3acJ_1_destruct_bufchan_r;
  assign q3acJ_1_destruct_r = ((! q3acJ_1_destruct_bufchan_d[0]) || q3acJ_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acJ_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acJ_1_destruct_r)
        q3acJ_1_destruct_bufchan_d <= q3acJ_1_destruct_d;
  Pointer_QTree_Int_t q3acJ_1_destruct_bufchan_buf;
  assign q3acJ_1_destruct_bufchan_r = (! q3acJ_1_destruct_bufchan_buf[0]);
  assign q3acJ_1_1_argbuf_d = (q3acJ_1_destruct_bufchan_buf[0] ? q3acJ_1_destruct_bufchan_buf :
                               q3acJ_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acJ_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acJ_1_1_argbuf_r && q3acJ_1_destruct_bufchan_buf[0]))
        q3acJ_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acJ_1_1_argbuf_r) && (! q3acJ_1_destruct_bufchan_buf[0])))
        q3acJ_1_destruct_bufchan_buf <= q3acJ_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3acS_1_destruct,Pointer_QTree_Int) > (q3acS_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3acS_1_destruct_bufchan_d;
  logic q3acS_1_destruct_bufchan_r;
  assign q3acS_1_destruct_r = ((! q3acS_1_destruct_bufchan_d[0]) || q3acS_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acS_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acS_1_destruct_r)
        q3acS_1_destruct_bufchan_d <= q3acS_1_destruct_d;
  Pointer_QTree_Int_t q3acS_1_destruct_bufchan_buf;
  assign q3acS_1_destruct_bufchan_r = (! q3acS_1_destruct_bufchan_buf[0]);
  assign q3acS_1_1_argbuf_d = (q3acS_1_destruct_bufchan_buf[0] ? q3acS_1_destruct_bufchan_buf :
                               q3acS_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acS_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acS_1_1_argbuf_r && q3acS_1_destruct_bufchan_buf[0]))
        q3acS_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acS_1_1_argbuf_r) && (! q3acS_1_destruct_bufchan_buf[0])))
        q3acS_1_destruct_bufchan_buf <= q3acS_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3acX_2_destruct,Pointer_QTree_Int) > (q3acX_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3acX_2_destruct_bufchan_d;
  logic q3acX_2_destruct_bufchan_r;
  assign q3acX_2_destruct_r = ((! q3acX_2_destruct_bufchan_d[0]) || q3acX_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acX_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acX_2_destruct_r)
        q3acX_2_destruct_bufchan_d <= q3acX_2_destruct_d;
  Pointer_QTree_Int_t q3acX_2_destruct_bufchan_buf;
  assign q3acX_2_destruct_bufchan_r = (! q3acX_2_destruct_bufchan_buf[0]);
  assign q3acX_2_1_argbuf_d = (q3acX_2_destruct_bufchan_buf[0] ? q3acX_2_destruct_bufchan_buf :
                               q3acX_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acX_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acX_2_1_argbuf_r && q3acX_2_destruct_bufchan_buf[0]))
        q3acX_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acX_2_1_argbuf_r) && (! q3acX_2_destruct_bufchan_buf[0])))
        q3acX_2_destruct_bufchan_buf <= q3acX_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3aco_1_destruct,Pointer_MaskQTree) > (q3aco_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3aco_1_destruct_bufchan_d;
  logic q3aco_1_destruct_bufchan_r;
  assign q3aco_1_destruct_r = ((! q3aco_1_destruct_bufchan_d[0]) || q3aco_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aco_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aco_1_destruct_r)
        q3aco_1_destruct_bufchan_d <= q3aco_1_destruct_d;
  Pointer_MaskQTree_t q3aco_1_destruct_bufchan_buf;
  assign q3aco_1_destruct_bufchan_r = (! q3aco_1_destruct_bufchan_buf[0]);
  assign q3aco_1_1_argbuf_d = (q3aco_1_destruct_bufchan_buf[0] ? q3aco_1_destruct_bufchan_buf :
                               q3aco_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aco_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aco_1_1_argbuf_r && q3aco_1_destruct_bufchan_buf[0]))
        q3aco_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aco_1_1_argbuf_r) && (! q3aco_1_destruct_bufchan_buf[0])))
        q3aco_1_destruct_bufchan_buf <= q3aco_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4acK_destruct,Pointer_QTree_Int) > (q4acK_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4acK_destruct_bufchan_d;
  logic q4acK_destruct_bufchan_r;
  assign q4acK_destruct_r = ((! q4acK_destruct_bufchan_d[0]) || q4acK_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acK_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acK_destruct_r) q4acK_destruct_bufchan_d <= q4acK_destruct_d;
  Pointer_QTree_Int_t q4acK_destruct_bufchan_buf;
  assign q4acK_destruct_bufchan_r = (! q4acK_destruct_bufchan_buf[0]);
  assign q4acK_1_argbuf_d = (q4acK_destruct_bufchan_buf[0] ? q4acK_destruct_bufchan_buf :
                             q4acK_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acK_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acK_1_argbuf_r && q4acK_destruct_bufchan_buf[0]))
        q4acK_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acK_1_argbuf_r) && (! q4acK_destruct_bufchan_buf[0])))
        q4acK_destruct_bufchan_buf <= q4acK_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4acT_destruct,Pointer_QTree_Int) > (q4acT_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4acT_destruct_bufchan_d;
  logic q4acT_destruct_bufchan_r;
  assign q4acT_destruct_r = ((! q4acT_destruct_bufchan_d[0]) || q4acT_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acT_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acT_destruct_r) q4acT_destruct_bufchan_d <= q4acT_destruct_d;
  Pointer_QTree_Int_t q4acT_destruct_bufchan_buf;
  assign q4acT_destruct_bufchan_r = (! q4acT_destruct_bufchan_buf[0]);
  assign q4acT_1_argbuf_d = (q4acT_destruct_bufchan_buf[0] ? q4acT_destruct_bufchan_buf :
                             q4acT_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acT_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acT_1_argbuf_r && q4acT_destruct_bufchan_buf[0]))
        q4acT_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acT_1_argbuf_r) && (! q4acT_destruct_bufchan_buf[0])))
        q4acT_destruct_bufchan_buf <= q4acT_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4acY_3_destruct,Pointer_QTree_Int) > (q4acY_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4acY_3_destruct_bufchan_d;
  logic q4acY_3_destruct_bufchan_r;
  assign q4acY_3_destruct_r = ((! q4acY_3_destruct_bufchan_d[0]) || q4acY_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acY_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acY_3_destruct_r)
        q4acY_3_destruct_bufchan_d <= q4acY_3_destruct_d;
  Pointer_QTree_Int_t q4acY_3_destruct_bufchan_buf;
  assign q4acY_3_destruct_bufchan_r = (! q4acY_3_destruct_bufchan_buf[0]);
  assign q4acY_3_1_argbuf_d = (q4acY_3_destruct_bufchan_buf[0] ? q4acY_3_destruct_bufchan_buf :
                               q4acY_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acY_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acY_3_1_argbuf_r && q4acY_3_destruct_bufchan_buf[0]))
        q4acY_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acY_3_1_argbuf_r) && (! q4acY_3_destruct_bufchan_buf[0])))
        q4acY_3_destruct_bufchan_buf <= q4acY_3_destruct_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int) > (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) */
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                             1'd0};
    else
      if (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf :
                                                           readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                               1'd0};
    else
      if ((readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
      else if (((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) > [(lizzieLet26_1,CT$wnnz_Int),
                                                                                      (lizzieLet26_2,CT$wnnz_Int),
                                                                                      (lizzieLet26_3,CT$wnnz_Int),
                                                                                      (lizzieLet26_4,CT$wnnz_Int)] */
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet26_1_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet26_2_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet26_3_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet26_4_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet26_4_d[0],
                                                                                                                       lizzieLet26_3_d[0],
                                                                                                                       lizzieLet26_2_d[0],
                                                                                                                       lizzieLet26_1_d[0]} & {lizzieLet26_4_r,
                                                                                                                                              lizzieLet26_3_r,
                                                                                                                                              lizzieLet26_2_r,
                                                                                                                                              lizzieLet26_1_r}));
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTkron_kron_Int_Int_Int) : (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf,CTkron_kron_Int_Int_Int) > (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTkron_kron_Int_Int_Int) */
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r = ((! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d <= {83'd0,
                                                                           1'd0};
    else
      if (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_r)
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_d;
  CTkron_kron_Int_Int_Int_t readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d = (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf :
                                                                         readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= {83'd0,
                                                                             1'd0};
    else
      if ((readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r && readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= {83'd0,
                                                                               1'd0};
      else if (((! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CTkron_kron_Int_Int_Int) : (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTkron_kron_Int_Int_Int) > [(lizzieLet30_1,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet30_2,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet30_3,CTkron_kron_Int_Int_Int),
                                                                                                                            (lizzieLet30_4,CTkron_kron_Int_Int_Int)] */
  logic [3:0] readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet30_1_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet30_2_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet30_3_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet30_4_d = {readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done = (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet30_4_d[0],
                                                                                                                                                   lizzieLet30_3_d[0],
                                                                                                                                                   lizzieLet30_2_d[0],
                                                                                                                                                   lizzieLet30_1_d[0]} & {lizzieLet30_4_r,
                                                                                                                                                                          lizzieLet30_3_r,
                                                                                                                                                                          lizzieLet30_2_r,
                                                                                                                                                                          lizzieLet30_1_r}));
  assign readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                                             readPointer_CTkron_kron_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_mask_Int) : (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf,CTmain_mask_Int) > (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb,CTmain_mask_Int) */
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r = ((! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d <= {115'd0,
                                                                   1'd0};
    else
      if (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_r)
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_d;
  CTmain_mask_Int_t readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf :
                                                                 readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                     1'd0};
    else
      if ((readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r && readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0,
                                                                       1'd0};
      else if (((! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTmain_mask_Int) : (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb,CTmain_mask_Int) > [(lizzieLet35_1,CTmain_mask_Int),
                                                                                                    (lizzieLet35_2,CTmain_mask_Int),
                                                                                                    (lizzieLet35_3,CTmain_mask_Int),
                                                                                                    (lizzieLet35_4,CTmain_mask_Int)] */
  logic [3:0] readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet35_1_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet35_2_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet35_3_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet35_4_d = {readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet35_4_d[0],
                                                                                                                                   lizzieLet35_3_d[0],
                                                                                                                                   lizzieLet35_2_d[0],
                                                                                                                                   lizzieLet35_1_d[0]} & {lizzieLet35_4_r,
                                                                                                                                                          lizzieLet35_3_r,
                                                                                                                                                          lizzieLet35_2_r,
                                                                                                                                                          lizzieLet35_1_r}));
  assign readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                                     readPointer_CTmain_mask_Intscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty CTmap''_map''_Int_Int_Int) : (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf,CTmap''_map''_Int_Int_Int) > (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb,CTmap''_map''_Int_Int_Int) */
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d ;
  logic \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r ;
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r  = ((! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d [0]) || \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d  <= {99'd0,
                                                                               1'd0};
    else
      if (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_r )
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d  <= \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_d ;
  \CTmap''_map''_Int_Int_Int_t  \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_r  = (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d  = (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0] ? \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  :
                                                                             \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= {99'd0,
                                                                                 1'd0};
    else
      if ((\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  && \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= {99'd0,
                                                                                   1'd0};
      else if (((! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r ) && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_buf  <= \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmap''_map''_Int_Int_Int) : (readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb,CTmap''_map''_Int_Int_Int) > [(lizzieLet40_1,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet40_2,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet40_3,CTmap''_map''_Int_Int_Int),
                                                                                                                                  (lizzieLet40_4,CTmap''_map''_Int_Int_Int)] */
  logic [3:0] \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done ;
  assign lizzieLet40_1_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet40_2_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet40_3_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet40_4_d = {\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done  = (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  | ({lizzieLet40_4_d[0],
                                                                                                                                                           lizzieLet40_3_d[0],
                                                                                                                                                           lizzieLet40_2_d[0],
                                                                                                                                                           lizzieLet40_1_d[0]} & {lizzieLet40_4_r,
                                                                                                                                                                                  lizzieLet40_3_r,
                                                                                                                                                                                  lizzieLet40_2_r,
                                                                                                                                                                                  lizzieLet40_1_r}));
  assign \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  = (& \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_emitted  <= (\readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_r  ? 4'd0 :
                                                                                 \readPointer_CTmap''_map''_Int_Int_Intscfarg_0_3_1_argbuf_rwb_done );
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreemskacl_1_argbuf,MaskQTree) > (readPointer_MaskQTreemskacl_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreemskacl_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreemskacl_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreemskacl_1_argbuf_r = ((! readPointer_MaskQTreemskacl_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreemskacl_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacl_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreemskacl_1_argbuf_r)
        readPointer_MaskQTreemskacl_1_argbuf_bufchan_d <= readPointer_MaskQTreemskacl_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreemskacl_1_argbuf_bufchan_r = (! readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreemskacl_1_argbuf_rwb_d = (readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf :
                                                       readPointer_MaskQTreemskacl_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreemskacl_1_argbuf_rwb_r && readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreemskacl_1_argbuf_rwb_r) && (! readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreemskacl_1_argbuf_bufchan_buf <= readPointer_MaskQTreemskacl_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreemskacl_1_argbuf_rwb,MaskQTree) > [(lizzieLet10_1_1,MaskQTree),
                                                                              (lizzieLet10_1_2,MaskQTree),
                                                                              (lizzieLet10_1_3,MaskQTree),
                                                                              (lizzieLet10_1_4,MaskQTree),
                                                                              (lizzieLet10_1_5,MaskQTree),
                                                                              (lizzieLet10_1_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreemskacl_1_argbuf_rwb_done;
  assign lizzieLet10_1_1_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet10_1_2_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet10_1_3_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet10_1_4_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet10_1_5_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet10_1_6_d = {readPointer_MaskQTreemskacl_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemskacl_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreemskacl_1_argbuf_rwb_done = (readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted | ({lizzieLet10_1_6_d[0],
                                                                                                               lizzieLet10_1_5_d[0],
                                                                                                               lizzieLet10_1_4_d[0],
                                                                                                               lizzieLet10_1_3_d[0],
                                                                                                               lizzieLet10_1_2_d[0],
                                                                                                               lizzieLet10_1_1_d[0]} & {lizzieLet10_1_6_r,
                                                                                                                                        lizzieLet10_1_5_r,
                                                                                                                                        lizzieLet10_1_4_r,
                                                                                                                                        lizzieLet10_1_3_r,
                                                                                                                                        lizzieLet10_1_2_r,
                                                                                                                                        lizzieLet10_1_1_r}));
  assign readPointer_MaskQTreemskacl_1_argbuf_rwb_r = (& readPointer_MaskQTreemskacl_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreemskacl_1_argbuf_rwb_emitted <= (readPointer_MaskQTreemskacl_1_argbuf_rwb_r ? 6'd0 :
                                                           readPointer_MaskQTreemskacl_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1acN_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1acN_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1acN_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1acN_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1acN_1_argbuf_r = ((! readPointer_QTree_Intm1acN_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1acN_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1acN_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1acN_1_argbuf_r)
        readPointer_QTree_Intm1acN_1_argbuf_bufchan_d <= readPointer_QTree_Intm1acN_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1acN_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1acN_1_argbuf_rwb_d = (readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1acN_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1acN_1_argbuf_rwb_r && readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1acN_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1acN_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1acN_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1acN_1_argbuf_rwb,QTree_Int) > [(lizzieLet6_1,QTree_Int),
                                                                             (lizzieLet6_2,QTree_Int),
                                                                             (lizzieLet6_3,QTree_Int),
                                                                             (lizzieLet6_4,QTree_Int),
                                                                             (lizzieLet6_5,QTree_Int),
                                                                             (lizzieLet6_6,QTree_Int),
                                                                             (lizzieLet6_7,QTree_Int)] */
  logic [6:0] readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Intm1acN_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet6_7_d = {readPointer_QTree_Intm1acN_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm1acN_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Intm1acN_1_argbuf_rwb_done = (readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted | ({lizzieLet6_7_d[0],
                                                                                                             lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_7_r,
                                                                                                                                   lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_Intm1acN_1_argbuf_rwb_r = (& readPointer_QTree_Intm1acN_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Intm1acN_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1acN_1_argbuf_rwb_r ? 7'd0 :
                                                          readPointer_QTree_Intm1acN_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntmacF_1_argbuf,QTree_Int) > (readPointer_QTree_IntmacF_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntmacF_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntmacF_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntmacF_1_argbuf_r = ((! readPointer_QTree_IntmacF_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntmacF_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacF_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntmacF_1_argbuf_r)
        readPointer_QTree_IntmacF_1_argbuf_bufchan_d <= readPointer_QTree_IntmacF_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntmacF_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntmacF_1_argbuf_bufchan_r = (! readPointer_QTree_IntmacF_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntmacF_1_argbuf_rwb_d = (readPointer_QTree_IntmacF_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntmacF_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_IntmacF_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacF_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntmacF_1_argbuf_rwb_r && readPointer_QTree_IntmacF_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntmacF_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntmacF_1_argbuf_rwb_r) && (! readPointer_QTree_IntmacF_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntmacF_1_argbuf_bufchan_buf <= readPointer_QTree_IntmacF_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntmacF_1_argbuf_rwb,QTree_Int) > [(lizzieLet17_1,QTree_Int),
                                                                            (lizzieLet17_2,QTree_Int),
                                                                            (lizzieLet17_3,QTree_Int),
                                                                            (lizzieLet17_4,QTree_Int),
                                                                            (lizzieLet17_5,QTree_Int),
                                                                            (lizzieLet17_6,QTree_Int),
                                                                            (lizzieLet17_7,QTree_Int)] */
  logic [6:0] readPointer_QTree_IntmacF_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_IntmacF_1_argbuf_rwb_done;
  assign lizzieLet17_1_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet17_2_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet17_3_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet17_4_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet17_5_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet17_6_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet17_7_d = {readPointer_QTree_IntmacF_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_IntmacF_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntmacF_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_IntmacF_1_argbuf_rwb_done = (readPointer_QTree_IntmacF_1_argbuf_rwb_emitted | ({lizzieLet17_7_d[0],
                                                                                                           lizzieLet17_6_d[0],
                                                                                                           lizzieLet17_5_d[0],
                                                                                                           lizzieLet17_4_d[0],
                                                                                                           lizzieLet17_3_d[0],
                                                                                                           lizzieLet17_2_d[0],
                                                                                                           lizzieLet17_1_d[0]} & {lizzieLet17_7_r,
                                                                                                                                  lizzieLet17_6_r,
                                                                                                                                  lizzieLet17_5_r,
                                                                                                                                  lizzieLet17_4_r,
                                                                                                                                  lizzieLet17_3_r,
                                                                                                                                  lizzieLet17_2_r,
                                                                                                                                  lizzieLet17_1_r}));
  assign readPointer_QTree_IntmacF_1_argbuf_rwb_r = (& readPointer_QTree_IntmacF_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntmacF_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_IntmacF_1_argbuf_rwb_emitted <= (readPointer_QTree_IntmacF_1_argbuf_rwb_r ? 7'd0 :
                                                         readPointer_QTree_IntmacF_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intmack_1_argbuf,QTree_Int) > (readPointer_QTree_Intmack_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intmack_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intmack_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intmack_1_argbuf_r = ((! readPointer_QTree_Intmack_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intmack_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intmack_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intmack_1_argbuf_r)
        readPointer_QTree_Intmack_1_argbuf_bufchan_d <= readPointer_QTree_Intmack_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intmack_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intmack_1_argbuf_bufchan_r = (! readPointer_QTree_Intmack_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intmack_1_argbuf_rwb_d = (readPointer_QTree_Intmack_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intmack_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_Intmack_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intmack_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intmack_1_argbuf_rwb_r && readPointer_QTree_Intmack_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intmack_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intmack_1_argbuf_rwb_r) && (! readPointer_QTree_Intmack_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intmack_1_argbuf_bufchan_buf <= readPointer_QTree_Intmack_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intwsxl_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intwsxl_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intwsxl_1_1_argbuf_r = ((! readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intwsxl_1_1_argbuf_r)
        readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d <= readPointer_QTree_Intwsxl_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d = (readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intwsxl_1_1_argbuf_rwb_r && readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intwsxl_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intwsxl_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intwsxl_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_Intwsxl_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_Intwsxl_1_1_argbuf_rwb_done = (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_Intwsxl_1_1_argbuf_rwb_r = (& readPointer_QTree_Intwsxl_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_Intwsxl_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intwsxl_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_Intwsxl_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (sc_0_11_destruct,Pointer_CTkron_kron_Int_Int_Int) > (sc_0_11_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_bufchan_d;
  logic sc_0_11_destruct_bufchan_r;
  assign sc_0_11_destruct_r = ((! sc_0_11_destruct_bufchan_d[0]) || sc_0_11_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_11_destruct_r)
        sc_0_11_destruct_bufchan_d <= sc_0_11_destruct_d;
  Pointer_CTkron_kron_Int_Int_Int_t sc_0_11_destruct_bufchan_buf;
  assign sc_0_11_destruct_bufchan_r = (! sc_0_11_destruct_bufchan_buf[0]);
  assign sc_0_11_1_argbuf_d = (sc_0_11_destruct_bufchan_buf[0] ? sc_0_11_destruct_bufchan_buf :
                               sc_0_11_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_11_1_argbuf_r && sc_0_11_destruct_bufchan_buf[0]))
        sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_11_1_argbuf_r) && (! sc_0_11_destruct_bufchan_buf[0])))
        sc_0_11_destruct_bufchan_buf <= sc_0_11_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (sc_0_15_destruct,Pointer_CTmain_mask_Int) > (sc_0_15_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t sc_0_15_destruct_bufchan_d;
  logic sc_0_15_destruct_bufchan_r;
  assign sc_0_15_destruct_r = ((! sc_0_15_destruct_bufchan_d[0]) || sc_0_15_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_15_destruct_r)
        sc_0_15_destruct_bufchan_d <= sc_0_15_destruct_d;
  Pointer_CTmain_mask_Int_t sc_0_15_destruct_bufchan_buf;
  assign sc_0_15_destruct_bufchan_r = (! sc_0_15_destruct_bufchan_buf[0]);
  assign sc_0_15_1_argbuf_d = (sc_0_15_destruct_bufchan_buf[0] ? sc_0_15_destruct_bufchan_buf :
                               sc_0_15_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_15_1_argbuf_r && sc_0_15_destruct_bufchan_buf[0]))
        sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_15_1_argbuf_r) && (! sc_0_15_destruct_bufchan_buf[0])))
        sc_0_15_destruct_bufchan_buf <= sc_0_15_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (sc_0_19_destruct,Pointer_CTmap''_map''_Int_Int_Int) > (sc_0_19_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_bufchan_d;
  logic sc_0_19_destruct_bufchan_r;
  assign sc_0_19_destruct_r = ((! sc_0_19_destruct_bufchan_d[0]) || sc_0_19_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_19_destruct_r)
        sc_0_19_destruct_bufchan_d <= sc_0_19_destruct_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  sc_0_19_destruct_bufchan_buf;
  assign sc_0_19_destruct_bufchan_r = (! sc_0_19_destruct_bufchan_buf[0]);
  assign sc_0_19_1_argbuf_d = (sc_0_19_destruct_bufchan_buf[0] ? sc_0_19_destruct_bufchan_buf :
                               sc_0_19_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_19_1_argbuf_r && sc_0_19_destruct_bufchan_buf[0]))
        sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_19_1_argbuf_r) && (! sc_0_19_destruct_bufchan_buf[0])))
        sc_0_19_destruct_bufchan_buf <= sc_0_19_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (sc_0_7_destruct,Pointer_CT$wnnz_Int) > (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_d;
  logic sc_0_7_destruct_bufchan_r;
  assign sc_0_7_destruct_r = ((! sc_0_7_destruct_bufchan_d[0]) || sc_0_7_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_7_destruct_r)
        sc_0_7_destruct_bufchan_d <= sc_0_7_destruct_d;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_buf;
  assign sc_0_7_destruct_bufchan_r = (! sc_0_7_destruct_bufchan_buf[0]);
  assign sc_0_7_1_argbuf_d = (sc_0_7_destruct_bufchan_buf[0] ? sc_0_7_destruct_bufchan_buf :
                              sc_0_7_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_7_1_argbuf_r && sc_0_7_destruct_bufchan_buf[0]))
        sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_7_1_argbuf_r) && (! sc_0_7_destruct_bufchan_buf[0])))
        sc_0_7_destruct_bufchan_buf <= sc_0_7_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (scfarg_0_1_goMux_mux,Pointer_CTkron_kron_Int_Int_Int) > (scfarg_0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CTkron_kron_Int_Int_Int_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (scfarg_0_2_goMux_mux,Pointer_CTmain_mask_Int) > (scfarg_0_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTmain_mask_Int_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (scfarg_0_3_goMux_mux,Pointer_CTmap''_map''_Int_Int_Int) > (scfarg_0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_bufchan_d;
  logic scfarg_0_3_goMux_mux_bufchan_r;
  assign scfarg_0_3_goMux_mux_r = ((! scfarg_0_3_goMux_mux_bufchan_d[0]) || scfarg_0_3_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_3_goMux_mux_r)
        scfarg_0_3_goMux_mux_bufchan_d <= scfarg_0_3_goMux_mux_d;
  \Pointer_CTmap''_map''_Int_Int_Int_t  scfarg_0_3_goMux_mux_bufchan_buf;
  assign scfarg_0_3_goMux_mux_bufchan_r = (! scfarg_0_3_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_3_1_argbuf_d = (scfarg_0_3_goMux_mux_bufchan_buf[0] ? scfarg_0_3_goMux_mux_bufchan_buf :
                                  scfarg_0_3_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_3_1_argbuf_r && scfarg_0_3_goMux_mux_bufchan_buf[0]))
        scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_3_1_argbuf_r) && (! scfarg_0_3_goMux_mux_bufchan_buf[0])))
        scfarg_0_3_goMux_mux_bufchan_buf <= scfarg_0_3_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) > (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1acr_3_destruct,Pointer_QTree_Int) > (t1acr_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1acr_3_destruct_bufchan_d;
  logic t1acr_3_destruct_bufchan_r;
  assign t1acr_3_destruct_r = ((! t1acr_3_destruct_bufchan_d[0]) || t1acr_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1acr_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1acr_3_destruct_r)
        t1acr_3_destruct_bufchan_d <= t1acr_3_destruct_d;
  Pointer_QTree_Int_t t1acr_3_destruct_bufchan_buf;
  assign t1acr_3_destruct_bufchan_r = (! t1acr_3_destruct_bufchan_buf[0]);
  assign t1acr_3_1_argbuf_d = (t1acr_3_destruct_bufchan_buf[0] ? t1acr_3_destruct_bufchan_buf :
                               t1acr_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1acr_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1acr_3_1_argbuf_r && t1acr_3_destruct_bufchan_buf[0]))
        t1acr_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1acr_3_1_argbuf_r) && (! t1acr_3_destruct_bufchan_buf[0])))
        t1acr_3_destruct_bufchan_buf <= t1acr_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2acs_2_destruct,Pointer_QTree_Int) > (t2acs_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2acs_2_destruct_bufchan_d;
  logic t2acs_2_destruct_bufchan_r;
  assign t2acs_2_destruct_r = ((! t2acs_2_destruct_bufchan_d[0]) || t2acs_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2acs_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2acs_2_destruct_r)
        t2acs_2_destruct_bufchan_d <= t2acs_2_destruct_d;
  Pointer_QTree_Int_t t2acs_2_destruct_bufchan_buf;
  assign t2acs_2_destruct_bufchan_r = (! t2acs_2_destruct_bufchan_buf[0]);
  assign t2acs_2_1_argbuf_d = (t2acs_2_destruct_bufchan_buf[0] ? t2acs_2_destruct_bufchan_buf :
                               t2acs_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2acs_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2acs_2_1_argbuf_r && t2acs_2_destruct_bufchan_buf[0]))
        t2acs_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2acs_2_1_argbuf_r) && (! t2acs_2_destruct_bufchan_buf[0])))
        t2acs_2_destruct_bufchan_buf <= t2acs_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3act_1_destruct,Pointer_QTree_Int) > (t3act_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3act_1_destruct_bufchan_d;
  logic t3act_1_destruct_bufchan_r;
  assign t3act_1_destruct_r = ((! t3act_1_destruct_bufchan_d[0]) || t3act_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3act_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3act_1_destruct_r)
        t3act_1_destruct_bufchan_d <= t3act_1_destruct_d;
  Pointer_QTree_Int_t t3act_1_destruct_bufchan_buf;
  assign t3act_1_destruct_bufchan_r = (! t3act_1_destruct_bufchan_buf[0]);
  assign t3act_1_1_argbuf_d = (t3act_1_destruct_bufchan_buf[0] ? t3act_1_destruct_bufchan_buf :
                               t3act_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3act_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3act_1_1_argbuf_r && t3act_1_destruct_bufchan_buf[0]))
        t3act_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3act_1_1_argbuf_r) && (! t3act_1_destruct_bufchan_buf[0])))
        t3act_1_destruct_bufchan_buf <= t3act_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4acu_destruct,Pointer_QTree_Int) > (t4acu_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4acu_destruct_bufchan_d;
  logic t4acu_destruct_bufchan_r;
  assign t4acu_destruct_r = ((! t4acu_destruct_bufchan_d[0]) || t4acu_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4acu_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4acu_destruct_r) t4acu_destruct_bufchan_d <= t4acu_destruct_d;
  Pointer_QTree_Int_t t4acu_destruct_bufchan_buf;
  assign t4acu_destruct_bufchan_r = (! t4acu_destruct_bufchan_buf[0]);
  assign t4acu_1_argbuf_d = (t4acu_destruct_bufchan_buf[0] ? t4acu_destruct_bufchan_buf :
                             t4acu_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4acu_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4acu_1_argbuf_r && t4acu_destruct_bufchan_buf[0]))
        t4acu_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4acu_1_argbuf_r) && (! t4acu_destruct_bufchan_buf[0])))
        t4acu_destruct_bufchan_buf <= t4acu_destruct_bufchan_d;
  
  /* buf (Ty Int) : (v'acE_2_2,Int) > (v'acE_2_2_argbuf,Int) */
  Int_t \v'acE_2_2_bufchan_d ;
  logic \v'acE_2_2_bufchan_r ;
  assign \v'acE_2_2_r  = ((! \v'acE_2_2_bufchan_d [0]) || \v'acE_2_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_2_2_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'acE_2_2_r ) \v'acE_2_2_bufchan_d  <= \v'acE_2_2_d ;
  Int_t \v'acE_2_2_bufchan_buf ;
  assign \v'acE_2_2_bufchan_r  = (! \v'acE_2_2_bufchan_buf [0]);
  assign \v'acE_2_2_argbuf_d  = (\v'acE_2_2_bufchan_buf [0] ? \v'acE_2_2_bufchan_buf  :
                                 \v'acE_2_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_2_2_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acE_2_2_argbuf_r  && \v'acE_2_2_bufchan_buf [0]))
        \v'acE_2_2_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acE_2_2_argbuf_r ) && (! \v'acE_2_2_bufchan_buf [0])))
        \v'acE_2_2_bufchan_buf  <= \v'acE_2_2_bufchan_d ;
  
  /* fork (Ty Int) : (v'acE_2_destruct,Int) > [(v'acE_2_1,Int),
                                          (v'acE_2_2,Int)] */
  logic [1:0] \v'acE_2_destruct_emitted ;
  logic [1:0] \v'acE_2_destruct_done ;
  assign \v'acE_2_1_d  = {\v'acE_2_destruct_d [32:1],
                          (\v'acE_2_destruct_d [0] && (! \v'acE_2_destruct_emitted [0]))};
  assign \v'acE_2_2_d  = {\v'acE_2_destruct_d [32:1],
                          (\v'acE_2_destruct_d [0] && (! \v'acE_2_destruct_emitted [1]))};
  assign \v'acE_2_destruct_done  = (\v'acE_2_destruct_emitted  | ({\v'acE_2_2_d [0],
                                                                   \v'acE_2_1_d [0]} & {\v'acE_2_2_r ,
                                                                                        \v'acE_2_1_r }));
  assign \v'acE_2_destruct_r  = (& \v'acE_2_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_2_destruct_emitted  <= 2'd0;
    else
      \v'acE_2_destruct_emitted  <= (\v'acE_2_destruct_r  ? 2'd0 :
                                     \v'acE_2_destruct_done );
  
  /* buf (Ty Int) : (v'acE_3_2,Int) > (v'acE_3_2_argbuf,Int) */
  Int_t \v'acE_3_2_bufchan_d ;
  logic \v'acE_3_2_bufchan_r ;
  assign \v'acE_3_2_r  = ((! \v'acE_3_2_bufchan_d [0]) || \v'acE_3_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_3_2_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'acE_3_2_r ) \v'acE_3_2_bufchan_d  <= \v'acE_3_2_d ;
  Int_t \v'acE_3_2_bufchan_buf ;
  assign \v'acE_3_2_bufchan_r  = (! \v'acE_3_2_bufchan_buf [0]);
  assign \v'acE_3_2_argbuf_d  = (\v'acE_3_2_bufchan_buf [0] ? \v'acE_3_2_bufchan_buf  :
                                 \v'acE_3_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_3_2_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acE_3_2_argbuf_r  && \v'acE_3_2_bufchan_buf [0]))
        \v'acE_3_2_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acE_3_2_argbuf_r ) && (! \v'acE_3_2_bufchan_buf [0])))
        \v'acE_3_2_bufchan_buf  <= \v'acE_3_2_bufchan_d ;
  
  /* fork (Ty Int) : (v'acE_3_destruct,Int) > [(v'acE_3_1,Int),
                                          (v'acE_3_2,Int)] */
  logic [1:0] \v'acE_3_destruct_emitted ;
  logic [1:0] \v'acE_3_destruct_done ;
  assign \v'acE_3_1_d  = {\v'acE_3_destruct_d [32:1],
                          (\v'acE_3_destruct_d [0] && (! \v'acE_3_destruct_emitted [0]))};
  assign \v'acE_3_2_d  = {\v'acE_3_destruct_d [32:1],
                          (\v'acE_3_destruct_d [0] && (! \v'acE_3_destruct_emitted [1]))};
  assign \v'acE_3_destruct_done  = (\v'acE_3_destruct_emitted  | ({\v'acE_3_2_d [0],
                                                                   \v'acE_3_1_d [0]} & {\v'acE_3_2_r ,
                                                                                        \v'acE_3_1_r }));
  assign \v'acE_3_destruct_r  = (& \v'acE_3_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_3_destruct_emitted  <= 2'd0;
    else
      \v'acE_3_destruct_emitted  <= (\v'acE_3_destruct_r  ? 2'd0 :
                                     \v'acE_3_destruct_done );
  
  /* buf (Ty Int) : (v'acE_4_destruct,Int) > (v'acE_4_1_argbuf,Int) */
  Int_t \v'acE_4_destruct_bufchan_d ;
  logic \v'acE_4_destruct_bufchan_r ;
  assign \v'acE_4_destruct_r  = ((! \v'acE_4_destruct_bufchan_d [0]) || \v'acE_4_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'acE_4_destruct_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\v'acE_4_destruct_r )
        \v'acE_4_destruct_bufchan_d  <= \v'acE_4_destruct_d ;
  Int_t \v'acE_4_destruct_bufchan_buf ;
  assign \v'acE_4_destruct_bufchan_r  = (! \v'acE_4_destruct_bufchan_buf [0]);
  assign \v'acE_4_1_argbuf_d  = (\v'acE_4_destruct_bufchan_buf [0] ? \v'acE_4_destruct_bufchan_buf  :
                                 \v'acE_4_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \v'acE_4_destruct_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'acE_4_1_argbuf_r  && \v'acE_4_destruct_bufchan_buf [0]))
        \v'acE_4_destruct_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'acE_4_1_argbuf_r ) && (! \v'acE_4_destruct_bufchan_buf [0])))
        \v'acE_4_destruct_bufchan_buf  <= \v'acE_4_destruct_bufchan_d ;
  
  /* buf (Ty Int) : (vacG_destruct,Int) > (vacG_1_argbuf,Int) */
  Int_t vacG_destruct_bufchan_d;
  logic vacG_destruct_bufchan_r;
  assign vacG_destruct_r = ((! vacG_destruct_bufchan_d[0]) || vacG_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacG_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vacG_destruct_r) vacG_destruct_bufchan_d <= vacG_destruct_d;
  Int_t vacG_destruct_bufchan_buf;
  assign vacG_destruct_bufchan_r = (! vacG_destruct_bufchan_buf[0]);
  assign vacG_1_argbuf_d = (vacG_destruct_bufchan_buf[0] ? vacG_destruct_bufchan_buf :
                            vacG_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacG_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vacG_1_argbuf_r && vacG_destruct_bufchan_buf[0]))
        vacG_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vacG_1_argbuf_r) && (! vacG_destruct_bufchan_buf[0])))
        vacG_destruct_bufchan_buf <= vacG_destruct_bufchan_d;
  
  /* buf (Ty Int) : (vacP_destruct,Int) > (vacP_1_argbuf,Int) */
  Int_t vacP_destruct_bufchan_d;
  logic vacP_destruct_bufchan_r;
  assign vacP_destruct_r = ((! vacP_destruct_bufchan_d[0]) || vacP_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacP_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vacP_destruct_r) vacP_destruct_bufchan_d <= vacP_destruct_d;
  Int_t vacP_destruct_bufchan_buf;
  assign vacP_destruct_bufchan_r = (! vacP_destruct_bufchan_buf[0]);
  assign vacP_1_argbuf_d = (vacP_destruct_bufchan_buf[0] ? vacP_destruct_bufchan_buf :
                            vacP_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacP_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vacP_1_argbuf_r && vacP_destruct_bufchan_buf[0]))
        vacP_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vacP_1_argbuf_r) && (! vacP_destruct_bufchan_buf[0])))
        vacP_destruct_bufchan_buf <= vacP_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (lizzieLet16_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet27_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet27_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet27_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca2_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet29_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet29_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet29_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca3_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (lizzieLet13_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf :
                                     writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca2_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca1_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf :
                                                                   writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca0_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                         1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) > (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d <= {16'd0,
                                                                    1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_r)
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d = (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf :
                                                                  writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0,
                                                                      1'd0};
    else
      if ((writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r && writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0,
                                                                        1'd0};
      else if (((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Int_Int_Int) : (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb,Pointer_CTkron_kron_Int_Int_Int) > (sca3_1_1_argbuf,Pointer_CTkron_kron_Int_Int_Int) */
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r = ((! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_r)
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Int_Int_Int_t writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf :
                              writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Int_Int_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet15_1_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet15_1_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf :
                                                             writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet15_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca3_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet15_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet24_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet24_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet24_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet24_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf :
                                    writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet24_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet36_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet36_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet36_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca2_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet37_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet37_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet37_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet37_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca1_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet37_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet38_1_argbuf,Pointer_CTmain_mask_Int) > (writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_r = ((! writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet38_1_argbuf_r)
        writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d <= writeCTmain_mask_IntlizzieLet38_1_argbuf_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_r = (! writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_d = (writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf :
                                                           writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_r && writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_r) && (! writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_buf <= writeCTmain_mask_IntlizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Int) : (writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb,Pointer_CTmain_mask_Int) > (sca0_2_1_argbuf,Pointer_CTmain_mask_Int) */
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_r = ((! writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                 1'd0};
    else
      if (writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_r)
        writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Int_t writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                     1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca3_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca3_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca3_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet21_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (lizzieLet9_1_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet9_1_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca2_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca2_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca2_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet41_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca1_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca1_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca1_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet42_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) > (writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_d  = (\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf  :
                                                                       \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_r  && \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Int_Int_Int) : (writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb,Pointer_CTmap''_map''_Int_Int_Int) > (sca0_3_1_argbuf,Pointer_CTmap''_map''_Int_Int_Int) */
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_r )
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Int_Int_Int_t  \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_3_1_argbuf_d = (\writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca0_3_1_argbuf_r && \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca0_3_1_argbuf_r) && (! \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Int_Int_IntlizzieLet43_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_r = ((! writeQTree_IntlizzieLet13_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_r)
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_d = (writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet13_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet13_1_argbuf_rwb_r && writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet13_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_2_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet14_2_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet14_2_1_argbuf_r = ((! writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_2_1_argbuf_r)
        writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet14_2_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet14_2_1_argbuf_rwb_d = (writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet14_2_1_argbuf_rwb_r && writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet14_2_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet14_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_2_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet14_2_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet14_2_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet14_2_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet14_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet16_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_1_argbuf_r = ((! writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_1_argbuf_r)
        writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet16_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet16_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet16_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet16_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet16_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet16_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet16_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_r = ((! writeQTree_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_r)
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_d = (writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet18_1_argbuf_rwb_r && writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet18_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet19_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet19_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet19_1_argbuf_r = ((! writeQTree_IntlizzieLet19_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet19_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet19_1_argbuf_r)
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet19_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet19_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_d = (writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet19_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet19_1_argbuf_rwb_r && writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet19_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet19_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet19_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet19_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet19_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet19_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet19_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_r = ((! writeQTree_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_r)
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_d = (writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet20_1_argbuf_rwb_r && writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet20_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_r = ((! writeQTree_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_r)
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_d = (writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet22_1_argbuf_rwb_r && writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet22_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_r = ((! writeQTree_IntlizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_r)
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_d = (writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet34_1_argbuf_rwb_r && writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet34_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet39_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_argbuf_r = ((! writeQTree_IntlizzieLet39_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_argbuf_r)
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet39_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_d = (writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet39_1_argbuf_rwb_r && writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet39_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet39_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet39_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet44_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet44_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet44_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet44_1_argbuf_r = ((! writeQTree_IntlizzieLet44_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet44_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet44_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet44_1_argbuf_r)
        writeQTree_IntlizzieLet44_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet44_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet44_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet44_1_argbuf_rwb_d = (writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet44_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet44_1_argbuf_rwb_r && writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet44_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet44_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet44_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet44_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet44_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet44_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet44_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_3_1_argbuf_d = (writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_3_1_argbuf_r && writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_3_1_argbuf_r) && (! writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet44_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet12_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsxl_1_goMux_mux,Pointer_QTree_Int) > (wsxl_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsxl_1_goMux_mux_bufchan_d;
  logic wsxl_1_goMux_mux_bufchan_r;
  assign wsxl_1_goMux_mux_r = ((! wsxl_1_goMux_mux_bufchan_d[0]) || wsxl_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsxl_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsxl_1_goMux_mux_r)
        wsxl_1_goMux_mux_bufchan_d <= wsxl_1_goMux_mux_d;
  Pointer_QTree_Int_t wsxl_1_goMux_mux_bufchan_buf;
  assign wsxl_1_goMux_mux_bufchan_r = (! wsxl_1_goMux_mux_bufchan_buf[0]);
  assign wsxl_1_1_argbuf_d = (wsxl_1_goMux_mux_bufchan_buf[0] ? wsxl_1_goMux_mux_bufchan_buf :
                              wsxl_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsxl_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsxl_1_1_argbuf_r && wsxl_1_goMux_mux_bufchan_buf[0]))
        wsxl_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsxl_1_1_argbuf_r) && (! wsxl_1_goMux_mux_bufchan_buf[0])))
        wsxl_1_goMux_mux_bufchan_buf <= wsxl_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) > (lizzieLet28_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d;
  logic wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_r;
  assign wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_r = ((! wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d[0]) || wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_r)
        wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d <= wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_d;
  CT$wnnz_Int_t wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf;
  assign wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_r = (! wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf[0] ? wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf :
                                   wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf[0]))
        wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf[0])))
        wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_buf <= wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int1) : [(wwsxo_2_destruct,Int#),
                                (lizzieLet26_4Lcall_$wnnz_Int2,Int#),
                                (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                (q4acY_2_destruct,Pointer_QTree_Int)] > (wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) */
  assign wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_d = Lcall_$wnnz_Int1_dc((& {wwsxo_2_destruct_d[0],
                                                                                                               lizzieLet26_4Lcall_$wnnz_Int2_d[0],
                                                                                                               sc_0_5_destruct_d[0],
                                                                                                               q4acY_2_destruct_d[0]}), wwsxo_2_destruct_d, lizzieLet26_4Lcall_$wnnz_Int2_d, sc_0_5_destruct_d, q4acY_2_destruct_d);
  assign {wwsxo_2_destruct_r,
          lizzieLet26_4Lcall_$wnnz_Int2_r,
          sc_0_5_destruct_r,
          q4acY_2_destruct_r} = {4 {(wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_r && wwsxo_2_1lizzieLet26_4Lcall_$wnnz_Int2_1sc_0_5_1q4acY_2_1Lcall_$wnnz_Int1_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) > (lizzieLet29_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  logic wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r;
  assign wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r = ((! wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d[0]) || wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= {115'd0,
                                                                                               1'd0};
    else
      if (wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r)
        wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  CT$wnnz_Int_t wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf;
  assign wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r = (! wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0] ? wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf :
                                   wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]))
        wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0])))
        wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int0) : [(wwsxo_3_destruct,Int#),
                                (ww1XyC_1_destruct,Int#),
                                (lizzieLet26_4Lcall_$wnnz_Int1,Int#),
                                (sc_0_6_destruct,Pointer_CT$wnnz_Int)] > (wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) */
  assign wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d = Lcall_$wnnz_Int0_dc((& {wwsxo_3_destruct_d[0],
                                                                                                                ww1XyC_1_destruct_d[0],
                                                                                                                lizzieLet26_4Lcall_$wnnz_Int1_d[0],
                                                                                                                sc_0_6_destruct_d[0]}), wwsxo_3_destruct_d, ww1XyC_1_destruct_d, lizzieLet26_4Lcall_$wnnz_Int1_d, sc_0_6_destruct_d);
  assign {wwsxo_3_destruct_r,
          ww1XyC_1_destruct_r,
          lizzieLet26_4Lcall_$wnnz_Int1_r,
          sc_0_6_destruct_r} = {4 {(wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r && wwsxo_3_1ww1XyC_1_1lizzieLet26_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsxo_4_1ww1XyC_2_1_Add32,Int#) (ww2XyF_1_destruct,Int#) > (es_6_1ww2XyF_1_1_Add32,Int#) */
  assign es_6_1ww2XyF_1_1_Add32_d = {(wwsxo_4_1ww1XyC_2_1_Add32_d[32:1] + ww2XyF_1_destruct_d[32:1]),
                                     (wwsxo_4_1ww1XyC_2_1_Add32_d[0] && ww2XyF_1_destruct_d[0])};
  assign {wwsxo_4_1ww1XyC_2_1_Add32_r,
          ww2XyF_1_destruct_r} = {2 {(es_6_1ww2XyF_1_1_Add32_r && es_6_1ww2XyF_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsxo_4_destruct,Int#) (ww1XyC_2_destruct,Int#) > (wwsxo_4_1ww1XyC_2_1_Add32,Int#) */
  assign wwsxo_4_1ww1XyC_2_1_Add32_d = {(wwsxo_4_destruct_d[32:1] + ww1XyC_2_destruct_d[32:1]),
                                        (wwsxo_4_destruct_d[0] && ww1XyC_2_destruct_d[0])};
  assign {wwsxo_4_destruct_r,
          ww1XyC_2_destruct_r} = {2 {(wwsxo_4_1ww1XyC_2_1_Add32_r && wwsxo_4_1ww1XyC_2_1_Add32_d[0])}};
  
  /* buf (Ty Int) : (xac0_1,Int) > (xac0_1_argbuf,Int) */
  Int_t xac0_1_bufchan_d;
  logic xac0_1_bufchan_r;
  assign xac0_1_r = ((! xac0_1_bufchan_d[0]) || xac0_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xac0_1_bufchan_d <= {32'd0, 1'd0};
    else if (xac0_1_r) xac0_1_bufchan_d <= xac0_1_d;
  Int_t xac0_1_bufchan_buf;
  assign xac0_1_bufchan_r = (! xac0_1_bufchan_buf[0]);
  assign xac0_1_argbuf_d = (xac0_1_bufchan_buf[0] ? xac0_1_bufchan_buf :
                            xac0_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xac0_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((xac0_1_argbuf_r && xac0_1_bufchan_buf[0]))
        xac0_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! xac0_1_argbuf_r) && (! xac0_1_bufchan_buf[0])))
        xac0_1_bufchan_buf <= xac0_1_bufchan_d;
endmodule