`timescale 1ns/1ns
import mMapAdd_package::*;

module mMapAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t m1aex_0_d,
  output logic m1aex_0_r,
  input Pointer_QTree_Int_t m2aey_1_d,
  output logic m2aey_1_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_1_1I#_dout ,
  input logic \es_1_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (m1aex_0, 16, 65536, Pointer_QTree_Int), (m2aey_1, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_1_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
CTf__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[16p,16p,16p,16p]) (3,[16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTf_f 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
TupGo___Pointer_QTree_Bool 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Bool___Pointer_CT__024wnnz 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_CTf__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,16p,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go__3_d;
  logic go__3_r;
  Go_t go__4_d;
  logic go__4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  \Word16#_t  initHP_CT$wnnz_d;
  logic initHP_CT$wnnz_r;
  \Word16#_t  incrHP_CT$wnnz_d;
  logic incrHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_d;
  logic incrHP_mergeCT$wnnz_r;
  Go_t incrHP_CT$wnnz1_d;
  logic incrHP_CT$wnnz1_r;
  Go_t incrHP_CT$wnnz2_d;
  logic incrHP_CT$wnnz2_r;
  \Word16#_t  addHP_CT$wnnz_d;
  logic addHP_CT$wnnz_r;
  \Word16#_t  mergeHP_CT$wnnz_d;
  logic mergeHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_buf_d;
  logic incrHP_mergeCT$wnnz_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_buf_d;
  logic mergeHP_CT$wnnz_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_d;
  logic forkHP1_CT$wnnz_r;
  \Word16#_t  forkHP1_CT$wnn2_d;
  logic forkHP1_CT$wnn2_r;
  \Word16#_t  forkHP1_CT$wnn3_d;
  logic forkHP1_CT$wnn3_r;
  C2_t memMergeChoice_CT$wnnz_d;
  logic memMergeChoice_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_d;
  logic memMergeIn_CT$wnnz_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_d;
  logic memOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memReadOut_CT$wnnz_d;
  logic memReadOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memWriteOut_CT$wnnz_d;
  logic memWriteOut_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_dbuf_d;
  logic memMergeIn_CT$wnnz_dbuf_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_rbuf_d;
  logic memMergeIn_CT$wnnz_rbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_dbuf_d;
  logic memOut_CT$wnnz_dbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_rbuf_d;
  logic memOut_CT$wnnz_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_d;
  logic destructReadIn_CT$wnnz_r;
  MemIn_CT$wnnz_t dconReadIn_CT$wnnz_d;
  logic dconReadIn_CT$wnnz_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_d;
  logic writeMerge_choice_CT$wnnz_r;
  CT$wnnz_t writeMerge_data_CT$wnnz_d;
  logic writeMerge_data_CT$wnnz_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_d;
  logic writeCT$wnnzlizzieLet2_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_d;
  logic writeCT$wnnzlizzieLet45_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_d;
  logic writeCT$wnnzlizzieLet46_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_d;
  logic writeCT$wnnzlizzieLet47_1_argbuf_r;
  MemIn_CT$wnnz_t dconWriteIn_CT$wnnz_d;
  logic dconWriteIn_CT$wnnz_r;
  Pointer_CT$wnnz_t dconPtr_CT$wnnz_d;
  logic dconPtr_CT$wnnz_r;
  Pointer_CT$wnnz_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Pointer_CT$wnnz_t demuxWriteResult_CT$wnnz_d;
  logic demuxWriteResult_CT$wnnz_r;
  \Word16#_t  \initHP_CTf''''''''_f''''''''_d ;
  logic \initHP_CTf''''''''_f''''''''_r ;
  \Word16#_t  \incrHP_CTf''''''''_f''''''''_d ;
  logic \incrHP_CTf''''''''_f''''''''_r ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_r ;
  Go_t \incrHP_CTf''''''''_f''''''''1_d ;
  logic \incrHP_CTf''''''''_f''''''''1_r ;
  Go_t \incrHP_CTf''''''''_f''''''''2_d ;
  logic \incrHP_CTf''''''''_f''''''''2_r ;
  \Word16#_t  \addHP_CTf''''''''_f''''''''_d ;
  logic \addHP_CTf''''''''_f''''''''_r ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_d ;
  logic \mergeHP_CTf''''''''_f''''''''_r ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_buf_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_buf_r ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_buf_d ;
  logic \mergeHP_CTf''''''''_f''''''''_buf_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f''''''''_d ;
  logic \forkHP1_CTf''''''''_f''''''''_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f'''''''2_d ;
  logic \forkHP1_CTf''''''''_f'''''''2_r ;
  \Word16#_t  \forkHP1_CTf''''''''_f'''''''3_d ;
  logic \forkHP1_CTf''''''''_f'''''''3_r ;
  C2_t \memMergeChoice_CTf''''''''_f''''''''_d ;
  logic \memMergeChoice_CTf''''''''_f''''''''_r ;
  \MemIn_CTf''''''''_f''''''''_t  \memMergeIn_CTf''''''''_f''''''''_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_r ;
  \MemOut_CTf''''''''_f''''''''_t  \memOut_CTf''''''''_f''''''''_d ;
  logic \memOut_CTf''''''''_f''''''''_r ;
  \MemOut_CTf''''''''_f''''''''_t  \memReadOut_CTf''''''''_f''''''''_d ;
  logic \memReadOut_CTf''''''''_f''''''''_r ;
  \MemOut_CTf''''''''_f''''''''_t  \memWriteOut_CTf''''''''_f''''''''_d ;
  logic \memWriteOut_CTf''''''''_f''''''''_r ;
  \MemIn_CTf''''''''_f''''''''_t  \memMergeIn_CTf''''''''_f''''''''_dbuf_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_dbuf_r ;
  \MemIn_CTf''''''''_f''''''''_t  \memMergeIn_CTf''''''''_f''''''''_rbuf_d ;
  logic \memMergeIn_CTf''''''''_f''''''''_rbuf_r ;
  \MemOut_CTf''''''''_f''''''''_t  \memOut_CTf''''''''_f''''''''_dbuf_d ;
  logic \memOut_CTf''''''''_f''''''''_dbuf_r ;
  \MemOut_CTf''''''''_f''''''''_t  \memOut_CTf''''''''_f''''''''_rbuf_d ;
  logic \memOut_CTf''''''''_f''''''''_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf''''''''_f''''''''_d ;
  logic \destructReadIn_CTf''''''''_f''''''''_r ;
  \MemIn_CTf''''''''_f''''''''_t  \dconReadIn_CTf''''''''_f''''''''_d ;
  logic \dconReadIn_CTf''''''''_f''''''''_r ;
  \CTf''''''''_f''''''''_t  \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf''''''''_f''''''''_d ;
  logic \writeMerge_choice_CTf''''''''_f''''''''_r ;
  \CTf''''''''_f''''''''_t  \writeMerge_data_CTf''''''''_f''''''''_d ;
  logic \writeMerge_data_CTf''''''''_f''''''''_r ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_r ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_r ;
  \MemIn_CTf''''''''_f''''''''_t  \dconWriteIn_CTf''''''''_f''''''''_d ;
  logic \dconWriteIn_CTf''''''''_f''''''''_r ;
  \Pointer_CTf''''''''_f''''''''_t  \dconPtr_CTf''''''''_f''''''''_d ;
  logic \dconPtr_CTf''''''''_f''''''''_r ;
  \Pointer_CTf''''''''_f''''''''_t  _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  \Pointer_CTf''''''''_f''''''''_t  \demuxWriteResult_CTf''''''''_f''''''''_d ;
  logic \demuxWriteResult_CTf''''''''_f''''''''_r ;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Boo2_d;
  logic forkHP1_QTree_Boo2_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_BoolwspF_1_1_argbuf_d;
  logic readPointer_QTree_BoolwspF_1_1_argbuf_r;
  C18_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet19_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet20_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_d;
  logic writeQTree_BoollizzieLet21_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_d;
  logic writeQTree_BoollizzieLet27_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_d;
  logic writeQTree_BoollizzieLet32_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet41_1_argbuf_d;
  logic writeQTree_BoollizzieLet41_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  initHP_CTf_f_d;
  logic initHP_CTf_f_r;
  \Word16#_t  incrHP_CTf_f_d;
  logic incrHP_CTf_f_r;
  Go_t incrHP_mergeCTf_f_d;
  logic incrHP_mergeCTf_f_r;
  Go_t incrHP_CTf_f1_d;
  logic incrHP_CTf_f1_r;
  Go_t incrHP_CTf_f2_d;
  logic incrHP_CTf_f2_r;
  \Word16#_t  addHP_CTf_f_d;
  logic addHP_CTf_f_r;
  \Word16#_t  mergeHP_CTf_f_d;
  logic mergeHP_CTf_f_r;
  Go_t incrHP_mergeCTf_f_buf_d;
  logic incrHP_mergeCTf_f_buf_r;
  \Word16#_t  mergeHP_CTf_f_buf_d;
  logic mergeHP_CTf_f_buf_r;
  \Word16#_t  forkHP1_CTf_f_d;
  logic forkHP1_CTf_f_r;
  \Word16#_t  forkHP1_CTf_2_d;
  logic forkHP1_CTf_2_r;
  \Word16#_t  forkHP1_CTf_3_d;
  logic forkHP1_CTf_3_r;
  C2_t memMergeChoice_CTf_f_d;
  logic memMergeChoice_CTf_f_r;
  MemIn_CTf_f_t memMergeIn_CTf_f_d;
  logic memMergeIn_CTf_f_r;
  MemOut_CTf_f_t memOut_CTf_f_d;
  logic memOut_CTf_f_r;
  MemOut_CTf_f_t memReadOut_CTf_f_d;
  logic memReadOut_CTf_f_r;
  MemOut_CTf_f_t memWriteOut_CTf_f_d;
  logic memWriteOut_CTf_f_r;
  MemIn_CTf_f_t memMergeIn_CTf_f_dbuf_d;
  logic memMergeIn_CTf_f_dbuf_r;
  MemIn_CTf_f_t memMergeIn_CTf_f_rbuf_d;
  logic memMergeIn_CTf_f_rbuf_r;
  MemOut_CTf_f_t memOut_CTf_f_dbuf_d;
  logic memOut_CTf_f_dbuf_r;
  MemOut_CTf_f_t memOut_CTf_f_rbuf_d;
  logic memOut_CTf_f_rbuf_r;
  \Word16#_t  destructReadIn_CTf_f_d;
  logic destructReadIn_CTf_f_r;
  MemIn_CTf_f_t dconReadIn_CTf_f_d;
  logic dconReadIn_CTf_f_r;
  CTf_f_t readPointer_CTf_fscfarg_0_2_1_argbuf_d;
  logic readPointer_CTf_fscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTf_f_d;
  logic writeMerge_choice_CTf_f_r;
  CTf_f_t writeMerge_data_CTf_f_d;
  logic writeMerge_data_CTf_f_r;
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_d;
  logic writeCTf_flizzieLet38_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_d;
  logic writeCTf_flizzieLet43_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_d;
  logic writeCTf_flizzieLet54_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_d;
  logic writeCTf_flizzieLet55_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_d;
  logic writeCTf_flizzieLet56_1_argbuf_r;
  MemIn_CTf_f_t dconWriteIn_CTf_f_d;
  logic dconWriteIn_CTf_f_r;
  Pointer_CTf_f_t dconPtr_CTf_f_d;
  logic dconPtr_CTf_f_r;
  Pointer_CTf_f_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_CTf_f_t demuxWriteResult_CTf_f_d;
  logic demuxWriteResult_CTf_f_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C3_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1ae6_1_argbuf_d;
  logic readPointer_QTree_Intm1ae6_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm2ae7_1_argbuf_d;
  logic readPointer_QTree_Intm2ae7_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  Go_t \$wnnzTupGo___Pointer_QTree_Boolgo_12_d ;
  logic \$wnnzTupGo___Pointer_QTree_Boolgo_12_r ;
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwspF_d ;
  logic \$wnnzTupGo___Pointer_QTree_BoolwspF_r ;
  Go_t go_12_1_d;
  logic go_12_1_r;
  Go_t go_12_2_d;
  logic go_12_2_r;
  Pointer_QTree_Bool_t wspF_1_argbuf_d;
  logic wspF_1_argbuf_r;
  Int_t \es_1_1I#_d ;
  logic \es_1_1I#_r ;
  Pointer_QTree_Int_t blae4_1_1_argbuf_d;
  logic blae4_1_1_argbuf_r;
  Pointer_QTree_Int_t blaec_1_argbuf_d;
  logic blaec_1_argbuf_r;
  Go_t boolConvert_1TupGo___Boolgo_4_d;
  logic boolConvert_1TupGo___Boolgo_4_r;
  Bool_t boolConvert_1TupGo___Boolbool_3_d;
  logic boolConvert_1TupGo___Boolbool_3_r;
  Bool_t bool_3_1_d;
  logic bool_3_1_r;
  Bool_t bool_3_2_d;
  logic bool_3_2_r;
  MyBool_t lizzieLet7_1_d;
  logic lizzieLet7_1_r;
  MyBool_t lizzieLet7_2_d;
  logic lizzieLet7_2_r;
  Go_t boolConvert_2TupGo___Boolgo_3_d;
  logic boolConvert_2TupGo___Boolgo_3_r;
  Bool_t boolConvert_2TupGo___Boolbool_2_d;
  logic boolConvert_2TupGo___Boolbool_2_r;
  Bool_t bool_2_1_d;
  logic bool_2_1_r;
  Bool_t bool_2_2_d;
  logic bool_2_2_r;
  MyBool_t lizzieLet17_1_d;
  logic lizzieLet17_1_r;
  MyBool_t lizzieLet17_2_d;
  logic lizzieLet17_2_r;
  Go_t boolConvert_3TupGo___Boolgo_2_d;
  logic boolConvert_3TupGo___Boolgo_2_r;
  Bool_t boolConvert_3TupGo___Boolbool_1_d;
  logic boolConvert_3TupGo___Boolbool_1_r;
  Bool_t bool_1_1_d;
  logic bool_1_1_r;
  Bool_t bool_1_2_d;
  logic bool_1_2_r;
  MyBool_t lizzieLet25_1_d;
  logic lizzieLet25_1_r;
  MyBool_t lizzieLet25_2_d;
  logic lizzieLet25_2_r;
  Go_t boolConvert_4TupGo___Boolgo_1_d;
  logic boolConvert_4TupGo___Boolgo_1_r;
  Bool_t boolConvert_4TupGo___Boolbool_d;
  logic boolConvert_4TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet30_1_d;
  logic lizzieLet30_1_r;
  MyBool_t lizzieLet30_2_d;
  logic lizzieLet30_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_4_resbuf_d;
  logic boolConvert_4_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  Go_t bool_1_1False_d;
  logic bool_1_1False_r;
  Go_t bool_1_1True_d;
  logic bool_1_1True_r;
  MyBool_t bool_1_1False_1MyFalse_d;
  logic bool_1_1False_1MyFalse_r;
  MyBool_t boolConvert_3_resbuf_d;
  logic boolConvert_3_resbuf_r;
  MyBool_t bool_1_1True_1MyTrue_d;
  logic bool_1_1True_1MyTrue_r;
  MyBool_t bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_d;
  logic bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t bool_2_1False_d;
  logic bool_2_1False_r;
  Go_t bool_2_1True_d;
  logic bool_2_1True_r;
  MyBool_t bool_2_1False_1MyFalse_d;
  logic bool_2_1False_1MyFalse_r;
  MyBool_t boolConvert_2_resbuf_d;
  logic boolConvert_2_resbuf_r;
  MyBool_t bool_2_1True_1MyTrue_d;
  logic bool_2_1True_1MyTrue_r;
  MyBool_t bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_d;
  logic bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_r;
  Go_t bool_3_1False_d;
  logic bool_3_1False_r;
  Go_t bool_3_1True_d;
  logic bool_3_1True_r;
  MyBool_t bool_3_1False_1MyFalse_d;
  logic bool_3_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_3_1True_1MyTrue_d;
  logic bool_3_1True_1MyTrue_r;
  MyBool_t bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_d;
  logic bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_r;
  Pointer_QTree_Int_t brae5_1_argbuf_d;
  logic brae5_1_argbuf_r;
  Pointer_QTree_Int_t braed_1_argbuf_d;
  logic braed_1_argbuf_r;
  Go_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_r;
  Pointer_QTree_Bool_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_r;
  Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_r;
  Go_t call_$wnnz_initBufi_d;
  logic call_$wnnz_initBufi_r;
  C5_t go_13_goMux_choice_d;
  logic go_13_goMux_choice_r;
  Go_t go_13_goMux_data_d;
  logic go_13_goMux_data_r;
  Go_t call_$wnnz_unlockFork1_d;
  logic call_$wnnz_unlockFork1_r;
  Go_t call_$wnnz_unlockFork2_d;
  logic call_$wnnz_unlockFork2_r;
  Go_t call_$wnnz_unlockFork3_d;
  logic call_$wnnz_unlockFork3_r;
  Go_t call_$wnnz_initBuf_d;
  logic call_$wnnz_initBuf_r;
  Go_t call_$wnnz_goMux1_d;
  logic call_$wnnz_goMux1_r;
  Pointer_QTree_Bool_t call_$wnnz_goMux2_d;
  logic call_$wnnz_goMux2_r;
  Pointer_CT$wnnz_t call_$wnnz_goMux3_d;
  logic call_$wnnz_goMux3_r;
  Go_t \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d ;
  logic \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_r ;
  Pointer_QTree_Int_t \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d ;
  logic \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_r ;
  \Pointer_CTf''''''''_f''''''''_t  \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d ;
  logic \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_r ;
  Go_t \call_f''''''''_f''''''''_initBufi_d ;
  logic \call_f''''''''_f''''''''_initBufi_r ;
  C5_t go_14_goMux_choice_d;
  logic go_14_goMux_choice_r;
  Go_t go_14_goMux_data_d;
  logic go_14_goMux_data_r;
  Go_t \call_f''''''''_f''''''''_unlockFork1_d ;
  logic \call_f''''''''_f''''''''_unlockFork1_r ;
  Go_t \call_f''''''''_f''''''''_unlockFork2_d ;
  logic \call_f''''''''_f''''''''_unlockFork2_r ;
  Go_t \call_f''''''''_f''''''''_unlockFork3_d ;
  logic \call_f''''''''_f''''''''_unlockFork3_r ;
  Go_t \call_f''''''''_f''''''''_initBuf_d ;
  logic \call_f''''''''_f''''''''_initBuf_r ;
  Go_t \call_f''''''''_f''''''''_goMux1_d ;
  logic \call_f''''''''_f''''''''_goMux1_r ;
  Pointer_QTree_Int_t \call_f''''''''_f''''''''_goMux2_d ;
  logic \call_f''''''''_f''''''''_goMux2_r ;
  \Pointer_CTf''''''''_f''''''''_t  \call_f''''''''_f''''''''_goMux3_d ;
  logic \call_f''''''''_f''''''''_goMux3_r ;
  Go_t call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d;
  logic call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_r;
  Pointer_QTree_Int_t call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d;
  logic call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_r;
  Pointer_QTree_Int_t call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d;
  logic call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_r;
  Pointer_CTf_f_t call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d;
  logic call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_r;
  Go_t call_f_f_initBufi_d;
  logic call_f_f_initBufi_r;
  C5_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t call_f_f_unlockFork1_d;
  logic call_f_f_unlockFork1_r;
  Go_t call_f_f_unlockFork2_d;
  logic call_f_f_unlockFork2_r;
  Go_t call_f_f_unlockFork3_d;
  logic call_f_f_unlockFork3_r;
  Go_t call_f_f_unlockFork4_d;
  logic call_f_f_unlockFork4_r;
  Go_t call_f_f_initBuf_d;
  logic call_f_f_initBuf_r;
  Go_t call_f_f_goMux1_d;
  logic call_f_f_goMux1_r;
  Pointer_QTree_Int_t call_f_f_goMux2_d;
  logic call_f_f_goMux2_r;
  Pointer_QTree_Int_t call_f_f_goMux3_d;
  logic call_f_f_goMux3_r;
  Pointer_CTf_f_t call_f_f_goMux4_d;
  logic call_f_f_goMux4_r;
  QTree_Bool_t lizzieLet20_1_1_argbuf_d;
  logic lizzieLet20_1_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  QTree_Bool_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  \Int#_t  es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_d;
  logic es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_r;
  C4_t \f''''''''1_choice_d ;
  logic \f''''''''1_choice_r ;
  TupGo_t \f''''''''1_data_d ;
  logic \f''''''''1_data_r ;
  MyBool_t go_16_1MyTrue_d;
  logic go_16_1MyTrue_r;
  Pointer_QTree_Bool_t \f''''''''1_resbuf_d ;
  logic \f''''''''1_resbuf_r ;
  Pointer_QTree_Bool_t \f''''''''1_2_argbuf_d ;
  logic \f''''''''1_2_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Bool_t \f''''''''1_3_argbuf_d ;
  logic \f''''''''1_3_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  Pointer_QTree_Bool_t \f''''''''1_4_argbuf_d ;
  logic \f''''''''1_4_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Pointer_QTree_Bool_t \f''''''''1_1_d ;
  logic \f''''''''1_1_r ;
  Pointer_QTree_Bool_t \f''''''''1_2_d ;
  logic \f''''''''1_2_r ;
  Pointer_QTree_Bool_t \f''''''''1_3_d ;
  logic \f''''''''1_3_r ;
  Pointer_QTree_Bool_t \f''''''''1_4_d ;
  logic \f''''''''1_4_r ;
  Go_t \f''''''''1TupGogo_16_d ;
  logic \f''''''''1TupGogo_16_r ;
  Pointer_QTree_Bool_t lizzieLet18_2_1_argbuf_d;
  logic lizzieLet18_2_1_argbuf_r;
  C8_t \f''''''''_f''''''''_choice_d ;
  logic \f''''''''_f''''''''_choice_r ;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''_data_d ;
  logic \f''''''''_f''''''''_data_r ;
  Go_t go_17_1_d;
  logic go_17_1_r;
  Go_t go_17_2_d;
  logic go_17_2_r;
  Pointer_QTree_Int_t q4a8u_1_1_argbuf_d;
  logic q4a8u_1_1_argbuf_r;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_resbuf_d ;
  logic \f''''''''_f''''''''_resbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_2_argbuf_d ;
  logic \f''''''''_f''''''''_2_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_3_argbuf_d ;
  logic \f''''''''_f''''''''_3_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_4_argbuf_d ;
  logic \f''''''''_f''''''''_4_argbuf_r ;
  QTree_Bool_t es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_d;
  logic es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_5_argbuf_d ;
  logic \f''''''''_f''''''''_5_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_6_argbuf_d ;
  logic \f''''''''_f''''''''_6_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_7_argbuf_d ;
  logic \f''''''''_f''''''''_7_argbuf_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_8_argbuf_d ;
  logic \f''''''''_f''''''''_8_argbuf_r ;
  QTree_Bool_t es_5_1es_6_1es_7_1es_8_1QNode_Bool_d;
  logic es_5_1es_6_1es_7_1es_8_1QNode_Bool_r;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_1_d ;
  logic \f''''''''_f''''''''_1_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_2_d ;
  logic \f''''''''_f''''''''_2_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_3_d ;
  logic \f''''''''_f''''''''_3_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_4_d ;
  logic \f''''''''_f''''''''_4_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_5_d ;
  logic \f''''''''_f''''''''_5_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_6_d ;
  logic \f''''''''_f''''''''_6_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_7_d ;
  logic \f''''''''_f''''''''_7_r ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_8_d ;
  logic \f''''''''_f''''''''_8_r ;
  Go_t \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_r ;
  Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_r ;
  Go_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_r;
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_r;
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_r;
  Go_t go_18_1_d;
  logic go_18_1_r;
  Go_t go_18_2_d;
  logic go_18_2_r;
  Pointer_QTree_Int_t m1ae6_1_1_argbuf_d;
  logic m1ae6_1_1_argbuf_r;
  Pointer_QTree_Int_t m2ae7_1_1_argbuf_d;
  logic m2ae7_1_1_argbuf_r;
  Pointer_QTree_Bool_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  Go_t go_1_argbuf_d;
  logic go_1_argbuf_r;
  CT$wnnz_t go_12_1L$wnnzsbos_d;
  logic go_12_1L$wnnzsbos_r;
  CT$wnnz_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_12_2_argbuf_d;
  logic go_12_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r;
  C5_t go_13_goMux_choice_1_d;
  logic go_13_goMux_choice_1_r;
  C5_t go_13_goMux_choice_2_d;
  logic go_13_goMux_choice_2_r;
  Pointer_QTree_Bool_t wspF_1_goMux_mux_d;
  logic wspF_1_goMux_mux_r;
  Pointer_CT$wnnz_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_14_goMux_choice_1_d;
  logic go_14_goMux_choice_1_r;
  C5_t go_14_goMux_choice_2_d;
  logic go_14_goMux_choice_2_r;
  Pointer_QTree_Int_t q4a8u_goMux_mux_d;
  logic q4a8u_goMux_mux_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C5_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  C5_t go_15_goMux_choice_3_d;
  logic go_15_goMux_choice_3_r;
  Pointer_QTree_Int_t m1ae6_goMux_mux_d;
  logic m1ae6_goMux_mux_r;
  Pointer_QTree_Int_t m2ae7_goMux_mux_d;
  logic m2ae7_goMux_mux_r;
  Pointer_CTf_f_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_d;
  logic lizzieLet0_1_1QVal_Bool_r;
  \CTf''''''''_f''''''''_t  \go_17_1Lf''''''''_f''''''''sbos_d ;
  logic \go_17_1Lf''''''''_f''''''''sbos_r ;
  \CTf''''''''_f''''''''_t  lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  Go_t go_17_2_argbuf_d;
  logic go_17_2_argbuf_r;
  \TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_t  \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d ;
  logic \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_r ;
  CTf_f_t go_18_1Lf_fsbos_d;
  logic go_18_1Lf_fsbos_r;
  CTf_f_t lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  Go_t go_18_2_argbuf_d;
  logic go_18_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_t call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d;
  logic call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_r;
  C4_t go_19_goMux_choice_1_d;
  logic go_19_goMux_choice_1_r;
  C4_t go_19_goMux_choice_2_d;
  logic go_19_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r;
  Go_t go_2_argbuf_d;
  logic go_2_argbuf_r;
  C5_t go_20_goMux_choice_1_d;
  logic go_20_goMux_choice_1_r;
  C5_t go_20_goMux_choice_2_d;
  logic go_20_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf''''''''_f''''''''_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C16_t go_21_goMux_choice_1_d;
  logic go_21_goMux_choice_1_r;
  C16_t go_21_goMux_choice_2_d;
  logic go_21_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTf_f_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  TupGo___Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_Bool_1_d ;
  logic \$wnnzTupGo___Pointer_QTree_Bool_1_r ;
  QTree_Bool_t lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Pointer_QTree_Int_t q1aen_destruct_d;
  logic q1aen_destruct_r;
  Pointer_QTree_Int_t q2aeo_destruct_d;
  logic q2aeo_destruct_r;
  Pointer_QTree_Int_t q3aep_destruct_d;
  logic q3aep_destruct_r;
  Pointer_QTree_Int_t q4aeq_destruct_d;
  logic q4aeq_destruct_r;
  Int_t v1aee_destruct_d;
  logic v1aee_destruct_r;
  QTree_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  QTree_Int_t lizzieLet12_1QVal_Int_d;
  logic lizzieLet12_1QVal_Int_r;
  QTree_Int_t lizzieLet12_1QNode_Int_d;
  logic lizzieLet12_1QNode_Int_r;
  QTree_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Go_t lizzieLet12_3QNone_Int_d;
  logic lizzieLet12_3QNone_Int_r;
  Go_t lizzieLet12_3QVal_Int_d;
  logic lizzieLet12_3QVal_Int_r;
  Go_t lizzieLet12_3QNode_Int_d;
  logic lizzieLet12_3QNode_Int_r;
  Go_t lizzieLet12_3QError_Int_d;
  logic lizzieLet12_3QError_Int_r;
  Go_t lizzieLet12_3QError_Int_1_d;
  logic lizzieLet12_3QError_Int_1_r;
  Go_t lizzieLet12_3QError_Int_2_d;
  logic lizzieLet12_3QError_Int_2_r;
  QTree_Bool_t lizzieLet12_3QError_Int_1QError_Bool_d;
  logic lizzieLet12_3QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Go_t lizzieLet12_3QError_Int_2_argbuf_d;
  logic lizzieLet12_3QError_Int_2_argbuf_r;
  QTree_Int_t lizzieLet12_4QNone_Int_d;
  logic lizzieLet12_4QNone_Int_r;
  QTree_Int_t lizzieLet12_4QVal_Int_d;
  logic lizzieLet12_4QVal_Int_r;
  QTree_Int_t lizzieLet12_4QNode_Int_d;
  logic lizzieLet12_4QNode_Int_r;
  QTree_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  QTree_Int_t lizzieLet12_4QNode_Int_1_d;
  logic lizzieLet12_4QNode_Int_1_r;
  QTree_Int_t lizzieLet12_4QNode_Int_2_d;
  logic lizzieLet12_4QNode_Int_2_r;
  QTree_Int_t lizzieLet12_4QNode_Int_3_d;
  logic lizzieLet12_4QNode_Int_3_r;
  QTree_Int_t lizzieLet12_4QNode_Int_4_d;
  logic lizzieLet12_4QNode_Int_4_r;
  QTree_Int_t lizzieLet12_4QNode_Int_5_d;
  logic lizzieLet12_4QNode_Int_5_r;
  QTree_Int_t lizzieLet12_4QNode_Int_6_d;
  logic lizzieLet12_4QNode_Int_6_r;
  QTree_Int_t lizzieLet12_4QNode_Int_7_d;
  logic lizzieLet12_4QNode_Int_7_r;
  QTree_Int_t lizzieLet12_4QNode_Int_8_d;
  logic lizzieLet12_4QNode_Int_8_r;
  Pointer_QTree_Int_t t1aes_destruct_d;
  logic t1aes_destruct_r;
  Pointer_QTree_Int_t t2aet_destruct_d;
  logic t2aet_destruct_r;
  Pointer_QTree_Int_t t3aeu_destruct_d;
  logic t3aeu_destruct_r;
  Pointer_QTree_Int_t t4aev_destruct_d;
  logic t4aev_destruct_r;
  QTree_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  QTree_Int_t lizzieLet12_4QNode_Int_1QNode_Int_d;
  logic lizzieLet12_4QNode_Int_1QNode_Int_r;
  QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_r;
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_r;
  Go_t lizzieLet12_4QNode_Int_3QNode_Int_d;
  logic lizzieLet12_4QNode_Int_3QNode_Int_r;
  Go_t lizzieLet12_4QNode_Int_3QError_Int_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_r;
  Go_t lizzieLet12_4QNode_Int_3QError_Int_1_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet12_4QNode_Int_3QError_Int_2_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_2_r;
  QTree_Bool_t lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  Go_t lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_1_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_1_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_2_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_2_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_3_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_3_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_4_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_4_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_5_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_5_r;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_r ;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_r ;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_r ;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int8_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int8_r ;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_r;
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_1_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_2_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_2_r;
  QTree_Bool_t lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QNone_Int_d;
  logic lizzieLet12_4QNode_Int_4QNone_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QVal_Int_d;
  logic lizzieLet12_4QNode_Int_4QVal_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QNode_Int_d;
  logic lizzieLet12_4QNode_Int_4QNode_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QError_Int_d;
  logic lizzieLet12_4QNode_Int_4QError_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_r;
  CTf_f_t lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_d;
  logic lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_r;
  CTf_f_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_5QNone_Int_d;
  logic lizzieLet12_4QNode_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_5QNode_Int_d;
  logic lizzieLet12_4QNode_Int_5QNode_Int_r;
  Pointer_QTree_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_6QNone_Int_d;
  logic lizzieLet12_4QNode_Int_6QNone_Int_r;
  Pointer_QTree_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_6QNode_Int_d;
  logic lizzieLet12_4QNode_Int_6QNode_Int_r;
  Pointer_QTree_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_7QNone_Int_d;
  logic lizzieLet12_4QNode_Int_7QNone_Int_r;
  Pointer_QTree_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_7QNode_Int_d;
  logic lizzieLet12_4QNode_Int_7QNode_Int_r;
  Pointer_QTree_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNone_Int_d;
  logic lizzieLet12_4QNode_Int_8QNone_Int_r;
  Pointer_QTree_Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNode_Int_d;
  logic lizzieLet12_4QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet12_4QNone_Int_1_d;
  logic lizzieLet12_4QNone_Int_1_r;
  QTree_Int_t lizzieLet12_4QNone_Int_2_d;
  logic lizzieLet12_4QNone_Int_2_r;
  QTree_Int_t lizzieLet12_4QNone_Int_3_d;
  logic lizzieLet12_4QNone_Int_3_r;
  QTree_Int_t lizzieLet12_4QNone_Int_4_d;
  logic lizzieLet12_4QNone_Int_4_r;
  Pointer_QTree_Int_t tlaea_destruct_d;
  logic tlaea_destruct_r;
  Pointer_QTree_Int_t traeb_destruct_d;
  logic traeb_destruct_r;
  Pointer_QTree_Int_t blaec_destruct_d;
  logic blaec_destruct_r;
  Pointer_QTree_Int_t braed_destruct_d;
  logic braed_destruct_r;
  Int_t vae8_destruct_d;
  logic vae8_destruct_r;
  QTree_Int_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  QTree_Int_t lizzieLet12_4QNone_Int_1QVal_Int_d;
  logic lizzieLet12_4QNone_Int_1QVal_Int_r;
  QTree_Int_t lizzieLet12_4QNone_Int_1QNode_Int_d;
  logic lizzieLet12_4QNone_Int_1QNode_Int_r;
  QTree_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_r;
  Go_t lizzieLet12_4QNone_Int_3QVal_Int_d;
  logic lizzieLet12_4QNone_Int_3QVal_Int_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_r;
  Go_t lizzieLet12_4QNone_Int_3QError_Int_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_r;
  Go_t lizzieLet12_4QNone_Int_3QError_Int_1_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_1_r;
  Go_t lizzieLet12_4QNone_Int_3QError_Int_2_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_2_r;
  QTree_Bool_t lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_1_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_1_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_2_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_2_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_3_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_3_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_4_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_4_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_5_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_5_r;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_r ;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_r ;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_r ;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_r;
  TupGo___Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_r ;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_r;
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_1_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_1_r;
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_2_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_2_r;
  QTree_Bool_t lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_r;
  QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_r;
  C16_t go_21_goMux_choice_d;
  logic go_21_goMux_choice_r;
  Go_t go_21_goMux_data_d;
  logic go_21_goMux_data_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNone_Int_d;
  logic lizzieLet12_4QNone_Int_4QNone_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QVal_Int_d;
  logic lizzieLet12_4QNone_Int_4QVal_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNode_Int_d;
  logic lizzieLet12_4QNone_Int_4QNode_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QError_Int_d;
  logic lizzieLet12_4QNone_Int_4QError_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet12_4QVal_Int_1_d;
  logic lizzieLet12_4QVal_Int_1_r;
  QTree_Int_t lizzieLet12_4QVal_Int_2_d;
  logic lizzieLet12_4QVal_Int_2_r;
  QTree_Int_t lizzieLet12_4QVal_Int_3_d;
  logic lizzieLet12_4QVal_Int_3_r;
  QTree_Int_t lizzieLet12_4QVal_Int_4_d;
  logic lizzieLet12_4QVal_Int_4_r;
  QTree_Int_t lizzieLet12_4QVal_Int_5_d;
  logic lizzieLet12_4QVal_Int_5_r;
  Int_t vaeg_destruct_d;
  logic vaeg_destruct_r;
  QTree_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  QTree_Int_t lizzieLet12_4QVal_Int_1QVal_Int_d;
  logic lizzieLet12_4QVal_Int_1QVal_Int_r;
  QTree_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  QTree_Int_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Go_t lizzieLet12_4QVal_Int_3QNone_Int_d;
  logic lizzieLet12_4QVal_Int_3QNone_Int_r;
  Go_t lizzieLet12_4QVal_Int_3QVal_Int_d;
  logic lizzieLet12_4QVal_Int_3QVal_Int_r;
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_r;
  Go_t lizzieLet12_4QVal_Int_3QError_Int_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_r;
  Go_t lizzieLet12_4QVal_Int_3QError_Int_1_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet12_4QVal_Int_3QError_Int_2_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_2_r;
  QTree_Bool_t lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Go_t lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_1_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_2_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_2_r;
  QTree_Bool_t lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QNone_Int_d;
  logic lizzieLet12_4QVal_Int_4QNone_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QVal_Int_d;
  logic lizzieLet12_4QVal_Int_4QVal_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QNode_Int_d;
  logic lizzieLet12_4QVal_Int_4QNode_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QError_Int_d;
  logic lizzieLet12_4QVal_Int_4QError_Int_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_r;
  Int_t lizzieLet12_4QVal_Int_5QNone_Int_d;
  logic lizzieLet12_4QVal_Int_5QNone_Int_r;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_r;
  Int_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Int_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Int_t lizzieLet12_4QVal_Int_5QNone_Int_1_d;
  logic lizzieLet12_4QVal_Int_5QNone_Int_1_r;
  Int_t lizzieLet12_4QVal_Int_5QNone_Int_2_d;
  logic lizzieLet12_4QVal_Int_5QNone_Int_2_r;
  Int_t lizzieLet12_4QVal_Int_5QNone_Int_3_d;
  logic lizzieLet12_4QVal_Int_5QNone_Int_3_r;
  Int_t lizzieLet12_4QVal_Int_5QNone_Int_4_d;
  logic lizzieLet12_4QVal_Int_5QNone_Int_4_r;
  \Int#_t  xakK_2_destruct_d;
  logic xakK_2_destruct_r;
  Int_t \lizzieLet12_4QVal_Int_5QNone_Int_1I#_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_1I#_r ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_r ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_r ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_r ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_r ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_r ;
  \Int#_t  \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet23_1wild3XR_1_1_Eq_d;
  logic lizzieLet23_1wild3XR_1_1_Eq_r;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_3TupGo___Bool_1_d;
  logic boolConvert_3TupGo___Bool_1_r;
  Pointer_CTf_f_t \lizzieLet12_4QVal_Int_5QNone_Int_4I#_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_4I#_r ;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_1_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_1_r;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_2_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_2_r;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_3_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_3_r;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_4_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_4_r;
  Int_t lizzieLet12_4QVal_Int_5QVal_Int_5_d;
  logic lizzieLet12_4QVal_Int_5QVal_Int_5_r;
  \Int#_t  xakw_destruct_d;
  logic xakw_destruct_r;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_1I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_1I#_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_3I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_3I#_r ;
  Pointer_CTf_f_t \lizzieLet12_4QVal_Int_5QVal_Int_4I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_4I#_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_r ;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_r ;
  \Int#_t  yakA_destruct_d;
  logic yakA_destruct_r;
  Int_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_r ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_r ;
  \Int#_t  \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet28_1wild4XU_1_Eq_d;
  logic lizzieLet28_1wild4XU_1_Eq_r;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_4TupGo___Bool_1_d;
  logic boolConvert_4TupGo___Bool_1_r;
  Pointer_CTf_f_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_r ;
  \Int#_t  \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_r ;
  \Int#_t  \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_r ;
  Pointer_CTf_f_t lizzieLet12_5QNone_Int_d;
  logic lizzieLet12_5QNone_Int_r;
  Pointer_CTf_f_t lizzieLet12_5QVal_Int_d;
  logic lizzieLet12_5QVal_Int_r;
  Pointer_CTf_f_t lizzieLet12_5QNode_Int_d;
  logic lizzieLet12_5QNode_Int_r;
  Pointer_CTf_f_t lizzieLet12_5QError_Int_d;
  logic lizzieLet12_5QError_Int_r;
  Pointer_CTf_f_t lizzieLet12_5QError_Int_1_argbuf_d;
  logic lizzieLet12_5QError_Int_1_argbuf_r;
  Bool_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t lizzieLet17_1MyFalse_d;
  logic lizzieLet17_1MyFalse_r;
  Go_t lizzieLet17_1MyTrue_d;
  logic lizzieLet17_1MyTrue_r;
  Go_t lizzieLet17_1MyFalse_1_d;
  logic lizzieLet17_1MyFalse_1_r;
  Go_t lizzieLet17_1MyFalse_2_d;
  logic lizzieLet17_1MyFalse_2_r;
  Go_t lizzieLet17_1MyFalse_1_argbuf_d;
  logic lizzieLet17_1MyFalse_1_argbuf_r;
  TupGo_t \f''''''''1TupGo_1_d ;
  logic \f''''''''1TupGo_1_r ;
  Go_t lizzieLet17_1MyFalse_2_argbuf_d;
  logic lizzieLet17_1MyFalse_2_argbuf_r;
  Go_t lizzieLet17_1MyTrue_1_d;
  logic lizzieLet17_1MyTrue_1_r;
  Go_t lizzieLet17_1MyTrue_2_d;
  logic lizzieLet17_1MyTrue_2_r;
  QTree_Bool_t lizzieLet17_1MyTrue_1QNone_Bool_d;
  logic lizzieLet17_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet19_1_1_argbuf_d;
  logic lizzieLet19_1_1_argbuf_r;
  Go_t lizzieLet17_1MyTrue_2_argbuf_d;
  logic lizzieLet17_1MyTrue_2_argbuf_r;
  Pointer_CTf_f_t lizzieLet17_2MyFalse_d;
  logic lizzieLet17_2MyFalse_r;
  Pointer_CTf_f_t lizzieLet17_2MyTrue_d;
  logic lizzieLet17_2MyTrue_r;
  Pointer_CTf_f_t lizzieLet17_2MyFalse_1_argbuf_d;
  logic lizzieLet17_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet17_2MyTrue_1_argbuf_d;
  logic lizzieLet17_2MyTrue_1_argbuf_r;
  Pointer_QTree_Bool_t q1a84_destruct_d;
  logic q1a84_destruct_r;
  Pointer_QTree_Bool_t q2a85_destruct_d;
  logic q2a85_destruct_r;
  Pointer_QTree_Bool_t q3a86_destruct_d;
  logic q3a86_destruct_r;
  Pointer_QTree_Bool_t q4a87_destruct_d;
  logic q4a87_destruct_r;
  QTree_Bool_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  QTree_Bool_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  QTree_Bool_t lizzieLet1_1QNode_Bool_d;
  logic lizzieLet1_1QNode_Bool_r;
  QTree_Bool_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Go_t lizzieLet1_3QNone_Bool_d;
  logic lizzieLet1_3QNone_Bool_r;
  Go_t lizzieLet1_3QVal_Bool_d;
  logic lizzieLet1_3QVal_Bool_r;
  Go_t lizzieLet1_3QNode_Bool_d;
  logic lizzieLet1_3QNode_Bool_r;
  Go_t lizzieLet1_3QError_Bool_d;
  logic lizzieLet1_3QError_Bool_r;
  Go_t lizzieLet1_3QError_Bool_1_d;
  logic lizzieLet1_3QError_Bool_1_r;
  Go_t lizzieLet1_3QError_Bool_2_d;
  logic lizzieLet1_3QError_Bool_2_r;
  Go_t lizzieLet1_3QError_Bool_1_argbuf_d;
  logic lizzieLet1_3QError_Bool_1_argbuf_r;
  \Int#_t  lizzieLet1_3QError_Bool_1_argbuf_0_d;
  logic lizzieLet1_3QError_Bool_1_argbuf_0_r;
  \Int#_t  lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Go_t lizzieLet1_3QError_Bool_2_argbuf_d;
  logic lizzieLet1_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet1_3QNode_Bool_1_argbuf_d;
  logic lizzieLet1_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet1_3QNone_Bool_1_d;
  logic lizzieLet1_3QNone_Bool_1_r;
  Go_t lizzieLet1_3QNone_Bool_2_d;
  logic lizzieLet1_3QNone_Bool_2_r;
  Go_t lizzieLet1_3QNone_Bool_1_argbuf_d;
  logic lizzieLet1_3QNone_Bool_1_argbuf_r;
  \Int#_t  lizzieLet1_3QNone_Bool_1_argbuf_0_d;
  logic lizzieLet1_3QNone_Bool_1_argbuf_0_r;
  \Int#_t  lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet1_3QNone_Bool_2_argbuf_d;
  logic lizzieLet1_3QNone_Bool_2_argbuf_r;
  C4_t go_19_goMux_choice_d;
  logic go_19_goMux_choice_r;
  Go_t go_19_goMux_data_d;
  logic go_19_goMux_data_r;
  Go_t lizzieLet1_3QVal_Bool_1_d;
  logic lizzieLet1_3QVal_Bool_1_r;
  Go_t lizzieLet1_3QVal_Bool_2_d;
  logic lizzieLet1_3QVal_Bool_2_r;
  Go_t lizzieLet1_3QVal_Bool_1_argbuf_d;
  logic lizzieLet1_3QVal_Bool_1_argbuf_r;
  \Int#_t  lizzieLet1_3QVal_Bool_1_argbuf_1_d;
  logic lizzieLet1_3QVal_Bool_1_argbuf_1_r;
  \Int#_t  lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Go_t lizzieLet1_3QVal_Bool_2_argbuf_d;
  logic lizzieLet1_3QVal_Bool_2_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet1_4QNone_Bool_d;
  logic lizzieLet1_4QNone_Bool_r;
  Pointer_CT$wnnz_t lizzieLet1_4QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_r;
  Pointer_CT$wnnz_t lizzieLet1_4QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_r;
  Pointer_CT$wnnz_t lizzieLet1_4QError_Bool_d;
  logic lizzieLet1_4QError_Bool_r;
  Pointer_CT$wnnz_t lizzieLet1_4QError_Bool_1_argbuf_d;
  logic lizzieLet1_4QError_Bool_1_argbuf_r;
  CT$wnnz_t lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d;
  logic lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet1_4QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QNone_Bool_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet1_4QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_1_argbuf_r;
  Bool_t lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Go_t lizzieLet25_1MyFalse_d;
  logic lizzieLet25_1MyFalse_r;
  Go_t lizzieLet25_1MyTrue_d;
  logic lizzieLet25_1MyTrue_r;
  Go_t lizzieLet25_1MyFalse_1_d;
  logic lizzieLet25_1MyFalse_1_r;
  Go_t lizzieLet25_1MyFalse_2_d;
  logic lizzieLet25_1MyFalse_2_r;
  Go_t lizzieLet25_1MyFalse_1_argbuf_d;
  logic lizzieLet25_1MyFalse_1_argbuf_r;
  TupGo_t \f''''''''1TupGo3_d ;
  logic \f''''''''1TupGo3_r ;
  Go_t lizzieLet25_1MyFalse_2_argbuf_d;
  logic lizzieLet25_1MyFalse_2_argbuf_r;
  Go_t lizzieLet25_1MyTrue_1_d;
  logic lizzieLet25_1MyTrue_1_r;
  Go_t lizzieLet25_1MyTrue_2_d;
  logic lizzieLet25_1MyTrue_2_r;
  QTree_Bool_t lizzieLet25_1MyTrue_1QNone_Bool_d;
  logic lizzieLet25_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  Go_t lizzieLet25_1MyTrue_2_argbuf_d;
  logic lizzieLet25_1MyTrue_2_argbuf_r;
  Pointer_CTf_f_t lizzieLet25_2MyFalse_d;
  logic lizzieLet25_2MyFalse_r;
  Pointer_CTf_f_t lizzieLet25_2MyTrue_d;
  logic lizzieLet25_2MyTrue_r;
  Pointer_CTf_f_t lizzieLet25_2MyFalse_1_argbuf_d;
  logic lizzieLet25_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet25_2MyTrue_1_argbuf_d;
  logic lizzieLet25_2MyTrue_1_argbuf_r;
  Bool_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Go_t lizzieLet30_1MyFalse_d;
  logic lizzieLet30_1MyFalse_r;
  Go_t lizzieLet30_1MyTrue_d;
  logic lizzieLet30_1MyTrue_r;
  Go_t lizzieLet30_1MyFalse_1_d;
  logic lizzieLet30_1MyFalse_1_r;
  Go_t lizzieLet30_1MyFalse_2_d;
  logic lizzieLet30_1MyFalse_2_r;
  Go_t lizzieLet30_1MyFalse_1_argbuf_d;
  logic lizzieLet30_1MyFalse_1_argbuf_r;
  TupGo_t \f''''''''1TupGo4_d ;
  logic \f''''''''1TupGo4_r ;
  Go_t lizzieLet30_1MyFalse_2_argbuf_d;
  logic lizzieLet30_1MyFalse_2_argbuf_r;
  Go_t lizzieLet30_1MyTrue_1_d;
  logic lizzieLet30_1MyTrue_1_r;
  Go_t lizzieLet30_1MyTrue_2_d;
  logic lizzieLet30_1MyTrue_2_r;
  QTree_Bool_t lizzieLet30_1MyTrue_1QNone_Bool_d;
  logic lizzieLet30_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  Go_t lizzieLet30_1MyTrue_2_argbuf_d;
  logic lizzieLet30_1MyTrue_2_argbuf_r;
  Pointer_CTf_f_t lizzieLet30_2MyFalse_d;
  logic lizzieLet30_2MyFalse_r;
  Pointer_CTf_f_t lizzieLet30_2MyTrue_d;
  logic lizzieLet30_2MyTrue_r;
  Pointer_CTf_f_t lizzieLet30_2MyFalse_1_argbuf_d;
  logic lizzieLet30_2MyFalse_1_argbuf_r;
  Pointer_CTf_f_t lizzieLet30_2MyTrue_1_argbuf_d;
  logic lizzieLet30_2MyTrue_1_argbuf_r;
  Pointer_QTree_Int_t tlae2_destruct_d;
  logic tlae2_destruct_r;
  Pointer_QTree_Int_t trae3_destruct_d;
  logic trae3_destruct_r;
  Pointer_QTree_Int_t blae4_destruct_d;
  logic blae4_destruct_r;
  Pointer_QTree_Int_t brae5_destruct_d;
  logic brae5_destruct_r;
  Int_t va8v_destruct_d;
  logic va8v_destruct_r;
  QTree_Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  QTree_Int_t lizzieLet3_1QVal_Int_d;
  logic lizzieLet3_1QVal_Int_r;
  QTree_Int_t lizzieLet3_1QNode_Int_d;
  logic lizzieLet3_1QNode_Int_r;
  QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Go_t lizzieLet3_3QNone_Int_d;
  logic lizzieLet3_3QNone_Int_r;
  Go_t lizzieLet3_3QVal_Int_d;
  logic lizzieLet3_3QVal_Int_r;
  Go_t lizzieLet3_3QNode_Int_d;
  logic lizzieLet3_3QNode_Int_r;
  Go_t lizzieLet3_3QError_Int_d;
  logic lizzieLet3_3QError_Int_r;
  Go_t lizzieLet3_3QError_Int_1_d;
  logic lizzieLet3_3QError_Int_1_r;
  Go_t lizzieLet3_3QError_Int_2_d;
  logic lizzieLet3_3QError_Int_2_r;
  QTree_Bool_t lizzieLet3_3QError_Int_1QError_Bool_d;
  logic lizzieLet3_3QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Go_t lizzieLet3_3QError_Int_2_argbuf_d;
  logic lizzieLet3_3QError_Int_2_argbuf_r;
  Go_t lizzieLet3_3QNode_Int_1_argbuf_d;
  logic lizzieLet3_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet3_3QNone_Int_1_d;
  logic lizzieLet3_3QNone_Int_1_r;
  Go_t lizzieLet3_3QNone_Int_2_d;
  logic lizzieLet3_3QNone_Int_2_r;
  QTree_Bool_t lizzieLet3_3QNone_Int_1QNone_Bool_d;
  logic lizzieLet3_3QNone_Int_1QNone_Bool_r;
  QTree_Bool_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  Go_t lizzieLet3_3QNone_Int_2_argbuf_d;
  logic lizzieLet3_3QNone_Int_2_argbuf_r;
  C5_t go_20_goMux_choice_d;
  logic go_20_goMux_choice_r;
  Go_t go_20_goMux_data_d;
  logic go_20_goMux_data_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QNone_Int_d;
  logic lizzieLet3_4QNone_Int_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QVal_Int_d;
  logic lizzieLet3_4QVal_Int_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QNode_Int_d;
  logic lizzieLet3_4QNode_Int_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QError_Int_d;
  logic lizzieLet3_4QError_Int_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QError_Int_1_argbuf_d;
  logic lizzieLet3_4QError_Int_1_argbuf_r;
  \CTf''''''''_f''''''''_t  \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_d ;
  logic \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_r ;
  \CTf''''''''_f''''''''_t  lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QNone_Int_1_argbuf_d;
  logic lizzieLet3_4QNone_Int_1_argbuf_r;
  \Int#_t  wwspI_4_destruct_d;
  logic wwspI_4_destruct_r;
  \Int#_t  ww1Xqr_2_destruct_d;
  logic ww1Xqr_2_destruct_r;
  \Int#_t  ww2Xqu_1_destruct_d;
  logic ww2Xqu_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  \Int#_t  wwspI_3_destruct_d;
  logic wwspI_3_destruct_r;
  \Int#_t  ww1Xqr_1_destruct_d;
  logic ww1Xqr_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Bool_t q4a87_3_destruct_d;
  logic q4a87_3_destruct_r;
  \Int#_t  wwspI_2_destruct_d;
  logic wwspI_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Bool_t q4a87_2_destruct_d;
  logic q4a87_2_destruct_r;
  Pointer_QTree_Bool_t q3a86_2_destruct_d;
  logic q3a86_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_QTree_Bool_t q4a87_1_destruct_d;
  logic q4a87_1_destruct_r;
  Pointer_QTree_Bool_t q3a86_1_destruct_d;
  logic q3a86_1_destruct_r;
  Pointer_QTree_Bool_t q2a85_1_destruct_d;
  logic q2a85_1_destruct_r;
  CT$wnnz_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  CT$wnnz_t lizzieLet44_1Lcall_$wnnz3_d;
  logic lizzieLet44_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet44_1Lcall_$wnnz2_d;
  logic lizzieLet44_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet44_1Lcall_$wnnz1_d;
  logic lizzieLet44_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet44_1Lcall_$wnnz0_d;
  logic lizzieLet44_1Lcall_$wnnz0_r;
  Go_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Go_t lizzieLet44_3Lcall_$wnnz3_d;
  logic lizzieLet44_3Lcall_$wnnz3_r;
  Go_t lizzieLet44_3Lcall_$wnnz2_d;
  logic lizzieLet44_3Lcall_$wnnz2_r;
  Go_t lizzieLet44_3Lcall_$wnnz1_d;
  logic lizzieLet44_3Lcall_$wnnz1_r;
  Go_t lizzieLet44_3Lcall_$wnnz0_d;
  logic lizzieLet44_3Lcall_$wnnz0_r;
  Go_t lizzieLet44_3Lcall_$wnnz0_1_argbuf_d;
  logic lizzieLet44_3Lcall_$wnnz0_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_$wnnz1_1_argbuf_d;
  logic lizzieLet44_3Lcall_$wnnz1_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_$wnnz2_1_argbuf_d;
  logic lizzieLet44_3Lcall_$wnnz2_1_argbuf_r;
  Go_t lizzieLet44_3Lcall_$wnnz3_1_argbuf_d;
  logic lizzieLet44_3Lcall_$wnnz3_1_argbuf_r;
  \Int#_t  lizzieLet44_4L$wnnzsbos_d;
  logic lizzieLet44_4L$wnnzsbos_r;
  \Int#_t  lizzieLet44_4Lcall_$wnnz3_d;
  logic lizzieLet44_4Lcall_$wnnz3_r;
  \Int#_t  lizzieLet44_4Lcall_$wnnz2_d;
  logic lizzieLet44_4Lcall_$wnnz2_r;
  \Int#_t  lizzieLet44_4Lcall_$wnnz1_d;
  logic lizzieLet44_4Lcall_$wnnz1_r;
  \Int#_t  lizzieLet44_4Lcall_$wnnz0_d;
  logic lizzieLet44_4Lcall_$wnnz0_r;
  \Int#_t  lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_d;
  logic lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_d;
  logic lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_goConst_d;
  logic call_$wnnz_goConst_r;
  \Int#_t  \$wnnz_resbuf_d ;
  logic \$wnnz_resbuf_r ;
  CT$wnnz_t lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d;
  logic lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet45_1_argbuf_d;
  logic lizzieLet45_1_argbuf_r;
  Pointer_QTree_Bool_t es_1_2_destruct_d;
  logic es_1_2_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Int_t tlae2_3_destruct_d;
  logic tlae2_3_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Int_t tlae2_2_destruct_d;
  logic tlae2_2_destruct_r;
  Pointer_QTree_Int_t trae3_2_destruct_d;
  logic trae3_2_destruct_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Int_t tlae2_1_destruct_d;
  logic tlae2_1_destruct_r;
  Pointer_QTree_Int_t trae3_1_destruct_d;
  logic trae3_1_destruct_r;
  Pointer_QTree_Int_t blae4_1_destruct_d;
  logic blae4_1_destruct_r;
  \CTf''''''''_f''''''''_t  _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  \CTf''''''''_f''''''''_t  \lizzieLet48_1Lcall_f''''''''_f''''''''3_d ;
  logic \lizzieLet48_1Lcall_f''''''''_f''''''''3_r ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_1Lcall_f''''''''_f''''''''2_d ;
  logic \lizzieLet48_1Lcall_f''''''''_f''''''''2_r ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_1Lcall_f''''''''_f''''''''1_d ;
  logic \lizzieLet48_1Lcall_f''''''''_f''''''''1_r ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_1Lcall_f''''''''_f''''''''0_d ;
  logic \lizzieLet48_1Lcall_f''''''''_f''''''''0_r ;
  Go_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''3_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''3_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''2_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''2_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''1_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''1_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''0_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''0_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_r ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf''''''''_f''''''''sbos_d ;
  logic \lizzieLet48_4Lf''''''''_f''''''''sbos_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''3_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''3_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''2_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''2_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''1_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''1_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''0_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''0_r ;
  QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet52_1_argbuf_d;
  logic lizzieLet52_1_argbuf_r;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_r ;
  \CTf''''''''_f''''''''_t  lizzieLet51_1_argbuf_d;
  logic lizzieLet51_1_argbuf_r;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_r ;
  \CTf''''''''_f''''''''_t  lizzieLet50_1_argbuf_d;
  logic lizzieLet50_1_argbuf_r;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_r ;
  \CTf''''''''_f''''''''_t  lizzieLet49_1_argbuf_d;
  logic lizzieLet49_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_r ;
  Go_t \call_f''''''''_f''''''''_goConst_d ;
  logic \call_f''''''''_f''''''''_goConst_r ;
  Pointer_QTree_Bool_t es_10_destruct_d;
  logic es_10_destruct_r;
  Pointer_QTree_Bool_t es_11_1_destruct_d;
  logic es_11_1_destruct_r;
  Pointer_QTree_Bool_t es_12_2_destruct_d;
  logic es_12_2_destruct_r;
  Pointer_CTf_f_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Bool_t es_11_destruct_d;
  logic es_11_destruct_r;
  Pointer_QTree_Bool_t es_12_1_destruct_d;
  logic es_12_1_destruct_r;
  Pointer_CTf_f_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t q1aen_3_destruct_d;
  logic q1aen_3_destruct_r;
  Pointer_QTree_Int_t t1aes_3_destruct_d;
  logic t1aes_3_destruct_r;
  Pointer_QTree_Bool_t es_12_destruct_d;
  logic es_12_destruct_r;
  Pointer_CTf_f_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t q1aen_2_destruct_d;
  logic q1aen_2_destruct_r;
  Pointer_QTree_Int_t t1aes_2_destruct_d;
  logic t1aes_2_destruct_r;
  Pointer_QTree_Int_t q2aeo_2_destruct_d;
  logic q2aeo_2_destruct_r;
  Pointer_QTree_Int_t t2aet_2_destruct_d;
  logic t2aet_2_destruct_r;
  Pointer_CTf_f_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t q1aen_1_destruct_d;
  logic q1aen_1_destruct_r;
  Pointer_QTree_Int_t t1aes_1_destruct_d;
  logic t1aes_1_destruct_r;
  Pointer_QTree_Int_t q2aeo_1_destruct_d;
  logic q2aeo_1_destruct_r;
  Pointer_QTree_Int_t t2aet_1_destruct_d;
  logic t2aet_1_destruct_r;
  Pointer_QTree_Int_t q3aep_1_destruct_d;
  logic q3aep_1_destruct_r;
  Pointer_QTree_Int_t t3aeu_1_destruct_d;
  logic t3aeu_1_destruct_r;
  CTf_f_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  CTf_f_t lizzieLet53_1Lcall_f_f3_d;
  logic lizzieLet53_1Lcall_f_f3_r;
  CTf_f_t lizzieLet53_1Lcall_f_f2_d;
  logic lizzieLet53_1Lcall_f_f2_r;
  CTf_f_t lizzieLet53_1Lcall_f_f1_d;
  logic lizzieLet53_1Lcall_f_f1_r;
  CTf_f_t lizzieLet53_1Lcall_f_f0_d;
  logic lizzieLet53_1Lcall_f_f0_r;
  Go_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Go_t lizzieLet53_3Lcall_f_f3_d;
  logic lizzieLet53_3Lcall_f_f3_r;
  Go_t lizzieLet53_3Lcall_f_f2_d;
  logic lizzieLet53_3Lcall_f_f2_r;
  Go_t lizzieLet53_3Lcall_f_f1_d;
  logic lizzieLet53_3Lcall_f_f1_r;
  Go_t lizzieLet53_3Lcall_f_f0_d;
  logic lizzieLet53_3Lcall_f_f0_r;
  Go_t lizzieLet53_3Lcall_f_f0_1_argbuf_d;
  logic lizzieLet53_3Lcall_f_f0_1_argbuf_r;
  Go_t lizzieLet53_3Lcall_f_f1_1_argbuf_d;
  logic lizzieLet53_3Lcall_f_f1_1_argbuf_r;
  Go_t lizzieLet53_3Lcall_f_f2_1_argbuf_d;
  logic lizzieLet53_3Lcall_f_f2_1_argbuf_r;
  Go_t lizzieLet53_3Lcall_f_f3_1_argbuf_d;
  logic lizzieLet53_3Lcall_f_f3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lf_fsbos_d;
  logic lizzieLet53_4Lf_fsbos_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lcall_f_f3_d;
  logic lizzieLet53_4Lcall_f_f3_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lcall_f_f2_d;
  logic lizzieLet53_4Lcall_f_f2_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lcall_f_f1_d;
  logic lizzieLet53_4Lcall_f_f1_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lcall_f_f0_d;
  logic lizzieLet53_4Lcall_f_f0_r;
  QTree_Bool_t lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_d;
  logic lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_r;
  QTree_Bool_t lizzieLet57_1_argbuf_d;
  logic lizzieLet57_1_argbuf_r;
  CTf_f_t lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_d;
  logic lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_r;
  CTf_f_t lizzieLet56_1_argbuf_d;
  logic lizzieLet56_1_argbuf_r;
  CTf_f_t lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_d;
  logic lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_r;
  CTf_f_t lizzieLet55_1_argbuf_d;
  logic lizzieLet55_1_argbuf_r;
  CTf_f_t lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_d;
  logic lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_r;
  CTf_f_t lizzieLet54_1_argbuf_d;
  logic lizzieLet54_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_d;
  logic lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_d;
  logic lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_r;
  Go_t call_f_f_goConst_d;
  logic call_f_f_goConst_r;
  Pointer_QTree_Bool_t f_f_resbuf_d;
  logic f_f_resbuf_r;
  Bool_t lizzieLet6_1_argbuf_d;
  logic lizzieLet6_1_argbuf_r;
  Go_t lizzieLet7_1MyFalse_d;
  logic lizzieLet7_1MyFalse_r;
  Go_t lizzieLet7_1MyTrue_d;
  logic lizzieLet7_1MyTrue_r;
  Go_t lizzieLet7_1MyFalse_1_d;
  logic lizzieLet7_1MyFalse_1_r;
  Go_t lizzieLet7_1MyFalse_2_d;
  logic lizzieLet7_1MyFalse_2_r;
  Go_t lizzieLet7_1MyFalse_1_argbuf_d;
  logic lizzieLet7_1MyFalse_1_argbuf_r;
  TupGo_t \f''''''''1TupGo2_d ;
  logic \f''''''''1TupGo2_r ;
  Go_t lizzieLet7_1MyFalse_2_argbuf_d;
  logic lizzieLet7_1MyFalse_2_argbuf_r;
  Go_t lizzieLet7_1MyTrue_1_d;
  logic lizzieLet7_1MyTrue_1_r;
  Go_t lizzieLet7_1MyTrue_2_d;
  logic lizzieLet7_1MyTrue_2_r;
  QTree_Bool_t lizzieLet7_1MyTrue_1QNone_Bool_d;
  logic lizzieLet7_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t lizzieLet7_1MyTrue_2_argbuf_d;
  logic lizzieLet7_1MyTrue_2_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyFalse_d;
  logic lizzieLet7_2MyFalse_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyTrue_d;
  logic lizzieLet7_2MyTrue_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyFalse_1_argbuf_d;
  logic lizzieLet7_2MyFalse_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyTrue_1_argbuf_d;
  logic lizzieLet7_2MyTrue_1_argbuf_r;
  Pointer_QTree_Int_t m1ae6_1_argbuf_d;
  logic m1ae6_1_argbuf_r;
  Pointer_QTree_Int_t m2ae7_1_argbuf_d;
  logic m2ae7_1_argbuf_r;
  Pointer_QTree_Bool_t q1a84_1_argbuf_d;
  logic q1a84_1_argbuf_r;
  Pointer_QTree_Int_t q1aen_3_1_argbuf_d;
  logic q1aen_3_1_argbuf_r;
  Pointer_QTree_Bool_t q2a85_1_1_argbuf_d;
  logic q2a85_1_1_argbuf_r;
  Pointer_QTree_Int_t q2aeo_2_1_argbuf_d;
  logic q2aeo_2_1_argbuf_r;
  Pointer_QTree_Bool_t q3a86_2_1_argbuf_d;
  logic q3a86_2_1_argbuf_r;
  Pointer_QTree_Int_t q3aep_1_1_argbuf_d;
  logic q3aep_1_1_argbuf_r;
  Pointer_QTree_Bool_t q4a87_3_1_argbuf_d;
  logic q4a87_3_1_argbuf_r;
  Pointer_QTree_Int_t q4a8u_1_argbuf_d;
  logic q4a8u_1_argbuf_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_t lizzieLet44_1_d;
  logic lizzieLet44_1_r;
  CT$wnnz_t lizzieLet44_2_d;
  logic lizzieLet44_2_r;
  CT$wnnz_t lizzieLet44_3_d;
  logic lizzieLet44_3_r;
  CT$wnnz_t lizzieLet44_4_d;
  logic lizzieLet44_4_r;
  \CTf''''''''_f''''''''_t  \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_r ;
  \CTf''''''''_f''''''''_t  lizzieLet48_1_d;
  logic lizzieLet48_1_r;
  \CTf''''''''_f''''''''_t  lizzieLet48_2_d;
  logic lizzieLet48_2_r;
  \CTf''''''''_f''''''''_t  lizzieLet48_3_d;
  logic lizzieLet48_3_r;
  \CTf''''''''_f''''''''_t  lizzieLet48_4_d;
  logic lizzieLet48_4_r;
  CTf_f_t readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_r;
  CTf_f_t lizzieLet53_1_d;
  logic lizzieLet53_1_r;
  CTf_f_t lizzieLet53_2_d;
  logic lizzieLet53_2_r;
  CTf_f_t lizzieLet53_3_d;
  logic lizzieLet53_3_r;
  CTf_f_t lizzieLet53_4_d;
  logic lizzieLet53_4_r;
  QTree_Bool_t readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d;
  logic readPointer_QTree_BoolwspF_1_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet1_1_d;
  logic lizzieLet1_1_r;
  QTree_Bool_t lizzieLet1_2_d;
  logic lizzieLet1_2_r;
  QTree_Bool_t lizzieLet1_3_d;
  logic lizzieLet1_3_r;
  QTree_Bool_t lizzieLet1_4_d;
  logic lizzieLet1_4_r;
  QTree_Int_t readPointer_QTree_Intm1ae6_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1ae6_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet12_1_d;
  logic lizzieLet12_1_r;
  QTree_Int_t lizzieLet12_2_d;
  logic lizzieLet12_2_r;
  QTree_Int_t lizzieLet12_3_d;
  logic lizzieLet12_3_r;
  QTree_Int_t lizzieLet12_4_d;
  logic lizzieLet12_4_r;
  QTree_Int_t lizzieLet12_5_d;
  logic lizzieLet12_5_r;
  QTree_Int_t readPointer_QTree_Intm2ae7_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2ae7_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_rwb_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  QTree_Int_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  QTree_Int_t lizzieLet3_3_d;
  logic lizzieLet3_3_r;
  QTree_Int_t lizzieLet3_4_d;
  logic lizzieLet3_4_r;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  Pointer_CTf_f_t sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wnnz_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTf_f_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wnnz_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1aes_3_1_argbuf_d;
  logic t1aes_3_1_argbuf_r;
  Pointer_QTree_Int_t t2aet_2_1_argbuf_d;
  logic t2aet_2_1_argbuf_r;
  Pointer_QTree_Int_t t3aeu_1_1_argbuf_d;
  logic t3aeu_1_1_argbuf_r;
  Pointer_QTree_Int_t t4aev_1_argbuf_d;
  logic t4aev_1_argbuf_r;
  Pointer_QTree_Int_t tlae2_3_1_argbuf_d;
  logic tlae2_3_1_argbuf_r;
  Pointer_QTree_Int_t tlaea_1_argbuf_d;
  logic tlaea_1_argbuf_r;
  Pointer_QTree_Int_t trae3_2_1_argbuf_d;
  logic trae3_2_1_argbuf_r;
  Pointer_QTree_Int_t traeb_1_argbuf_d;
  logic traeb_1_argbuf_r;
  \Int#_t  xakK_destruct_d;
  logic xakK_destruct_r;
  Int_t \va8v_1I#_d ;
  logic \va8v_1I#_r ;
  Go_t \va8v_3I#_d ;
  logic \va8v_3I#_r ;
  Go_t \va8v_3I#_1_d ;
  logic \va8v_3I#_1_r ;
  Go_t \va8v_3I#_2_d ;
  logic \va8v_3I#_2_r ;
  Go_t \va8v_3I#_3_d ;
  logic \va8v_3I#_3_r ;
  Go_t \va8v_3I#_1_argbuf_d ;
  logic \va8v_3I#_1_argbuf_r ;
  \Int#_t  \va8v_3I#_1_argbuf_0_d ;
  logic \va8v_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet5_1wild2XE_1_Eq_d;
  logic lizzieLet5_1wild2XE_1_Eq_r;
  Go_t \va8v_3I#_2_argbuf_d ;
  logic \va8v_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  \Pointer_CTf''''''''_f''''''''_t  \va8v_4I#_d ;
  logic \va8v_4I#_r ;
  Int_t va8v_1_d;
  logic va8v_1_r;
  Int_t va8v_2_d;
  logic va8v_2_r;
  Int_t va8v_3_d;
  logic va8v_3_r;
  Int_t va8v_4_d;
  logic va8v_4_r;
  \Int#_t  xakK_1_destruct_d;
  logic xakK_1_destruct_r;
  Int_t \vae8_1I#_d ;
  logic \vae8_1I#_r ;
  Go_t \vae8_3I#_d ;
  logic \vae8_3I#_r ;
  Go_t \vae8_3I#_1_d ;
  logic \vae8_3I#_1_r ;
  Go_t \vae8_3I#_2_d ;
  logic \vae8_3I#_2_r ;
  Go_t \vae8_3I#_3_d ;
  logic \vae8_3I#_3_r ;
  Go_t \vae8_3I#_1_argbuf_d ;
  logic \vae8_3I#_1_argbuf_r ;
  \Int#_t  \vae8_3I#_1_argbuf_0_d ;
  logic \vae8_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet15_1wild3XR_1_Eq_d;
  logic lizzieLet15_1wild3XR_1_Eq_r;
  Go_t \vae8_3I#_2_argbuf_d ;
  logic \vae8_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_2TupGo___Bool_1_d;
  logic boolConvert_2TupGo___Bool_1_r;
  Pointer_CTf_f_t \vae8_4I#_d ;
  logic \vae8_4I#_r ;
  Int_t vae8_1_d;
  logic vae8_1_r;
  Int_t vae8_2_d;
  logic vae8_2_r;
  Int_t vae8_3_d;
  logic vae8_3_r;
  Int_t vae8_4_d;
  logic vae8_4_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet2_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet45_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet46_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet47_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_r ;
  \Pointer_CTf''''''''_f''''''''_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_rwb_d;
  logic writeCTf_flizzieLet38_1_argbuf_rwb_r;
  Pointer_CTf_f_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_rwb_d;
  logic writeCTf_flizzieLet43_1_argbuf_rwb_r;
  Pointer_CTf_f_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_rwb_d;
  logic writeCTf_flizzieLet54_1_argbuf_rwb_r;
  Pointer_CTf_f_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_rwb_d;
  logic writeCTf_flizzieLet55_1_argbuf_rwb_r;
  Pointer_CTf_f_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_rwb_d;
  logic writeCTf_flizzieLet56_1_argbuf_rwb_r;
  Pointer_CTf_f_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet19_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet20_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet21_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet27_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet32_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet41_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet41_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Bool_t wspF_1_1_argbuf_d;
  logic wspF_1_1_argbuf_r;
  CT$wnnz_t lizzieLet46_1_argbuf_d;
  logic lizzieLet46_1_argbuf_r;
  CT$wnnz_t wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d;
  logic wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  CT$wnnz_t wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  logic wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r;
  \Int#_t  es_6_1_1ww2Xqu_1_1_Add32_d;
  logic es_6_1_1ww2Xqu_1_1_Add32_r;
  \Int#_t  wwspI_4_1ww1Xqr_2_1_Add32_d;
  logic wwspI_4_1ww1Xqr_2_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go__3,Go),
                                (go__4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go)] */
  logic [9:0] sourceGo_emitted;
  logic [9:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go__3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go__4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign sourceGo_done = (sourceGo_emitted | ({go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go__4_d[0],
                                               go__3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go__4_r,
                                                             go__3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 10'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 10'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,Lit 0) : (go__3,Go) > (initHP_CT$wnnz,Word16#) */
  assign initHP_CT$wnnz_d = {16'd0, go__3_d[0]};
  assign go__3_r = initHP_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz1,Go) > (incrHP_CT$wnnz,Word16#) */
  assign incrHP_CT$wnnz_d = {16'd1, incrHP_CT$wnnz1_d[0]};
  assign incrHP_CT$wnnz1_r = incrHP_CT$wnnz_r;
  
  /* merge (Ty Go) : [(go__4,Go),
                 (incrHP_CT$wnnz2,Go)] > (incrHP_mergeCT$wnnz,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_selected;
  logic [1:0] incrHP_mergeCT$wnnz_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_select))
        incrHP_mergeCT$wnnz_selected = incrHP_mergeCT$wnnz_select;
      else
        if (go__4_d[0]) incrHP_mergeCT$wnnz_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz2_d[0])
          incrHP_mergeCT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_select <= (incrHP_mergeCT$wnnz_r ? 2'd0 :
                                     incrHP_mergeCT$wnnz_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_selected[0])
      incrHP_mergeCT$wnnz_d = go__4_d;
    else if (incrHP_mergeCT$wnnz_selected[1])
      incrHP_mergeCT$wnnz_d = incrHP_CT$wnnz2_d;
    else incrHP_mergeCT$wnnz_d = 1'd0;
  assign {incrHP_CT$wnnz2_r,
          go__4_r} = (incrHP_mergeCT$wnnz_r ? incrHP_mergeCT$wnnz_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_buf,Go) > [(incrHP_CT$wnnz1,Go),
                                               (incrHP_CT$wnnz2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_buf_done;
  assign incrHP_CT$wnnz1_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[0]));
  assign incrHP_CT$wnnz2_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_buf_done = (incrHP_mergeCT$wnnz_buf_emitted | ({incrHP_CT$wnnz2_d[0],
                                                                             incrHP_CT$wnnz1_d[0]} & {incrHP_CT$wnnz2_r,
                                                                                                      incrHP_CT$wnnz1_r}));
  assign incrHP_mergeCT$wnnz_buf_r = (& incrHP_mergeCT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_buf_emitted <= (incrHP_mergeCT$wnnz_buf_r ? 2'd0 :
                                          incrHP_mergeCT$wnnz_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz,Word16#) (forkHP1_CT$wnnz,Word16#) > (addHP_CT$wnnz,Word16#) */
  assign addHP_CT$wnnz_d = {(incrHP_CT$wnnz_d[16:1] + forkHP1_CT$wnnz_d[16:1]),
                            (incrHP_CT$wnnz_d[0] && forkHP1_CT$wnnz_d[0])};
  assign {incrHP_CT$wnnz_r,
          forkHP1_CT$wnnz_r} = {2 {(addHP_CT$wnnz_r && addHP_CT$wnnz_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz,Word16#),
                      (addHP_CT$wnnz,Word16#)] > (mergeHP_CT$wnnz,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_selected;
  logic [1:0] mergeHP_CT$wnnz_select;
  always_comb
    begin
      mergeHP_CT$wnnz_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_select))
        mergeHP_CT$wnnz_selected = mergeHP_CT$wnnz_select;
      else
        if (initHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_select <= 2'd0;
    else
      mergeHP_CT$wnnz_select <= (mergeHP_CT$wnnz_r ? 2'd0 :
                                 mergeHP_CT$wnnz_selected);
  always_comb
    if (mergeHP_CT$wnnz_selected[0])
      mergeHP_CT$wnnz_d = initHP_CT$wnnz_d;
    else if (mergeHP_CT$wnnz_selected[1])
      mergeHP_CT$wnnz_d = addHP_CT$wnnz_d;
    else mergeHP_CT$wnnz_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_r,
          initHP_CT$wnnz_r} = (mergeHP_CT$wnnz_r ? mergeHP_CT$wnnz_selected :
                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz,Go) > (incrHP_mergeCT$wnnz_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_bufchan_d;
  logic incrHP_mergeCT$wnnz_bufchan_r;
  assign incrHP_mergeCT$wnnz_r = ((! incrHP_mergeCT$wnnz_bufchan_d[0]) || incrHP_mergeCT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_r)
        incrHP_mergeCT$wnnz_bufchan_d <= incrHP_mergeCT$wnnz_d;
  Go_t incrHP_mergeCT$wnnz_bufchan_buf;
  assign incrHP_mergeCT$wnnz_bufchan_r = (! incrHP_mergeCT$wnnz_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_buf_d = (incrHP_mergeCT$wnnz_bufchan_buf[0] ? incrHP_mergeCT$wnnz_bufchan_buf :
                                      incrHP_mergeCT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_buf_r && incrHP_mergeCT$wnnz_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_buf_r) && (! incrHP_mergeCT$wnnz_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_bufchan_buf <= incrHP_mergeCT$wnnz_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz,Word16#) > (mergeHP_CT$wnnz_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_bufchan_d;
  logic mergeHP_CT$wnnz_bufchan_r;
  assign mergeHP_CT$wnnz_r = ((! mergeHP_CT$wnnz_bufchan_d[0]) || mergeHP_CT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_r)
        mergeHP_CT$wnnz_bufchan_d <= mergeHP_CT$wnnz_d;
  \Word16#_t  mergeHP_CT$wnnz_bufchan_buf;
  assign mergeHP_CT$wnnz_bufchan_r = (! mergeHP_CT$wnnz_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_buf_d = (mergeHP_CT$wnnz_bufchan_buf[0] ? mergeHP_CT$wnnz_bufchan_buf :
                                  mergeHP_CT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_buf_r && mergeHP_CT$wnnz_bufchan_buf[0]))
        mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_buf_r) && (! mergeHP_CT$wnnz_bufchan_buf[0])))
        mergeHP_CT$wnnz_bufchan_buf <= mergeHP_CT$wnnz_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_buf,Word16#) > [(forkHP1_CT$wnnz,Word16#),
                                                     (forkHP1_CT$wnn2,Word16#),
                                                     (forkHP1_CT$wnn3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_buf_done;
  assign forkHP1_CT$wnnz_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[0]))};
  assign forkHP1_CT$wnn2_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[1]))};
  assign forkHP1_CT$wnn3_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_buf_done = (mergeHP_CT$wnnz_buf_emitted | ({forkHP1_CT$wnn3_d[0],
                                                                     forkHP1_CT$wnn2_d[0],
                                                                     forkHP1_CT$wnnz_d[0]} & {forkHP1_CT$wnn3_r,
                                                                                              forkHP1_CT$wnn2_r,
                                                                                              forkHP1_CT$wnnz_r}));
  assign mergeHP_CT$wnnz_buf_r = (& mergeHP_CT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_buf_emitted <= (mergeHP_CT$wnnz_buf_r ? 3'd0 :
                                      mergeHP_CT$wnnz_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz) : [(dconReadIn_CT$wnnz,MemIn_CT$wnnz),
                                (dconWriteIn_CT$wnnz,MemIn_CT$wnnz)] > (memMergeChoice_CT$wnnz,C2) (memMergeIn_CT$wnnz,MemIn_CT$wnnz) */
  logic [1:0] dconReadIn_CT$wnnz_select_d;
  assign dconReadIn_CT$wnnz_select_d = ((| dconReadIn_CT$wnnz_select_q) ? dconReadIn_CT$wnnz_select_q :
                                        (dconReadIn_CT$wnnz_d[0] ? 2'd1 :
                                         (dconWriteIn_CT$wnnz_d[0] ? 2'd2 :
                                          2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_select_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                      dconReadIn_CT$wnnz_select_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_emit_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                    dconReadIn_CT$wnnz_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_d;
  assign dconReadIn_CT$wnnz_emit_d = (dconReadIn_CT$wnnz_emit_q | ({memMergeChoice_CT$wnnz_d[0],
                                                                    memMergeIn_CT$wnnz_d[0]} & {memMergeChoice_CT$wnnz_r,
                                                                                                memMergeIn_CT$wnnz_r}));
  logic dconReadIn_CT$wnnz_done;
  assign dconReadIn_CT$wnnz_done = (& dconReadIn_CT$wnnz_emit_d);
  assign {dconWriteIn_CT$wnnz_r,
          dconReadIn_CT$wnnz_r} = (dconReadIn_CT$wnnz_done ? dconReadIn_CT$wnnz_select_d :
                                   2'd0);
  assign memMergeIn_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconReadIn_CT$wnnz_d :
                                 ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconWriteIn_CT$wnnz_d :
                                  {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C1_2_dc(1'd1) :
                                     ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C2_2_dc(1'd1) :
                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz,
      Ty MemOut_CT$wnnz) : (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) > (memOut_CT$wnnz,MemOut_CT$wnnz) */
  logic [114:0] memMergeIn_CT$wnnz_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_dbuf_din;
  logic [114:0] memOut_CT$wnnz_q;
  logic memOut_CT$wnnz_valid;
  logic memMergeIn_CT$wnnz_dbuf_we;
  logic memOut_CT$wnnz_we;
  assign memMergeIn_CT$wnnz_dbuf_din = memMergeIn_CT$wnnz_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_dbuf_address = memMergeIn_CT$wnnz_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_dbuf_we = (memMergeIn_CT$wnnz_dbuf_d[1:1] && memMergeIn_CT$wnnz_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_we <= 1'd0;
        memOut_CT$wnnz_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_we <= memMergeIn_CT$wnnz_dbuf_we;
        memOut_CT$wnnz_valid <= memMergeIn_CT$wnnz_dbuf_d[0];
        if (memMergeIn_CT$wnnz_dbuf_we)
          begin
            memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address] <= memMergeIn_CT$wnnz_dbuf_din;
            memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_din;
          end
        else
          memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address];
      end
  assign memOut_CT$wnnz_d = {memOut_CT$wnnz_q,
                             memOut_CT$wnnz_we,
                             memOut_CT$wnnz_valid};
  assign memMergeIn_CT$wnnz_dbuf_r = ((! memOut_CT$wnnz_valid) || memOut_CT$wnnz_r);
  logic [31:0] profiling_MemIn_CT$wnnz_read;
  logic [31:0] profiling_MemIn_CT$wnnz_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_write <= 0;
        profiling_MemIn_CT$wnnz_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_write <= (profiling_MemIn_CT$wnnz_write + 1);
      else
        if ((memOut_CT$wnnz_valid == 1'd1))
          profiling_MemIn_CT$wnnz_read <= (profiling_MemIn_CT$wnnz_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz) : (memMergeChoice_CT$wnnz,C2) (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) > [(memReadOut_CT$wnnz,MemOut_CT$wnnz),
                                                                                                (memWriteOut_CT$wnnz,MemOut_CT$wnnz)] */
  logic [1:0] memOut_CT$wnnz_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_d[0] && memOut_CT$wnnz_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_d[1:1])
        1'd0: memOut_CT$wnnz_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                 memOut_CT$wnnz_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                  memOut_CT$wnnz_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_dbuf_r = (| (memOut_CT$wnnz_dbuf_onehotd & {memWriteOut_CT$wnnz_r,
                                                                    memReadOut_CT$wnnz_r}));
  assign memMergeChoice_CT$wnnz_r = memOut_CT$wnnz_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) */
  assign memMergeIn_CT$wnnz_rbuf_r = ((! memMergeIn_CT$wnnz_dbuf_d[0]) || memMergeIn_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_rbuf_r)
        memMergeIn_CT$wnnz_dbuf_d <= memMergeIn_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) */
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_buf;
  assign memMergeIn_CT$wnnz_r = (! memMergeIn_CT$wnnz_buf[0]);
  assign memMergeIn_CT$wnnz_rbuf_d = (memMergeIn_CT$wnnz_buf[0] ? memMergeIn_CT$wnnz_buf :
                                      memMergeIn_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_rbuf_r && memMergeIn_CT$wnnz_buf[0]))
        memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_rbuf_r) && (! memMergeIn_CT$wnnz_buf[0])))
        memMergeIn_CT$wnnz_buf <= memMergeIn_CT$wnnz_d;
  
  /* dbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) > (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) */
  assign memOut_CT$wnnz_rbuf_r = ((! memOut_CT$wnnz_dbuf_d[0]) || memOut_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_rbuf_r)
        memOut_CT$wnnz_dbuf_d <= memOut_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz,MemOut_CT$wnnz) > (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) */
  MemOut_CT$wnnz_t memOut_CT$wnnz_buf;
  assign memOut_CT$wnnz_r = (! memOut_CT$wnnz_buf[0]);
  assign memOut_CT$wnnz_rbuf_d = (memOut_CT$wnnz_buf[0] ? memOut_CT$wnnz_buf :
                                  memOut_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_rbuf_r && memOut_CT$wnnz_buf[0]))
        memOut_CT$wnnz_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_rbuf_r) && (! memOut_CT$wnnz_buf[0])))
        memOut_CT$wnnz_buf <= memOut_CT$wnnz_d;
  
  /* destruct (Ty Pointer_CT$wnnz,
          Dcon Pointer_CT$wnnz) : (scfarg_0_1_argbuf,Pointer_CT$wnnz) > [(destructReadIn_CT$wnnz,Word16#)] */
  assign destructReadIn_CT$wnnz_d = {scfarg_0_1_argbuf_d[16:1],
                                     scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon ReadIn_CT$wnnz) : [(destructReadIn_CT$wnnz,Word16#)] > (dconReadIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconReadIn_CT$wnnz_d = ReadIn_CT$wnnz_dc((& {destructReadIn_CT$wnnz_d[0]}), destructReadIn_CT$wnnz_d);
  assign {destructReadIn_CT$wnnz_r} = {1 {(dconReadIn_CT$wnnz_r && dconReadIn_CT$wnnz_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz,
          Dcon ReadOut_CT$wnnz) : (memReadOut_CT$wnnz,MemOut_CT$wnnz) > [(readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz)] */
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_d[116:2],
                                                   memReadOut_CT$wnnz_d[0]};
  assign memReadOut_CT$wnnz_r = readPointer_CT$wnnzscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CT$wnnz) : [(lizzieLet0_1_argbuf,CT$wnnz),
                                (lizzieLet2_1_argbuf,CT$wnnz),
                                (lizzieLet45_1_argbuf,CT$wnnz),
                                (lizzieLet46_1_argbuf,CT$wnnz),
                                (lizzieLet47_1_argbuf,CT$wnnz)] > (writeMerge_choice_CT$wnnz,C5) (writeMerge_data_CT$wnnz,CT$wnnz) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet2_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet45_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet46_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet47_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_d[0],
                                                                      writeMerge_data_CT$wnnz_d[0]} & {writeMerge_choice_CT$wnnz_r,
                                                                                                       writeMerge_data_CT$wnnz_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet47_1_argbuf_r,
          lizzieLet46_1_argbuf_r,
          lizzieLet45_1_argbuf_r,
          lizzieLet2_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                      ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet2_1_argbuf_d :
                                       ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet45_1_argbuf_d :
                                        ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet46_1_argbuf_d :
                                         ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                          {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                        ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                         ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                          ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                           ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz) : (writeMerge_choice_CT$wnnz,C5) (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz) > [(writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet2_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet45_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet46_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet47_1_argbuf,Pointer_CT$wnnz)] */
  logic [4:0] demuxWriteResult_CT$wnnz_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_d[0] && demuxWriteResult_CT$wnnz_d[0]))
      unique case (writeMerge_choice_CT$wnnz_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_onehotd = 5'd0;
  assign writeCT$wnnzlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[0]};
  assign writeCT$wnnzlizzieLet2_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[1]};
  assign writeCT$wnnzlizzieLet45_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[2]};
  assign writeCT$wnnzlizzieLet46_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[3]};
  assign writeCT$wnnzlizzieLet47_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_r = (| (demuxWriteResult_CT$wnnz_onehotd & {writeCT$wnnzlizzieLet47_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet46_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet45_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet2_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_r = demuxWriteResult_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon WriteIn_CT$wnnz) : [(forkHP1_CT$wnn2,Word16#),
                               (writeMerge_data_CT$wnnz,CT$wnnz)] > (dconWriteIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconWriteIn_CT$wnnz_d = WriteIn_CT$wnnz_dc((& {forkHP1_CT$wnn2_d[0],
                                                        writeMerge_data_CT$wnnz_d[0]}), forkHP1_CT$wnn2_d, writeMerge_data_CT$wnnz_d);
  assign {forkHP1_CT$wnn2_r,
          writeMerge_data_CT$wnnz_r} = {2 {(dconWriteIn_CT$wnnz_r && dconWriteIn_CT$wnnz_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz,
      Dcon Pointer_CT$wnnz) : [(forkHP1_CT$wnn3,Word16#)] > (dconPtr_CT$wnnz,Pointer_CT$wnnz) */
  assign dconPtr_CT$wnnz_d = Pointer_CT$wnnz_dc((& {forkHP1_CT$wnn3_d[0]}), forkHP1_CT$wnn3_d);
  assign {forkHP1_CT$wnn3_r} = {1 {(dconPtr_CT$wnnz_r && dconPtr_CT$wnnz_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz,
       Ty Pointer_CT$wnnz) : (memWriteOut_CT$wnnz,MemOut_CT$wnnz) (dconPtr_CT$wnnz,Pointer_CT$wnnz) > [(_36,Pointer_CT$wnnz),
                                                                                                       (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz)] */
  logic [1:0] dconPtr_CT$wnnz_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_d[0] && dconPtr_CT$wnnz_d[0]))
      unique case (memWriteOut_CT$wnnz_d[1:1])
        1'd0: dconPtr_CT$wnnz_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_onehotd = 2'd0;
  assign _36_d = {dconPtr_CT$wnnz_d[16:1],
                  dconPtr_CT$wnnz_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_d = {dconPtr_CT$wnnz_d[16:1],
                                       dconPtr_CT$wnnz_onehotd[1]};
  assign dconPtr_CT$wnnz_r = (| (dconPtr_CT$wnnz_onehotd & {demuxWriteResult_CT$wnnz_r,
                                                            _36_r}));
  assign memWriteOut_CT$wnnz_r = dconPtr_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__5,Go) > (initHP_CTf''''''''_f'''''''',Word16#) */
  assign \initHP_CTf''''''''_f''''''''_d  = {16'd0, go__5_d[0]};
  assign go__5_r = \initHP_CTf''''''''_f''''''''_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf''''''''_f''''''''1,Go) > (incrHP_CTf''''''''_f'''''''',Word16#) */
  assign \incrHP_CTf''''''''_f''''''''_d  = {16'd1,
                                             \incrHP_CTf''''''''_f''''''''1_d [0]};
  assign \incrHP_CTf''''''''_f''''''''1_r  = \incrHP_CTf''''''''_f''''''''_r ;
  
  /* merge (Ty Go) : [(go__6,Go),
                 (incrHP_CTf''''''''_f''''''''2,Go)] > (incrHP_mergeCTf''''''''_f'''''''',Go) */
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_selected ;
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_select ;
  always_comb
    begin
      \incrHP_mergeCTf''''''''_f''''''''_selected  = 2'd0;
      if ((| \incrHP_mergeCTf''''''''_f''''''''_select ))
        \incrHP_mergeCTf''''''''_f''''''''_selected  = \incrHP_mergeCTf''''''''_f''''''''_select ;
      else
        if (go__6_d[0])
          \incrHP_mergeCTf''''''''_f''''''''_selected [0] = 1'd1;
        else if (\incrHP_CTf''''''''_f''''''''2_d [0])
          \incrHP_mergeCTf''''''''_f''''''''_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_select  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''_f''''''''_select  <= (\incrHP_mergeCTf''''''''_f''''''''_r  ? 2'd0 :
                                                     \incrHP_mergeCTf''''''''_f''''''''_selected );
  always_comb
    if (\incrHP_mergeCTf''''''''_f''''''''_selected [0])
      \incrHP_mergeCTf''''''''_f''''''''_d  = go__6_d;
    else if (\incrHP_mergeCTf''''''''_f''''''''_selected [1])
      \incrHP_mergeCTf''''''''_f''''''''_d  = \incrHP_CTf''''''''_f''''''''2_d ;
    else \incrHP_mergeCTf''''''''_f''''''''_d  = 1'd0;
  assign {\incrHP_CTf''''''''_f''''''''2_r ,
          go__6_r} = (\incrHP_mergeCTf''''''''_f''''''''_r  ? \incrHP_mergeCTf''''''''_f''''''''_selected  :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf''''''''_f''''''''_buf,Go) > [(incrHP_CTf''''''''_f''''''''1,Go),
                                                             (incrHP_CTf''''''''_f''''''''2,Go)] */
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf''''''''_f''''''''_buf_done ;
  assign \incrHP_CTf''''''''_f''''''''1_d  = (\incrHP_mergeCTf''''''''_f''''''''_buf_d [0] && (! \incrHP_mergeCTf''''''''_f''''''''_buf_emitted [0]));
  assign \incrHP_CTf''''''''_f''''''''2_d  = (\incrHP_mergeCTf''''''''_f''''''''_buf_d [0] && (! \incrHP_mergeCTf''''''''_f''''''''_buf_emitted [1]));
  assign \incrHP_mergeCTf''''''''_f''''''''_buf_done  = (\incrHP_mergeCTf''''''''_f''''''''_buf_emitted  | ({\incrHP_CTf''''''''_f''''''''2_d [0],
                                                                                                             \incrHP_CTf''''''''_f''''''''1_d [0]} & {\incrHP_CTf''''''''_f''''''''2_r ,
                                                                                                                                                      \incrHP_CTf''''''''_f''''''''1_r }));
  assign \incrHP_mergeCTf''''''''_f''''''''_buf_r  = (& \incrHP_mergeCTf''''''''_f''''''''_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf''''''''_f''''''''_buf_emitted  <= (\incrHP_mergeCTf''''''''_f''''''''_buf_r  ? 2'd0 :
                                                          \incrHP_mergeCTf''''''''_f''''''''_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf''''''''_f'''''''',Word16#) (forkHP1_CTf''''''''_f'''''''',Word16#) > (addHP_CTf''''''''_f'''''''',Word16#) */
  assign \addHP_CTf''''''''_f''''''''_d  = {(\incrHP_CTf''''''''_f''''''''_d [16:1] + \forkHP1_CTf''''''''_f''''''''_d [16:1]),
                                            (\incrHP_CTf''''''''_f''''''''_d [0] && \forkHP1_CTf''''''''_f''''''''_d [0])};
  assign {\incrHP_CTf''''''''_f''''''''_r ,
          \forkHP1_CTf''''''''_f''''''''_r } = {2 {(\addHP_CTf''''''''_f''''''''_r  && \addHP_CTf''''''''_f''''''''_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf''''''''_f'''''''',Word16#),
                      (addHP_CTf''''''''_f'''''''',Word16#)] > (mergeHP_CTf''''''''_f'''''''',Word16#) */
  logic [1:0] \mergeHP_CTf''''''''_f''''''''_selected ;
  logic [1:0] \mergeHP_CTf''''''''_f''''''''_select ;
  always_comb
    begin
      \mergeHP_CTf''''''''_f''''''''_selected  = 2'd0;
      if ((| \mergeHP_CTf''''''''_f''''''''_select ))
        \mergeHP_CTf''''''''_f''''''''_selected  = \mergeHP_CTf''''''''_f''''''''_select ;
      else
        if (\initHP_CTf''''''''_f''''''''_d [0])
          \mergeHP_CTf''''''''_f''''''''_selected [0] = 1'd1;
        else if (\addHP_CTf''''''''_f''''''''_d [0])
          \mergeHP_CTf''''''''_f''''''''_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_select  <= 2'd0;
    else
      \mergeHP_CTf''''''''_f''''''''_select  <= (\mergeHP_CTf''''''''_f''''''''_r  ? 2'd0 :
                                                 \mergeHP_CTf''''''''_f''''''''_selected );
  always_comb
    if (\mergeHP_CTf''''''''_f''''''''_selected [0])
      \mergeHP_CTf''''''''_f''''''''_d  = \initHP_CTf''''''''_f''''''''_d ;
    else if (\mergeHP_CTf''''''''_f''''''''_selected [1])
      \mergeHP_CTf''''''''_f''''''''_d  = \addHP_CTf''''''''_f''''''''_d ;
    else \mergeHP_CTf''''''''_f''''''''_d  = {16'd0, 1'd0};
  assign {\addHP_CTf''''''''_f''''''''_r ,
          \initHP_CTf''''''''_f''''''''_r } = (\mergeHP_CTf''''''''_f''''''''_r  ? \mergeHP_CTf''''''''_f''''''''_selected  :
                                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf''''''''_f'''''''',Go) > (incrHP_mergeCTf''''''''_f''''''''_buf,Go) */
  Go_t \incrHP_mergeCTf''''''''_f''''''''_bufchan_d ;
  logic \incrHP_mergeCTf''''''''_f''''''''_bufchan_r ;
  assign \incrHP_mergeCTf''''''''_f''''''''_r  = ((! \incrHP_mergeCTf''''''''_f''''''''_bufchan_d [0]) || \incrHP_mergeCTf''''''''_f''''''''_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf''''''''_f''''''''_r )
        \incrHP_mergeCTf''''''''_f''''''''_bufchan_d  <= \incrHP_mergeCTf''''''''_f''''''''_d ;
  Go_t \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf ;
  assign \incrHP_mergeCTf''''''''_f''''''''_bufchan_r  = (! \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf [0]);
  assign \incrHP_mergeCTf''''''''_f''''''''_buf_d  = (\incrHP_mergeCTf''''''''_f''''''''_bufchan_buf [0] ? \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf  :
                                                      \incrHP_mergeCTf''''''''_f''''''''_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf''''''''_f''''''''_buf_r  && \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf [0]))
        \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf''''''''_f''''''''_buf_r ) && (! \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf [0])))
        \incrHP_mergeCTf''''''''_f''''''''_bufchan_buf  <= \incrHP_mergeCTf''''''''_f''''''''_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf''''''''_f'''''''',Word16#) > (mergeHP_CTf''''''''_f''''''''_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_bufchan_d ;
  logic \mergeHP_CTf''''''''_f''''''''_bufchan_r ;
  assign \mergeHP_CTf''''''''_f''''''''_r  = ((! \mergeHP_CTf''''''''_f''''''''_bufchan_d [0]) || \mergeHP_CTf''''''''_f''''''''_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf''''''''_f''''''''_r )
        \mergeHP_CTf''''''''_f''''''''_bufchan_d  <= \mergeHP_CTf''''''''_f''''''''_d ;
  \Word16#_t  \mergeHP_CTf''''''''_f''''''''_bufchan_buf ;
  assign \mergeHP_CTf''''''''_f''''''''_bufchan_r  = (! \mergeHP_CTf''''''''_f''''''''_bufchan_buf [0]);
  assign \mergeHP_CTf''''''''_f''''''''_buf_d  = (\mergeHP_CTf''''''''_f''''''''_bufchan_buf [0] ? \mergeHP_CTf''''''''_f''''''''_bufchan_buf  :
                                                  \mergeHP_CTf''''''''_f''''''''_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf''''''''_f''''''''_buf_r  && \mergeHP_CTf''''''''_f''''''''_bufchan_buf [0]))
        \mergeHP_CTf''''''''_f''''''''_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf''''''''_f''''''''_buf_r ) && (! \mergeHP_CTf''''''''_f''''''''_bufchan_buf [0])))
        \mergeHP_CTf''''''''_f''''''''_bufchan_buf  <= \mergeHP_CTf''''''''_f''''''''_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf''''''''_f''''''''_buf,Word16#) > [(forkHP1_CTf''''''''_f'''''''',Word16#),
                                                                   (forkHP1_CTf''''''''_f'''''''2,Word16#),
                                                                   (forkHP1_CTf''''''''_f'''''''3,Word16#)] */
  logic [2:0] \mergeHP_CTf''''''''_f''''''''_buf_emitted ;
  logic [2:0] \mergeHP_CTf''''''''_f''''''''_buf_done ;
  assign \forkHP1_CTf''''''''_f''''''''_d  = {\mergeHP_CTf''''''''_f''''''''_buf_d [16:1],
                                              (\mergeHP_CTf''''''''_f''''''''_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_buf_emitted [0]))};
  assign \forkHP1_CTf''''''''_f'''''''2_d  = {\mergeHP_CTf''''''''_f''''''''_buf_d [16:1],
                                              (\mergeHP_CTf''''''''_f''''''''_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_buf_emitted [1]))};
  assign \forkHP1_CTf''''''''_f'''''''3_d  = {\mergeHP_CTf''''''''_f''''''''_buf_d [16:1],
                                              (\mergeHP_CTf''''''''_f''''''''_buf_d [0] && (! \mergeHP_CTf''''''''_f''''''''_buf_emitted [2]))};
  assign \mergeHP_CTf''''''''_f''''''''_buf_done  = (\mergeHP_CTf''''''''_f''''''''_buf_emitted  | ({\forkHP1_CTf''''''''_f'''''''3_d [0],
                                                                                                     \forkHP1_CTf''''''''_f'''''''2_d [0],
                                                                                                     \forkHP1_CTf''''''''_f''''''''_d [0]} & {\forkHP1_CTf''''''''_f'''''''3_r ,
                                                                                                                                              \forkHP1_CTf''''''''_f'''''''2_r ,
                                                                                                                                              \forkHP1_CTf''''''''_f''''''''_r }));
  assign \mergeHP_CTf''''''''_f''''''''_buf_r  = (& \mergeHP_CTf''''''''_f''''''''_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf''''''''_f''''''''_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf''''''''_f''''''''_buf_emitted  <= (\mergeHP_CTf''''''''_f''''''''_buf_r  ? 3'd0 :
                                                      \mergeHP_CTf''''''''_f''''''''_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf''''''''_f'''''''') : [(dconReadIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f''''''''),
                                              (dconWriteIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f'''''''')] > (memMergeChoice_CTf''''''''_f'''''''',C2) (memMergeIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f'''''''') */
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_select_d ;
  assign \dconReadIn_CTf''''''''_f''''''''_select_d  = ((| \dconReadIn_CTf''''''''_f''''''''_select_q ) ? \dconReadIn_CTf''''''''_f''''''''_select_q  :
                                                        (\dconReadIn_CTf''''''''_f''''''''_d [0] ? 2'd1 :
                                                         (\dconWriteIn_CTf''''''''_f''''''''_d [0] ? 2'd2 :
                                                          2'd0)));
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''_f''''''''_select_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''_f''''''''_select_q  <= (\dconReadIn_CTf''''''''_f''''''''_done  ? 2'd0 :
                                                      \dconReadIn_CTf''''''''_f''''''''_select_d );
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf''''''''_f''''''''_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf''''''''_f''''''''_emit_q  <= (\dconReadIn_CTf''''''''_f''''''''_done  ? 2'd0 :
                                                    \dconReadIn_CTf''''''''_f''''''''_emit_d );
  logic [1:0] \dconReadIn_CTf''''''''_f''''''''_emit_d ;
  assign \dconReadIn_CTf''''''''_f''''''''_emit_d  = (\dconReadIn_CTf''''''''_f''''''''_emit_q  | ({\memMergeChoice_CTf''''''''_f''''''''_d [0],
                                                                                                    \memMergeIn_CTf''''''''_f''''''''_d [0]} & {\memMergeChoice_CTf''''''''_f''''''''_r ,
                                                                                                                                                \memMergeIn_CTf''''''''_f''''''''_r }));
  logic \dconReadIn_CTf''''''''_f''''''''_done ;
  assign \dconReadIn_CTf''''''''_f''''''''_done  = (& \dconReadIn_CTf''''''''_f''''''''_emit_d );
  assign {\dconWriteIn_CTf''''''''_f''''''''_r ,
          \dconReadIn_CTf''''''''_f''''''''_r } = (\dconReadIn_CTf''''''''_f''''''''_done  ? \dconReadIn_CTf''''''''_f''''''''_select_d  :
                                                   2'd0);
  assign \memMergeIn_CTf''''''''_f''''''''_d  = ((\dconReadIn_CTf''''''''_f''''''''_select_d [0] && (! \dconReadIn_CTf''''''''_f''''''''_emit_q [0])) ? \dconReadIn_CTf''''''''_f''''''''_d  :
                                                 ((\dconReadIn_CTf''''''''_f''''''''_select_d [1] && (! \dconReadIn_CTf''''''''_f''''''''_emit_q [0])) ? \dconWriteIn_CTf''''''''_f''''''''_d  :
                                                  {84'd0, 1'd0}));
  assign \memMergeChoice_CTf''''''''_f''''''''_d  = ((\dconReadIn_CTf''''''''_f''''''''_select_d [0] && (! \dconReadIn_CTf''''''''_f''''''''_emit_q [1])) ? C1_2_dc(1'd1) :
                                                     ((\dconReadIn_CTf''''''''_f''''''''_select_d [1] && (! \dconReadIn_CTf''''''''_f''''''''_emit_q [1])) ? C2_2_dc(1'd1) :
                                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf''''''''_f'''''''',
      Ty MemOut_CTf''''''''_f'''''''') : (memMergeIn_CTf''''''''_f''''''''_dbuf,MemIn_CTf''''''''_f'''''''') > (memOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f'''''''') */
  logic [66:0] \memMergeIn_CTf''''''''_f''''''''_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf''''''''_f''''''''_dbuf_address ;
  logic [66:0] \memMergeIn_CTf''''''''_f''''''''_dbuf_din ;
  logic [66:0] \memOut_CTf''''''''_f''''''''_q ;
  logic \memOut_CTf''''''''_f''''''''_valid ;
  logic \memMergeIn_CTf''''''''_f''''''''_dbuf_we ;
  logic \memOut_CTf''''''''_f''''''''_we ;
  assign \memMergeIn_CTf''''''''_f''''''''_dbuf_din  = \memMergeIn_CTf''''''''_f''''''''_dbuf_d [84:18];
  assign \memMergeIn_CTf''''''''_f''''''''_dbuf_address  = \memMergeIn_CTf''''''''_f''''''''_dbuf_d [17:2];
  assign \memMergeIn_CTf''''''''_f''''''''_dbuf_we  = (\memMergeIn_CTf''''''''_f''''''''_dbuf_d [1:1] && \memMergeIn_CTf''''''''_f''''''''_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf''''''''_f''''''''_we  <= 1'd0;
        \memOut_CTf''''''''_f''''''''_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf''''''''_f''''''''_we  <= \memMergeIn_CTf''''''''_f''''''''_dbuf_we ;
        \memOut_CTf''''''''_f''''''''_valid  <= \memMergeIn_CTf''''''''_f''''''''_dbuf_d [0];
        if (\memMergeIn_CTf''''''''_f''''''''_dbuf_we )
          begin
            \memMergeIn_CTf''''''''_f''''''''_dbuf_mem [\memMergeIn_CTf''''''''_f''''''''_dbuf_address ] <= \memMergeIn_CTf''''''''_f''''''''_dbuf_din ;
            \memOut_CTf''''''''_f''''''''_q  <= \memMergeIn_CTf''''''''_f''''''''_dbuf_din ;
          end
        else
          \memOut_CTf''''''''_f''''''''_q  <= \memMergeIn_CTf''''''''_f''''''''_dbuf_mem [\memMergeIn_CTf''''''''_f''''''''_dbuf_address ];
      end
  assign \memOut_CTf''''''''_f''''''''_d  = {\memOut_CTf''''''''_f''''''''_q ,
                                             \memOut_CTf''''''''_f''''''''_we ,
                                             \memOut_CTf''''''''_f''''''''_valid };
  assign \memMergeIn_CTf''''''''_f''''''''_dbuf_r  = ((! \memOut_CTf''''''''_f''''''''_valid ) || \memOut_CTf''''''''_f''''''''_r );
  logic [31:0] \profiling_MemIn_CTf''''''''_f''''''''_read ;
  logic [31:0] \profiling_MemIn_CTf''''''''_f''''''''_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf''''''''_f''''''''_write  <= 0;
        \profiling_MemIn_CTf''''''''_f''''''''_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf''''''''_f''''''''_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf''''''''_f''''''''_write  <= (\profiling_MemIn_CTf''''''''_f''''''''_write  + 1);
      else
        if ((\memOut_CTf''''''''_f''''''''_valid  == 1'd1))
          \profiling_MemIn_CTf''''''''_f''''''''_read  <= (\profiling_MemIn_CTf''''''''_f''''''''_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf''''''''_f'''''''') : (memMergeChoice_CTf''''''''_f'''''''',C2) (memOut_CTf''''''''_f''''''''_dbuf,MemOut_CTf''''''''_f'''''''') > [(memReadOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f''''''''),
                                                                                                                                                        (memWriteOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f'''''''')] */
  logic [1:0] \memOut_CTf''''''''_f''''''''_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf''''''''_f''''''''_d [0] && \memOut_CTf''''''''_f''''''''_dbuf_d [0]))
      unique case (\memMergeChoice_CTf''''''''_f''''''''_d [1:1])
        1'd0: \memOut_CTf''''''''_f''''''''_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf''''''''_f''''''''_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf''''''''_f''''''''_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf''''''''_f''''''''_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf''''''''_f''''''''_d  = {\memOut_CTf''''''''_f''''''''_dbuf_d [68:1],
                                                 \memOut_CTf''''''''_f''''''''_dbuf_onehotd [0]};
  assign \memWriteOut_CTf''''''''_f''''''''_d  = {\memOut_CTf''''''''_f''''''''_dbuf_d [68:1],
                                                  \memOut_CTf''''''''_f''''''''_dbuf_onehotd [1]};
  assign \memOut_CTf''''''''_f''''''''_dbuf_r  = (| (\memOut_CTf''''''''_f''''''''_dbuf_onehotd  & {\memWriteOut_CTf''''''''_f''''''''_r ,
                                                                                                    \memReadOut_CTf''''''''_f''''''''_r }));
  assign \memMergeChoice_CTf''''''''_f''''''''_r  = \memOut_CTf''''''''_f''''''''_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf''''''''_f'''''''') : (memMergeIn_CTf''''''''_f''''''''_rbuf,MemIn_CTf''''''''_f'''''''') > (memMergeIn_CTf''''''''_f''''''''_dbuf,MemIn_CTf''''''''_f'''''''') */
  assign \memMergeIn_CTf''''''''_f''''''''_rbuf_r  = ((! \memMergeIn_CTf''''''''_f''''''''_dbuf_d [0]) || \memMergeIn_CTf''''''''_f''''''''_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''_f''''''''_dbuf_d  <= {84'd0, 1'd0};
    else
      if (\memMergeIn_CTf''''''''_f''''''''_rbuf_r )
        \memMergeIn_CTf''''''''_f''''''''_dbuf_d  <= \memMergeIn_CTf''''''''_f''''''''_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf''''''''_f'''''''') : (memMergeIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f'''''''') > (memMergeIn_CTf''''''''_f''''''''_rbuf,MemIn_CTf''''''''_f'''''''') */
  \MemIn_CTf''''''''_f''''''''_t  \memMergeIn_CTf''''''''_f''''''''_buf ;
  assign \memMergeIn_CTf''''''''_f''''''''_r  = (! \memMergeIn_CTf''''''''_f''''''''_buf [0]);
  assign \memMergeIn_CTf''''''''_f''''''''_rbuf_d  = (\memMergeIn_CTf''''''''_f''''''''_buf [0] ? \memMergeIn_CTf''''''''_f''''''''_buf  :
                                                      \memMergeIn_CTf''''''''_f''''''''_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf''''''''_f''''''''_buf  <= {84'd0, 1'd0};
    else
      if ((\memMergeIn_CTf''''''''_f''''''''_rbuf_r  && \memMergeIn_CTf''''''''_f''''''''_buf [0]))
        \memMergeIn_CTf''''''''_f''''''''_buf  <= {84'd0, 1'd0};
      else if (((! \memMergeIn_CTf''''''''_f''''''''_rbuf_r ) && (! \memMergeIn_CTf''''''''_f''''''''_buf [0])))
        \memMergeIn_CTf''''''''_f''''''''_buf  <= \memMergeIn_CTf''''''''_f''''''''_d ;
  
  /* dbuf (Ty MemOut_CTf''''''''_f'''''''') : (memOut_CTf''''''''_f''''''''_rbuf,MemOut_CTf''''''''_f'''''''') > (memOut_CTf''''''''_f''''''''_dbuf,MemOut_CTf''''''''_f'''''''') */
  assign \memOut_CTf''''''''_f''''''''_rbuf_r  = ((! \memOut_CTf''''''''_f''''''''_dbuf_d [0]) || \memOut_CTf''''''''_f''''''''_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''_f''''''''_dbuf_d  <= {68'd0, 1'd0};
    else
      if (\memOut_CTf''''''''_f''''''''_rbuf_r )
        \memOut_CTf''''''''_f''''''''_dbuf_d  <= \memOut_CTf''''''''_f''''''''_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf''''''''_f'''''''') : (memOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f'''''''') > (memOut_CTf''''''''_f''''''''_rbuf,MemOut_CTf''''''''_f'''''''') */
  \MemOut_CTf''''''''_f''''''''_t  \memOut_CTf''''''''_f''''''''_buf ;
  assign \memOut_CTf''''''''_f''''''''_r  = (! \memOut_CTf''''''''_f''''''''_buf [0]);
  assign \memOut_CTf''''''''_f''''''''_rbuf_d  = (\memOut_CTf''''''''_f''''''''_buf [0] ? \memOut_CTf''''''''_f''''''''_buf  :
                                                  \memOut_CTf''''''''_f''''''''_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf''''''''_f''''''''_buf  <= {68'd0, 1'd0};
    else
      if ((\memOut_CTf''''''''_f''''''''_rbuf_r  && \memOut_CTf''''''''_f''''''''_buf [0]))
        \memOut_CTf''''''''_f''''''''_buf  <= {68'd0, 1'd0};
      else if (((! \memOut_CTf''''''''_f''''''''_rbuf_r ) && (! \memOut_CTf''''''''_f''''''''_buf [0])))
        \memOut_CTf''''''''_f''''''''_buf  <= \memOut_CTf''''''''_f''''''''_d ;
  
  /* destruct (Ty Pointer_CTf''''''''_f'''''''',
          Dcon Pointer_CTf''''''''_f'''''''') : (scfarg_0_1_1_argbuf,Pointer_CTf''''''''_f'''''''') > [(destructReadIn_CTf''''''''_f'''''''',Word16#)] */
  assign \destructReadIn_CTf''''''''_f''''''''_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                     scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf''''''''_f''''''''_r ;
  
  /* dcon (Ty MemIn_CTf''''''''_f'''''''',
      Dcon ReadIn_CTf''''''''_f'''''''') : [(destructReadIn_CTf''''''''_f'''''''',Word16#)] > (dconReadIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f'''''''') */
  assign \dconReadIn_CTf''''''''_f''''''''_d  = \ReadIn_CTf''''''''_f''''''''_dc ((& {\destructReadIn_CTf''''''''_f''''''''_d [0]}), \destructReadIn_CTf''''''''_f''''''''_d );
  assign {\destructReadIn_CTf''''''''_f''''''''_r } = {1 {(\dconReadIn_CTf''''''''_f''''''''_r  && \dconReadIn_CTf''''''''_f''''''''_d [0])}};
  
  /* destruct (Ty MemOut_CTf''''''''_f'''''''',
          Dcon ReadOut_CTf''''''''_f'''''''') : (memReadOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f'''''''') > [(readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf,CTf''''''''_f'''''''')] */
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_d  = {\memReadOut_CTf''''''''_f''''''''_d [68:2],
                                                                     \memReadOut_CTf''''''''_f''''''''_d [0]};
  assign \memReadOut_CTf''''''''_f''''''''_r  = \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf''''''''_f'''''''') : [(lizzieLet10_1_argbuf,CTf''''''''_f''''''''),
                                        (lizzieLet42_1_argbuf,CTf''''''''_f''''''''),
                                        (lizzieLet49_1_argbuf,CTf''''''''_f''''''''),
                                        (lizzieLet50_1_argbuf,CTf''''''''_f''''''''),
                                        (lizzieLet51_1_argbuf,CTf''''''''_f'''''''')] > (writeMerge_choice_CTf''''''''_f'''''''',C5) (writeMerge_data_CTf''''''''_f'''''''',CTf''''''''_f'''''''') */
  logic [4:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet42_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet49_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet50_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet51_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 5'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({\writeMerge_choice_CTf''''''''_f''''''''_d [0],
                                                                        \writeMerge_data_CTf''''''''_f''''''''_d [0]} & {\writeMerge_choice_CTf''''''''_f''''''''_r ,
                                                                                                                         \writeMerge_data_CTf''''''''_f''''''''_r }));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {lizzieLet51_1_argbuf_r,
          lizzieLet50_1_argbuf_r,
          lizzieLet49_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf''''''''_f''''''''_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                                      ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                       ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet49_1_argbuf_d :
                                                        ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet50_1_argbuf_d :
                                                         ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet51_1_argbuf_d :
                                                          {67'd0, 1'd0})))));
  assign \writeMerge_choice_CTf''''''''_f''''''''_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                        ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                         ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                          ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                           ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf''''''''_f'''''''') : (writeMerge_choice_CTf''''''''_f'''''''',C5) (demuxWriteResult_CTf''''''''_f'''''''',Pointer_CTf''''''''_f'''''''') > [(writeCTf''''''''_f''''''''lizzieLet10_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                                                                                                                  (writeCTf''''''''_f''''''''lizzieLet42_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                                                                                                                  (writeCTf''''''''_f''''''''lizzieLet49_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                                                                                                                  (writeCTf''''''''_f''''''''lizzieLet50_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                                                                                                                  (writeCTf''''''''_f''''''''lizzieLet51_1_argbuf,Pointer_CTf''''''''_f'''''''')] */
  logic [4:0] \demuxWriteResult_CTf''''''''_f''''''''_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf''''''''_f''''''''_d [0] && \demuxWriteResult_CTf''''''''_f''''''''_d [0]))
      unique case (\writeMerge_choice_CTf''''''''_f''''''''_d [3:1])
        3'd0: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd16;
        default: \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf''''''''_f''''''''_onehotd  = 5'd0;
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_d [16:1],
                                                               \demuxWriteResult_CTf''''''''_f''''''''_onehotd [0]};
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_d [16:1],
                                                               \demuxWriteResult_CTf''''''''_f''''''''_onehotd [1]};
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_d [16:1],
                                                               \demuxWriteResult_CTf''''''''_f''''''''_onehotd [2]};
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_d [16:1],
                                                               \demuxWriteResult_CTf''''''''_f''''''''_onehotd [3]};
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_d  = {\demuxWriteResult_CTf''''''''_f''''''''_d [16:1],
                                                               \demuxWriteResult_CTf''''''''_f''''''''_onehotd [4]};
  assign \demuxWriteResult_CTf''''''''_f''''''''_r  = (| (\demuxWriteResult_CTf''''''''_f''''''''_onehotd  & {\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_r ,
                                                                                                              \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_r ,
                                                                                                              \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_r ,
                                                                                                              \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_r ,
                                                                                                              \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_r }));
  assign \writeMerge_choice_CTf''''''''_f''''''''_r  = \demuxWriteResult_CTf''''''''_f''''''''_r ;
  
  /* dcon (Ty MemIn_CTf''''''''_f'''''''',
      Dcon WriteIn_CTf''''''''_f'''''''') : [(forkHP1_CTf''''''''_f'''''''2,Word16#),
                                             (writeMerge_data_CTf''''''''_f'''''''',CTf''''''''_f'''''''')] > (dconWriteIn_CTf''''''''_f'''''''',MemIn_CTf''''''''_f'''''''') */
  assign \dconWriteIn_CTf''''''''_f''''''''_d  = \WriteIn_CTf''''''''_f''''''''_dc ((& {\forkHP1_CTf''''''''_f'''''''2_d [0],
                                                                                        \writeMerge_data_CTf''''''''_f''''''''_d [0]}), \forkHP1_CTf''''''''_f'''''''2_d , \writeMerge_data_CTf''''''''_f''''''''_d );
  assign {\forkHP1_CTf''''''''_f'''''''2_r ,
          \writeMerge_data_CTf''''''''_f''''''''_r } = {2 {(\dconWriteIn_CTf''''''''_f''''''''_r  && \dconWriteIn_CTf''''''''_f''''''''_d [0])}};
  
  /* dcon (Ty Pointer_CTf''''''''_f'''''''',
      Dcon Pointer_CTf''''''''_f'''''''') : [(forkHP1_CTf''''''''_f'''''''3,Word16#)] > (dconPtr_CTf''''''''_f'''''''',Pointer_CTf''''''''_f'''''''') */
  assign \dconPtr_CTf''''''''_f''''''''_d  = \Pointer_CTf''''''''_f''''''''_dc ((& {\forkHP1_CTf''''''''_f'''''''3_d [0]}), \forkHP1_CTf''''''''_f'''''''3_d );
  assign {\forkHP1_CTf''''''''_f'''''''3_r } = {1 {(\dconPtr_CTf''''''''_f''''''''_r  && \dconPtr_CTf''''''''_f''''''''_d [0])}};
  
  /* demux (Ty MemOut_CTf''''''''_f'''''''',
       Ty Pointer_CTf''''''''_f'''''''') : (memWriteOut_CTf''''''''_f'''''''',MemOut_CTf''''''''_f'''''''') (dconPtr_CTf''''''''_f'''''''',Pointer_CTf''''''''_f'''''''') > [(_35,Pointer_CTf''''''''_f''''''''),
                                                                                                                                                                             (demuxWriteResult_CTf''''''''_f'''''''',Pointer_CTf''''''''_f'''''''')] */
  logic [1:0] \dconPtr_CTf''''''''_f''''''''_onehotd ;
  always_comb
    if ((\memWriteOut_CTf''''''''_f''''''''_d [0] && \dconPtr_CTf''''''''_f''''''''_d [0]))
      unique case (\memWriteOut_CTf''''''''_f''''''''_d [1:1])
        1'd0: \dconPtr_CTf''''''''_f''''''''_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf''''''''_f''''''''_onehotd  = 2'd2;
        default: \dconPtr_CTf''''''''_f''''''''_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf''''''''_f''''''''_onehotd  = 2'd0;
  assign _35_d = {\dconPtr_CTf''''''''_f''''''''_d [16:1],
                  \dconPtr_CTf''''''''_f''''''''_onehotd [0]};
  assign \demuxWriteResult_CTf''''''''_f''''''''_d  = {\dconPtr_CTf''''''''_f''''''''_d [16:1],
                                                       \dconPtr_CTf''''''''_f''''''''_onehotd [1]};
  assign \dconPtr_CTf''''''''_f''''''''_r  = (| (\dconPtr_CTf''''''''_f''''''''_onehotd  & {\demuxWriteResult_CTf''''''''_f''''''''_r ,
                                                                                            _35_r}));
  assign \memWriteOut_CTf''''''''_f''''''''_r  = \dconPtr_CTf''''''''_f''''''''_r ;
  
  /* const (Ty Word16#,Lit 0) : (go__7,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go__8_d[0]) incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go__8_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go__8_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Boo2,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#)] */
  logic [2:0] mergeHP_QTree_Bool_buf_emitted;
  logic [2:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Boo2_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Boo2_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Boo2_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 3'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (wspF_1_1_argbuf,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {wspF_1_1_argbuf_d[16:1],
                                        wspF_1_1_argbuf_d[0]};
  assign wspF_1_1_argbuf_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(readPointer_QTree_BoolwspF_1_1_argbuf,QTree_Bool)] */
  assign readPointer_QTree_BoolwspF_1_1_argbuf_d = {memReadOut_QTree_Bool_d[67:2],
                                                    memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = readPointer_QTree_BoolwspF_1_1_argbuf_r;
  
  /* mergectrl (Ty C18,
           Ty QTree_Bool) : [(lizzieLet11_1_argbuf,QTree_Bool),
                             (lizzieLet14_1_argbuf,QTree_Bool),
                             (lizzieLet19_1_1_argbuf,QTree_Bool),
                             (lizzieLet20_1_1_argbuf,QTree_Bool),
                             (lizzieLet21_1_argbuf,QTree_Bool),
                             (lizzieLet27_1_argbuf,QTree_Bool),
                             (lizzieLet32_1_argbuf,QTree_Bool),
                             (lizzieLet33_1_argbuf,QTree_Bool),
                             (lizzieLet34_1_argbuf,QTree_Bool),
                             (lizzieLet36_1_argbuf,QTree_Bool),
                             (lizzieLet37_1_argbuf,QTree_Bool),
                             (lizzieLet39_1_argbuf,QTree_Bool),
                             (lizzieLet40_1_argbuf,QTree_Bool),
                             (lizzieLet41_1_argbuf,QTree_Bool),
                             (lizzieLet4_1_argbuf,QTree_Bool),
                             (lizzieLet52_1_argbuf,QTree_Bool),
                             (lizzieLet57_1_argbuf,QTree_Bool),
                             (lizzieLet9_1_argbuf,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C18) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [17:0] lizzieLet11_1_argbuf_select_d;
  assign lizzieLet11_1_argbuf_select_d = ((| lizzieLet11_1_argbuf_select_q) ? lizzieLet11_1_argbuf_select_q :
                                          (lizzieLet11_1_argbuf_d[0] ? 18'd1 :
                                           (lizzieLet14_1_argbuf_d[0] ? 18'd2 :
                                            (lizzieLet19_1_1_argbuf_d[0] ? 18'd4 :
                                             (lizzieLet20_1_1_argbuf_d[0] ? 18'd8 :
                                              (lizzieLet21_1_argbuf_d[0] ? 18'd16 :
                                               (lizzieLet27_1_argbuf_d[0] ? 18'd32 :
                                                (lizzieLet32_1_argbuf_d[0] ? 18'd64 :
                                                 (lizzieLet33_1_argbuf_d[0] ? 18'd128 :
                                                  (lizzieLet34_1_argbuf_d[0] ? 18'd256 :
                                                   (lizzieLet36_1_argbuf_d[0] ? 18'd512 :
                                                    (lizzieLet37_1_argbuf_d[0] ? 18'd1024 :
                                                     (lizzieLet39_1_argbuf_d[0] ? 18'd2048 :
                                                      (lizzieLet40_1_argbuf_d[0] ? 18'd4096 :
                                                       (lizzieLet41_1_argbuf_d[0] ? 18'd8192 :
                                                        (lizzieLet4_1_argbuf_d[0] ? 18'd16384 :
                                                         (lizzieLet52_1_argbuf_d[0] ? 18'd32768 :
                                                          (lizzieLet57_1_argbuf_d[0] ? 18'd65536 :
                                                           (lizzieLet9_1_argbuf_d[0] ? 18'd131072 :
                                                            18'd0)))))))))))))))))));
  logic [17:0] lizzieLet11_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_select_q <= 18'd0;
    else
      lizzieLet11_1_argbuf_select_q <= (lizzieLet11_1_argbuf_done ? 18'd0 :
                                        lizzieLet11_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_argbuf_emit_q <= (lizzieLet11_1_argbuf_done ? 2'd0 :
                                      lizzieLet11_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_d;
  assign lizzieLet11_1_argbuf_emit_d = (lizzieLet11_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                        writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                            writeMerge_data_QTree_Bool_r}));
  logic lizzieLet11_1_argbuf_done;
  assign lizzieLet11_1_argbuf_done = (& lizzieLet11_1_argbuf_emit_d);
  assign {lizzieLet9_1_argbuf_r,
          lizzieLet57_1_argbuf_r,
          lizzieLet52_1_argbuf_r,
          lizzieLet4_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet40_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_1_argbuf_r,
          lizzieLet19_1_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (lizzieLet11_1_argbuf_done ? lizzieLet11_1_argbuf_select_d :
                                     18'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet11_1_argbuf_d :
                                         ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                          ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet19_1_1_argbuf_d :
                                           ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet20_1_1_argbuf_d :
                                            ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                             ((lizzieLet11_1_argbuf_select_d[5] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                              ((lizzieLet11_1_argbuf_select_d[6] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                               ((lizzieLet11_1_argbuf_select_d[7] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                ((lizzieLet11_1_argbuf_select_d[8] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                 ((lizzieLet11_1_argbuf_select_d[9] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                  ((lizzieLet11_1_argbuf_select_d[10] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                   ((lizzieLet11_1_argbuf_select_d[11] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                                    ((lizzieLet11_1_argbuf_select_d[12] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                                     ((lizzieLet11_1_argbuf_select_d[13] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                      ((lizzieLet11_1_argbuf_select_d[14] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet4_1_argbuf_d :
                                                       ((lizzieLet11_1_argbuf_select_d[15] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet52_1_argbuf_d :
                                                        ((lizzieLet11_1_argbuf_select_d[16] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet57_1_argbuf_d :
                                                         ((lizzieLet11_1_argbuf_select_d[17] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                          {66'd0, 1'd0}))))))))))))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C1_18_dc(1'd1) :
                                           ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C2_18_dc(1'd1) :
                                            ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C3_18_dc(1'd1) :
                                             ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C4_18_dc(1'd1) :
                                              ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C5_18_dc(1'd1) :
                                               ((lizzieLet11_1_argbuf_select_d[5] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C6_18_dc(1'd1) :
                                                ((lizzieLet11_1_argbuf_select_d[6] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C7_18_dc(1'd1) :
                                                 ((lizzieLet11_1_argbuf_select_d[7] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C8_18_dc(1'd1) :
                                                  ((lizzieLet11_1_argbuf_select_d[8] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C9_18_dc(1'd1) :
                                                   ((lizzieLet11_1_argbuf_select_d[9] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C10_18_dc(1'd1) :
                                                    ((lizzieLet11_1_argbuf_select_d[10] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C11_18_dc(1'd1) :
                                                     ((lizzieLet11_1_argbuf_select_d[11] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C12_18_dc(1'd1) :
                                                      ((lizzieLet11_1_argbuf_select_d[12] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C13_18_dc(1'd1) :
                                                       ((lizzieLet11_1_argbuf_select_d[13] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C14_18_dc(1'd1) :
                                                        ((lizzieLet11_1_argbuf_select_d[14] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C15_18_dc(1'd1) :
                                                         ((lizzieLet11_1_argbuf_select_d[15] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C16_18_dc(1'd1) :
                                                          ((lizzieLet11_1_argbuf_select_d[16] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C17_18_dc(1'd1) :
                                                           ((lizzieLet11_1_argbuf_select_d[17] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C18_18_dc(1'd1) :
                                                            {5'd0, 1'd0}))))))))))))))))));
  
  /* demux (Ty C18,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C18) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet11_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet19_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet20_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet21_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet27_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet32_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet33_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet39_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet40_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet41_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet52_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet57_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet9_1_argbuf,Pointer_QTree_Bool)] */
  logic [17:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[5:1])
        5'd0: demuxWriteResult_QTree_Bool_onehotd = 18'd1;
        5'd1: demuxWriteResult_QTree_Bool_onehotd = 18'd2;
        5'd2: demuxWriteResult_QTree_Bool_onehotd = 18'd4;
        5'd3: demuxWriteResult_QTree_Bool_onehotd = 18'd8;
        5'd4: demuxWriteResult_QTree_Bool_onehotd = 18'd16;
        5'd5: demuxWriteResult_QTree_Bool_onehotd = 18'd32;
        5'd6: demuxWriteResult_QTree_Bool_onehotd = 18'd64;
        5'd7: demuxWriteResult_QTree_Bool_onehotd = 18'd128;
        5'd8: demuxWriteResult_QTree_Bool_onehotd = 18'd256;
        5'd9: demuxWriteResult_QTree_Bool_onehotd = 18'd512;
        5'd10: demuxWriteResult_QTree_Bool_onehotd = 18'd1024;
        5'd11: demuxWriteResult_QTree_Bool_onehotd = 18'd2048;
        5'd12: demuxWriteResult_QTree_Bool_onehotd = 18'd4096;
        5'd13: demuxWriteResult_QTree_Bool_onehotd = 18'd8192;
        5'd14: demuxWriteResult_QTree_Bool_onehotd = 18'd16384;
        5'd15: demuxWriteResult_QTree_Bool_onehotd = 18'd32768;
        5'd16: demuxWriteResult_QTree_Bool_onehotd = 18'd65536;
        5'd17: demuxWriteResult_QTree_Bool_onehotd = 18'd131072;
        default: demuxWriteResult_QTree_Bool_onehotd = 18'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 18'd0;
  assign writeQTree_BoollizzieLet11_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet19_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet20_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet21_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet27_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet32_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[7]};
  assign writeQTree_BoollizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[8]};
  assign writeQTree_BoollizzieLet36_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[9]};
  assign writeQTree_BoollizzieLet37_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[10]};
  assign writeQTree_BoollizzieLet39_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[11]};
  assign writeQTree_BoollizzieLet40_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[12]};
  assign writeQTree_BoollizzieLet41_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[13]};
  assign writeQTree_BoollizzieLet4_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[14]};
  assign writeQTree_BoollizzieLet52_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[15]};
  assign writeQTree_BoollizzieLet57_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[16]};
  assign writeQTree_BoollizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[17]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {writeQTree_BoollizzieLet9_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet57_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet52_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet4_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet41_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet40_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet39_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet37_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet36_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet34_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet33_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet32_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet27_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet21_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet20_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet19_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet14_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet11_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo2,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo2_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo2_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo2_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0]}), forkHP1_QTree_Boo3_d);
  assign {forkHP1_QTree_Boo3_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_34,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _34_d = {dconPtr_QTree_Bool_d[16:1],
                  dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _34_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,Lit 0) : (go__9,Go) > (initHP_CTf_f,Word16#) */
  assign initHP_CTf_f_d = {16'd0, go__9_d[0]};
  assign go__9_r = initHP_CTf_f_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf_f1,Go) > (incrHP_CTf_f,Word16#) */
  assign incrHP_CTf_f_d = {16'd1, incrHP_CTf_f1_d[0]};
  assign incrHP_CTf_f1_r = incrHP_CTf_f_r;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTf_f2,Go)] > (incrHP_mergeCTf_f,Go) */
  logic [1:0] incrHP_mergeCTf_f_selected;
  logic [1:0] incrHP_mergeCTf_f_select;
  always_comb
    begin
      incrHP_mergeCTf_f_selected = 2'd0;
      if ((| incrHP_mergeCTf_f_select))
        incrHP_mergeCTf_f_selected = incrHP_mergeCTf_f_select;
      else
        if (go__10_d[0]) incrHP_mergeCTf_f_selected[0] = 1'd1;
        else if (incrHP_CTf_f2_d[0]) incrHP_mergeCTf_f_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_select <= 2'd0;
    else
      incrHP_mergeCTf_f_select <= (incrHP_mergeCTf_f_r ? 2'd0 :
                                   incrHP_mergeCTf_f_selected);
  always_comb
    if (incrHP_mergeCTf_f_selected[0]) incrHP_mergeCTf_f_d = go__10_d;
    else if (incrHP_mergeCTf_f_selected[1])
      incrHP_mergeCTf_f_d = incrHP_CTf_f2_d;
    else incrHP_mergeCTf_f_d = 1'd0;
  assign {incrHP_CTf_f2_r,
          go__10_r} = (incrHP_mergeCTf_f_r ? incrHP_mergeCTf_f_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_f_buf,Go) > [(incrHP_CTf_f1,Go),
                                             (incrHP_CTf_f2,Go)] */
  logic [1:0] incrHP_mergeCTf_f_buf_emitted;
  logic [1:0] incrHP_mergeCTf_f_buf_done;
  assign incrHP_CTf_f1_d = (incrHP_mergeCTf_f_buf_d[0] && (! incrHP_mergeCTf_f_buf_emitted[0]));
  assign incrHP_CTf_f2_d = (incrHP_mergeCTf_f_buf_d[0] && (! incrHP_mergeCTf_f_buf_emitted[1]));
  assign incrHP_mergeCTf_f_buf_done = (incrHP_mergeCTf_f_buf_emitted | ({incrHP_CTf_f2_d[0],
                                                                         incrHP_CTf_f1_d[0]} & {incrHP_CTf_f2_r,
                                                                                                incrHP_CTf_f1_r}));
  assign incrHP_mergeCTf_f_buf_r = (& incrHP_mergeCTf_f_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_f_buf_emitted <= (incrHP_mergeCTf_f_buf_r ? 2'd0 :
                                        incrHP_mergeCTf_f_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf_f,Word16#) (forkHP1_CTf_f,Word16#) > (addHP_CTf_f,Word16#) */
  assign addHP_CTf_f_d = {(incrHP_CTf_f_d[16:1] + forkHP1_CTf_f_d[16:1]),
                          (incrHP_CTf_f_d[0] && forkHP1_CTf_f_d[0])};
  assign {incrHP_CTf_f_r,
          forkHP1_CTf_f_r} = {2 {(addHP_CTf_f_r && addHP_CTf_f_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf_f,Word16#),
                      (addHP_CTf_f,Word16#)] > (mergeHP_CTf_f,Word16#) */
  logic [1:0] mergeHP_CTf_f_selected;
  logic [1:0] mergeHP_CTf_f_select;
  always_comb
    begin
      mergeHP_CTf_f_selected = 2'd0;
      if ((| mergeHP_CTf_f_select))
        mergeHP_CTf_f_selected = mergeHP_CTf_f_select;
      else
        if (initHP_CTf_f_d[0]) mergeHP_CTf_f_selected[0] = 1'd1;
        else if (addHP_CTf_f_d[0]) mergeHP_CTf_f_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_select <= 2'd0;
    else
      mergeHP_CTf_f_select <= (mergeHP_CTf_f_r ? 2'd0 :
                               mergeHP_CTf_f_selected);
  always_comb
    if (mergeHP_CTf_f_selected[0]) mergeHP_CTf_f_d = initHP_CTf_f_d;
    else if (mergeHP_CTf_f_selected[1])
      mergeHP_CTf_f_d = addHP_CTf_f_d;
    else mergeHP_CTf_f_d = {16'd0, 1'd0};
  assign {addHP_CTf_f_r,
          initHP_CTf_f_r} = (mergeHP_CTf_f_r ? mergeHP_CTf_f_selected :
                             2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf_f,Go) > (incrHP_mergeCTf_f_buf,Go) */
  Go_t incrHP_mergeCTf_f_bufchan_d;
  logic incrHP_mergeCTf_f_bufchan_r;
  assign incrHP_mergeCTf_f_r = ((! incrHP_mergeCTf_f_bufchan_d[0]) || incrHP_mergeCTf_f_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_f_r)
        incrHP_mergeCTf_f_bufchan_d <= incrHP_mergeCTf_f_d;
  Go_t incrHP_mergeCTf_f_bufchan_buf;
  assign incrHP_mergeCTf_f_bufchan_r = (! incrHP_mergeCTf_f_bufchan_buf[0]);
  assign incrHP_mergeCTf_f_buf_d = (incrHP_mergeCTf_f_bufchan_buf[0] ? incrHP_mergeCTf_f_bufchan_buf :
                                    incrHP_mergeCTf_f_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_f_buf_r && incrHP_mergeCTf_f_bufchan_buf[0]))
        incrHP_mergeCTf_f_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_f_buf_r) && (! incrHP_mergeCTf_f_bufchan_buf[0])))
        incrHP_mergeCTf_f_bufchan_buf <= incrHP_mergeCTf_f_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf_f,Word16#) > (mergeHP_CTf_f_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_f_bufchan_d;
  logic mergeHP_CTf_f_bufchan_r;
  assign mergeHP_CTf_f_r = ((! mergeHP_CTf_f_bufchan_d[0]) || mergeHP_CTf_f_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTf_f_r) mergeHP_CTf_f_bufchan_d <= mergeHP_CTf_f_d;
  \Word16#_t  mergeHP_CTf_f_bufchan_buf;
  assign mergeHP_CTf_f_bufchan_r = (! mergeHP_CTf_f_bufchan_buf[0]);
  assign mergeHP_CTf_f_buf_d = (mergeHP_CTf_f_bufchan_buf[0] ? mergeHP_CTf_f_bufchan_buf :
                                mergeHP_CTf_f_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_f_buf_r && mergeHP_CTf_f_bufchan_buf[0]))
        mergeHP_CTf_f_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_f_buf_r) && (! mergeHP_CTf_f_bufchan_buf[0])))
        mergeHP_CTf_f_bufchan_buf <= mergeHP_CTf_f_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_f_buf,Word16#) > [(forkHP1_CTf_f,Word16#),
                                                   (forkHP1_CTf_2,Word16#),
                                                   (forkHP1_CTf_3,Word16#)] */
  logic [2:0] mergeHP_CTf_f_buf_emitted;
  logic [2:0] mergeHP_CTf_f_buf_done;
  assign forkHP1_CTf_f_d = {mergeHP_CTf_f_buf_d[16:1],
                            (mergeHP_CTf_f_buf_d[0] && (! mergeHP_CTf_f_buf_emitted[0]))};
  assign forkHP1_CTf_2_d = {mergeHP_CTf_f_buf_d[16:1],
                            (mergeHP_CTf_f_buf_d[0] && (! mergeHP_CTf_f_buf_emitted[1]))};
  assign forkHP1_CTf_3_d = {mergeHP_CTf_f_buf_d[16:1],
                            (mergeHP_CTf_f_buf_d[0] && (! mergeHP_CTf_f_buf_emitted[2]))};
  assign mergeHP_CTf_f_buf_done = (mergeHP_CTf_f_buf_emitted | ({forkHP1_CTf_3_d[0],
                                                                 forkHP1_CTf_2_d[0],
                                                                 forkHP1_CTf_f_d[0]} & {forkHP1_CTf_3_r,
                                                                                        forkHP1_CTf_2_r,
                                                                                        forkHP1_CTf_f_r}));
  assign mergeHP_CTf_f_buf_r = (& mergeHP_CTf_f_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_f_buf_emitted <= (mergeHP_CTf_f_buf_r ? 3'd0 :
                                    mergeHP_CTf_f_buf_done);
  
  /* mergectrl (Ty C2,Ty MemIn_CTf_f) : [(dconReadIn_CTf_f,MemIn_CTf_f),
                                    (dconWriteIn_CTf_f,MemIn_CTf_f)] > (memMergeChoice_CTf_f,C2) (memMergeIn_CTf_f,MemIn_CTf_f) */
  logic [1:0] dconReadIn_CTf_f_select_d;
  assign dconReadIn_CTf_f_select_d = ((| dconReadIn_CTf_f_select_q) ? dconReadIn_CTf_f_select_q :
                                      (dconReadIn_CTf_f_d[0] ? 2'd1 :
                                       (dconWriteIn_CTf_f_d[0] ? 2'd2 :
                                        2'd0)));
  logic [1:0] dconReadIn_CTf_f_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_select_q <= 2'd0;
    else
      dconReadIn_CTf_f_select_q <= (dconReadIn_CTf_f_done ? 2'd0 :
                                    dconReadIn_CTf_f_select_d);
  logic [1:0] dconReadIn_CTf_f_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_emit_q <= 2'd0;
    else
      dconReadIn_CTf_f_emit_q <= (dconReadIn_CTf_f_done ? 2'd0 :
                                  dconReadIn_CTf_f_emit_d);
  logic [1:0] dconReadIn_CTf_f_emit_d;
  assign dconReadIn_CTf_f_emit_d = (dconReadIn_CTf_f_emit_q | ({memMergeChoice_CTf_f_d[0],
                                                                memMergeIn_CTf_f_d[0]} & {memMergeChoice_CTf_f_r,
                                                                                          memMergeIn_CTf_f_r}));
  logic dconReadIn_CTf_f_done;
  assign dconReadIn_CTf_f_done = (& dconReadIn_CTf_f_emit_d);
  assign {dconWriteIn_CTf_f_r,
          dconReadIn_CTf_f_r} = (dconReadIn_CTf_f_done ? dconReadIn_CTf_f_select_d :
                                 2'd0);
  assign memMergeIn_CTf_f_d = ((dconReadIn_CTf_f_select_d[0] && (! dconReadIn_CTf_f_emit_q[0])) ? dconReadIn_CTf_f_d :
                               ((dconReadIn_CTf_f_select_d[1] && (! dconReadIn_CTf_f_emit_q[0])) ? dconWriteIn_CTf_f_d :
                                {132'd0, 1'd0}));
  assign memMergeChoice_CTf_f_d = ((dconReadIn_CTf_f_select_d[0] && (! dconReadIn_CTf_f_emit_q[1])) ? C1_2_dc(1'd1) :
                                   ((dconReadIn_CTf_f_select_d[1] && (! dconReadIn_CTf_f_emit_q[1])) ? C2_2_dc(1'd1) :
                                    {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf_f,
      Ty MemOut_CTf_f) : (memMergeIn_CTf_f_dbuf,MemIn_CTf_f) > (memOut_CTf_f,MemOut_CTf_f) */
  logic [114:0] memMergeIn_CTf_f_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_f_dbuf_address;
  logic [114:0] memMergeIn_CTf_f_dbuf_din;
  logic [114:0] memOut_CTf_f_q;
  logic memOut_CTf_f_valid;
  logic memMergeIn_CTf_f_dbuf_we;
  logic memOut_CTf_f_we;
  assign memMergeIn_CTf_f_dbuf_din = memMergeIn_CTf_f_dbuf_d[132:18];
  assign memMergeIn_CTf_f_dbuf_address = memMergeIn_CTf_f_dbuf_d[17:2];
  assign memMergeIn_CTf_f_dbuf_we = (memMergeIn_CTf_f_dbuf_d[1:1] && memMergeIn_CTf_f_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_f_we <= 1'd0;
        memOut_CTf_f_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_f_we <= memMergeIn_CTf_f_dbuf_we;
        memOut_CTf_f_valid <= memMergeIn_CTf_f_dbuf_d[0];
        if (memMergeIn_CTf_f_dbuf_we)
          begin
            memMergeIn_CTf_f_dbuf_mem[memMergeIn_CTf_f_dbuf_address] <= memMergeIn_CTf_f_dbuf_din;
            memOut_CTf_f_q <= memMergeIn_CTf_f_dbuf_din;
          end
        else
          memOut_CTf_f_q <= memMergeIn_CTf_f_dbuf_mem[memMergeIn_CTf_f_dbuf_address];
      end
  assign memOut_CTf_f_d = {memOut_CTf_f_q,
                           memOut_CTf_f_we,
                           memOut_CTf_f_valid};
  assign memMergeIn_CTf_f_dbuf_r = ((! memOut_CTf_f_valid) || memOut_CTf_f_r);
  logic [31:0] profiling_MemIn_CTf_f_read;
  logic [31:0] profiling_MemIn_CTf_f_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_f_write <= 0;
        profiling_MemIn_CTf_f_read <= 0;
      end
    else
      if ((memMergeIn_CTf_f_dbuf_we == 1'd1))
        profiling_MemIn_CTf_f_write <= (profiling_MemIn_CTf_f_write + 1);
      else
        if ((memOut_CTf_f_valid == 1'd1))
          profiling_MemIn_CTf_f_read <= (profiling_MemIn_CTf_f_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf_f) : (memMergeChoice_CTf_f,C2) (memOut_CTf_f_dbuf,MemOut_CTf_f) > [(memReadOut_CTf_f,MemOut_CTf_f),
                                                                                        (memWriteOut_CTf_f,MemOut_CTf_f)] */
  logic [1:0] memOut_CTf_f_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_f_d[0] && memOut_CTf_f_dbuf_d[0]))
      unique case (memMergeChoice_CTf_f_d[1:1])
        1'd0: memOut_CTf_f_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_f_dbuf_onehotd = 2'd2;
        default: memOut_CTf_f_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_f_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_f_d = {memOut_CTf_f_dbuf_d[116:1],
                               memOut_CTf_f_dbuf_onehotd[0]};
  assign memWriteOut_CTf_f_d = {memOut_CTf_f_dbuf_d[116:1],
                                memOut_CTf_f_dbuf_onehotd[1]};
  assign memOut_CTf_f_dbuf_r = (| (memOut_CTf_f_dbuf_onehotd & {memWriteOut_CTf_f_r,
                                                                memReadOut_CTf_f_r}));
  assign memMergeChoice_CTf_f_r = memOut_CTf_f_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf_f) : (memMergeIn_CTf_f_rbuf,MemIn_CTf_f) > (memMergeIn_CTf_f_dbuf,MemIn_CTf_f) */
  assign memMergeIn_CTf_f_rbuf_r = ((! memMergeIn_CTf_f_dbuf_d[0]) || memMergeIn_CTf_f_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTf_f_rbuf_r)
        memMergeIn_CTf_f_dbuf_d <= memMergeIn_CTf_f_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf_f) : (memMergeIn_CTf_f,MemIn_CTf_f) > (memMergeIn_CTf_f_rbuf,MemIn_CTf_f) */
  MemIn_CTf_f_t memMergeIn_CTf_f_buf;
  assign memMergeIn_CTf_f_r = (! memMergeIn_CTf_f_buf[0]);
  assign memMergeIn_CTf_f_rbuf_d = (memMergeIn_CTf_f_buf[0] ? memMergeIn_CTf_f_buf :
                                    memMergeIn_CTf_f_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTf_f_rbuf_r && memMergeIn_CTf_f_buf[0]))
        memMergeIn_CTf_f_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTf_f_rbuf_r) && (! memMergeIn_CTf_f_buf[0])))
        memMergeIn_CTf_f_buf <= memMergeIn_CTf_f_d;
  
  /* dbuf (Ty MemOut_CTf_f) : (memOut_CTf_f_rbuf,MemOut_CTf_f) > (memOut_CTf_f_dbuf,MemOut_CTf_f) */
  assign memOut_CTf_f_rbuf_r = ((! memOut_CTf_f_dbuf_d[0]) || memOut_CTf_f_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTf_f_rbuf_r)
        memOut_CTf_f_dbuf_d <= memOut_CTf_f_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf_f) : (memOut_CTf_f,MemOut_CTf_f) > (memOut_CTf_f_rbuf,MemOut_CTf_f) */
  MemOut_CTf_f_t memOut_CTf_f_buf;
  assign memOut_CTf_f_r = (! memOut_CTf_f_buf[0]);
  assign memOut_CTf_f_rbuf_d = (memOut_CTf_f_buf[0] ? memOut_CTf_f_buf :
                                memOut_CTf_f_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTf_f_rbuf_r && memOut_CTf_f_buf[0]))
        memOut_CTf_f_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTf_f_rbuf_r) && (! memOut_CTf_f_buf[0])))
        memOut_CTf_f_buf <= memOut_CTf_f_d;
  
  /* destruct (Ty Pointer_CTf_f,
          Dcon Pointer_CTf_f) : (scfarg_0_2_1_argbuf,Pointer_CTf_f) > [(destructReadIn_CTf_f,Word16#)] */
  assign destructReadIn_CTf_f_d = {scfarg_0_2_1_argbuf_d[16:1],
                                   scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTf_f_r;
  
  /* dcon (Ty MemIn_CTf_f,
      Dcon ReadIn_CTf_f) : [(destructReadIn_CTf_f,Word16#)] > (dconReadIn_CTf_f,MemIn_CTf_f) */
  assign dconReadIn_CTf_f_d = ReadIn_CTf_f_dc((& {destructReadIn_CTf_f_d[0]}), destructReadIn_CTf_f_d);
  assign {destructReadIn_CTf_f_r} = {1 {(dconReadIn_CTf_f_r && dconReadIn_CTf_f_d[0])}};
  
  /* destruct (Ty MemOut_CTf_f,
          Dcon ReadOut_CTf_f) : (memReadOut_CTf_f,MemOut_CTf_f) > [(readPointer_CTf_fscfarg_0_2_1_argbuf,CTf_f)] */
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_d = {memReadOut_CTf_f_d[116:2],
                                                   memReadOut_CTf_f_d[0]};
  assign memReadOut_CTf_f_r = readPointer_CTf_fscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CTf_f) : [(lizzieLet38_1_argbuf,CTf_f),
                              (lizzieLet43_1_argbuf,CTf_f),
                              (lizzieLet54_1_argbuf,CTf_f),
                              (lizzieLet55_1_argbuf,CTf_f),
                              (lizzieLet56_1_argbuf,CTf_f)] > (writeMerge_choice_CTf_f,C5) (writeMerge_data_CTf_f,CTf_f) */
  logic [4:0] lizzieLet38_1_argbuf_select_d;
  assign lizzieLet38_1_argbuf_select_d = ((| lizzieLet38_1_argbuf_select_q) ? lizzieLet38_1_argbuf_select_q :
                                          (lizzieLet38_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet43_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet54_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet55_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet56_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet38_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet38_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet38_1_argbuf_select_q <= (lizzieLet38_1_argbuf_done ? 5'd0 :
                                        lizzieLet38_1_argbuf_select_d);
  logic [1:0] lizzieLet38_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet38_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet38_1_argbuf_emit_q <= (lizzieLet38_1_argbuf_done ? 2'd0 :
                                      lizzieLet38_1_argbuf_emit_d);
  logic [1:0] lizzieLet38_1_argbuf_emit_d;
  assign lizzieLet38_1_argbuf_emit_d = (lizzieLet38_1_argbuf_emit_q | ({writeMerge_choice_CTf_f_d[0],
                                                                        writeMerge_data_CTf_f_d[0]} & {writeMerge_choice_CTf_f_r,
                                                                                                       writeMerge_data_CTf_f_r}));
  logic lizzieLet38_1_argbuf_done;
  assign lizzieLet38_1_argbuf_done = (& lizzieLet38_1_argbuf_emit_d);
  assign {lizzieLet56_1_argbuf_r,
          lizzieLet55_1_argbuf_r,
          lizzieLet54_1_argbuf_r,
          lizzieLet43_1_argbuf_r,
          lizzieLet38_1_argbuf_r} = (lizzieLet38_1_argbuf_done ? lizzieLet38_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_f_d = ((lizzieLet38_1_argbuf_select_d[0] && (! lizzieLet38_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                    ((lizzieLet38_1_argbuf_select_d[1] && (! lizzieLet38_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                     ((lizzieLet38_1_argbuf_select_d[2] && (! lizzieLet38_1_argbuf_emit_q[0])) ? lizzieLet54_1_argbuf_d :
                                      ((lizzieLet38_1_argbuf_select_d[3] && (! lizzieLet38_1_argbuf_emit_q[0])) ? lizzieLet55_1_argbuf_d :
                                       ((lizzieLet38_1_argbuf_select_d[4] && (! lizzieLet38_1_argbuf_emit_q[0])) ? lizzieLet56_1_argbuf_d :
                                        {115'd0, 1'd0})))));
  assign writeMerge_choice_CTf_f_d = ((lizzieLet38_1_argbuf_select_d[0] && (! lizzieLet38_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                      ((lizzieLet38_1_argbuf_select_d[1] && (! lizzieLet38_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                       ((lizzieLet38_1_argbuf_select_d[2] && (! lizzieLet38_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                        ((lizzieLet38_1_argbuf_select_d[3] && (! lizzieLet38_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                         ((lizzieLet38_1_argbuf_select_d[4] && (! lizzieLet38_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                          {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf_f) : (writeMerge_choice_CTf_f,C5) (demuxWriteResult_CTf_f,Pointer_CTf_f) > [(writeCTf_flizzieLet38_1_argbuf,Pointer_CTf_f),
                                                                                                  (writeCTf_flizzieLet43_1_argbuf,Pointer_CTf_f),
                                                                                                  (writeCTf_flizzieLet54_1_argbuf,Pointer_CTf_f),
                                                                                                  (writeCTf_flizzieLet55_1_argbuf,Pointer_CTf_f),
                                                                                                  (writeCTf_flizzieLet56_1_argbuf,Pointer_CTf_f)] */
  logic [4:0] demuxWriteResult_CTf_f_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_f_d[0] && demuxWriteResult_CTf_f_d[0]))
      unique case (writeMerge_choice_CTf_f_d[3:1])
        3'd0: demuxWriteResult_CTf_f_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_f_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_f_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_f_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_f_onehotd = 5'd16;
        default: demuxWriteResult_CTf_f_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_f_onehotd = 5'd0;
  assign writeCTf_flizzieLet38_1_argbuf_d = {demuxWriteResult_CTf_f_d[16:1],
                                             demuxWriteResult_CTf_f_onehotd[0]};
  assign writeCTf_flizzieLet43_1_argbuf_d = {demuxWriteResult_CTf_f_d[16:1],
                                             demuxWriteResult_CTf_f_onehotd[1]};
  assign writeCTf_flizzieLet54_1_argbuf_d = {demuxWriteResult_CTf_f_d[16:1],
                                             demuxWriteResult_CTf_f_onehotd[2]};
  assign writeCTf_flizzieLet55_1_argbuf_d = {demuxWriteResult_CTf_f_d[16:1],
                                             demuxWriteResult_CTf_f_onehotd[3]};
  assign writeCTf_flizzieLet56_1_argbuf_d = {demuxWriteResult_CTf_f_d[16:1],
                                             demuxWriteResult_CTf_f_onehotd[4]};
  assign demuxWriteResult_CTf_f_r = (| (demuxWriteResult_CTf_f_onehotd & {writeCTf_flizzieLet56_1_argbuf_r,
                                                                          writeCTf_flizzieLet55_1_argbuf_r,
                                                                          writeCTf_flizzieLet54_1_argbuf_r,
                                                                          writeCTf_flizzieLet43_1_argbuf_r,
                                                                          writeCTf_flizzieLet38_1_argbuf_r}));
  assign writeMerge_choice_CTf_f_r = demuxWriteResult_CTf_f_r;
  
  /* dcon (Ty MemIn_CTf_f,
      Dcon WriteIn_CTf_f) : [(forkHP1_CTf_2,Word16#),
                             (writeMerge_data_CTf_f,CTf_f)] > (dconWriteIn_CTf_f,MemIn_CTf_f) */
  assign dconWriteIn_CTf_f_d = WriteIn_CTf_f_dc((& {forkHP1_CTf_2_d[0],
                                                    writeMerge_data_CTf_f_d[0]}), forkHP1_CTf_2_d, writeMerge_data_CTf_f_d);
  assign {forkHP1_CTf_2_r,
          writeMerge_data_CTf_f_r} = {2 {(dconWriteIn_CTf_f_r && dconWriteIn_CTf_f_d[0])}};
  
  /* dcon (Ty Pointer_CTf_f,
      Dcon Pointer_CTf_f) : [(forkHP1_CTf_3,Word16#)] > (dconPtr_CTf_f,Pointer_CTf_f) */
  assign dconPtr_CTf_f_d = Pointer_CTf_f_dc((& {forkHP1_CTf_3_d[0]}), forkHP1_CTf_3_d);
  assign {forkHP1_CTf_3_r} = {1 {(dconPtr_CTf_f_r && dconPtr_CTf_f_d[0])}};
  
  /* demux (Ty MemOut_CTf_f,
       Ty Pointer_CTf_f) : (memWriteOut_CTf_f,MemOut_CTf_f) (dconPtr_CTf_f,Pointer_CTf_f) > [(_33,Pointer_CTf_f),
                                                                                             (demuxWriteResult_CTf_f,Pointer_CTf_f)] */
  logic [1:0] dconPtr_CTf_f_onehotd;
  always_comb
    if ((memWriteOut_CTf_f_d[0] && dconPtr_CTf_f_d[0]))
      unique case (memWriteOut_CTf_f_d[1:1])
        1'd0: dconPtr_CTf_f_onehotd = 2'd1;
        1'd1: dconPtr_CTf_f_onehotd = 2'd2;
        default: dconPtr_CTf_f_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_f_onehotd = 2'd0;
  assign _33_d = {dconPtr_CTf_f_d[16:1], dconPtr_CTf_f_onehotd[0]};
  assign demuxWriteResult_CTf_f_d = {dconPtr_CTf_f_d[16:1],
                                     dconPtr_CTf_f_onehotd[1]};
  assign dconPtr_CTf_f_r = (| (dconPtr_CTf_f_onehotd & {demuxWriteResult_CTf_f_r,
                                                        _33_r}));
  assign memWriteOut_CTf_f_r = dconPtr_CTf_f_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Int) : [(m1ae6_1_argbuf,Pointer_QTree_Int),
                                    (m2ae7_1_argbuf,Pointer_QTree_Int),
                                    (q4a8u_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C3) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [2:0] m1ae6_1_argbuf_select_d;
  assign m1ae6_1_argbuf_select_d = ((| m1ae6_1_argbuf_select_q) ? m1ae6_1_argbuf_select_q :
                                    (m1ae6_1_argbuf_d[0] ? 3'd1 :
                                     (m2ae7_1_argbuf_d[0] ? 3'd2 :
                                      (q4a8u_1_argbuf_d[0] ? 3'd4 :
                                       3'd0))));
  logic [2:0] m1ae6_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae6_1_argbuf_select_q <= 3'd0;
    else
      m1ae6_1_argbuf_select_q <= (m1ae6_1_argbuf_done ? 3'd0 :
                                  m1ae6_1_argbuf_select_d);
  logic [1:0] m1ae6_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae6_1_argbuf_emit_q <= 2'd0;
    else
      m1ae6_1_argbuf_emit_q <= (m1ae6_1_argbuf_done ? 2'd0 :
                                m1ae6_1_argbuf_emit_d);
  logic [1:0] m1ae6_1_argbuf_emit_d;
  assign m1ae6_1_argbuf_emit_d = (m1ae6_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1ae6_1_argbuf_done;
  assign m1ae6_1_argbuf_done = (& m1ae6_1_argbuf_emit_d);
  assign {q4a8u_1_argbuf_r,
          m2ae7_1_argbuf_r,
          m1ae6_1_argbuf_r} = (m1ae6_1_argbuf_done ? m1ae6_1_argbuf_select_d :
                               3'd0);
  assign readMerge_data_QTree_Int_d = ((m1ae6_1_argbuf_select_d[0] && (! m1ae6_1_argbuf_emit_q[0])) ? m1ae6_1_argbuf_d :
                                       ((m1ae6_1_argbuf_select_d[1] && (! m1ae6_1_argbuf_emit_q[0])) ? m2ae7_1_argbuf_d :
                                        ((m1ae6_1_argbuf_select_d[2] && (! m1ae6_1_argbuf_emit_q[0])) ? q4a8u_1_argbuf_d :
                                         {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Int_d = ((m1ae6_1_argbuf_select_d[0] && (! m1ae6_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                         ((m1ae6_1_argbuf_select_d[1] && (! m1ae6_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                          ((m1ae6_1_argbuf_select_d[2] && (! m1ae6_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                           {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C3) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1ae6_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm2ae7_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intq4a8u_1_argbuf,QTree_Int)] */
  logic [2:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 3'd4;
        default: destructReadOut_QTree_Int_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 3'd0;
  assign readPointer_QTree_Intm1ae6_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intm2ae7_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intq4a8u_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[2]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intq4a8u_1_argbuf_r,
                                                                                readPointer_QTree_Intm2ae7_1_argbuf_r,
                                                                                readPointer_QTree_Intm1ae6_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (dummy_write_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            dummy_write_QTree_Int_d[0]}), forkHP1_QTree_In3_d, dummy_write_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          dummy_write_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_32,Pointer_QTree_Int),
                                                                                                                 (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _32_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign dummy_write_QTree_Int_sink_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                _32_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (m1aex_0,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2aey_1,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_QTree_Bool) : ($wnnzTupGo___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool) > [($wnnzTupGo___Pointer_QTree_Boolgo_12,Go),
                                                                                                               ($wnnzTupGo___Pointer_QTree_BoolwspF,Pointer_QTree_Bool)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Bool_1_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Bool_1_done ;
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_12_d  = (\$wnnzTupGo___Pointer_QTree_Bool_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Bool_1_emitted [0]));
  assign \$wnnzTupGo___Pointer_QTree_BoolwspF_d  = {\$wnnzTupGo___Pointer_QTree_Bool_1_d [16:1],
                                                    (\$wnnzTupGo___Pointer_QTree_Bool_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Bool_1_emitted [1]))};
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_done  = (\$wnnzTupGo___Pointer_QTree_Bool_1_emitted  | ({\$wnnzTupGo___Pointer_QTree_BoolwspF_d [0],
                                                                                                     \$wnnzTupGo___Pointer_QTree_Boolgo_12_d [0]} & {\$wnnzTupGo___Pointer_QTree_BoolwspF_r ,
                                                                                                                                                     \$wnnzTupGo___Pointer_QTree_Boolgo_12_r }));
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_r  = (& \$wnnzTupGo___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Bool_1_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Bool_1_emitted  <= (\$wnnzTupGo___Pointer_QTree_Bool_1_r  ? 2'd0 :
                                                      \$wnnzTupGo___Pointer_QTree_Bool_1_done );
  
  /* fork (Ty Go) : ($wnnzTupGo___Pointer_QTree_Boolgo_12,Go) > [(go_12_1,Go),
                                                            (go_12_2,Go)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Boolgo_12_done ;
  assign go_12_1_d = (\$wnnzTupGo___Pointer_QTree_Boolgo_12_d [0] && (! \$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted [0]));
  assign go_12_2_d = (\$wnnzTupGo___Pointer_QTree_Boolgo_12_d [0] && (! \$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted [1]));
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_12_done  = (\$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted  | ({go_12_2_d[0],
                                                                                                           go_12_1_d[0]} & {go_12_2_r,
                                                                                                                            go_12_1_r}));
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_12_r  = (& \$wnnzTupGo___Pointer_QTree_Boolgo_12_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Boolgo_12_emitted  <= (\$wnnzTupGo___Pointer_QTree_Boolgo_12_r  ? 2'd0 :
                                                         \$wnnzTupGo___Pointer_QTree_Boolgo_12_done );
  
  /* buf (Ty Pointer_QTree_Bool) : ($wnnzTupGo___Pointer_QTree_BoolwspF,Pointer_QTree_Bool) > (wspF_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d ;
  logic \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_r ;
  assign \$wnnzTupGo___Pointer_QTree_BoolwspF_r  = ((! \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d [0]) || \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wnnzTupGo___Pointer_QTree_BoolwspF_r )
        \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d  <= \$wnnzTupGo___Pointer_QTree_BoolwspF_d ;
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf ;
  assign \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_r  = (! \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf [0]);
  assign wspF_1_argbuf_d = (\$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf [0] ? \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf  :
                            \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((wspF_1_argbuf_r && \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf [0]))
        \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! wspF_1_argbuf_r) && (! \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf [0])))
        \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_buf  <= \$wnnzTupGo___Pointer_QTree_BoolwspF_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_resbuf,Int#)] > (es_1_1I#,Int) */
  assign \es_1_1I#_d  = \I#_dc ((& {\$wnnz_resbuf_d [0]}), \$wnnz_resbuf_d );
  assign {\$wnnz_resbuf_r } = {1 {(\es_1_1I#_r  && \es_1_1I#_d [0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (blae4_1_destruct,Pointer_QTree_Int) > (blae4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t blae4_1_destruct_bufchan_d;
  logic blae4_1_destruct_bufchan_r;
  assign blae4_1_destruct_r = ((! blae4_1_destruct_bufchan_d[0]) || blae4_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) blae4_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (blae4_1_destruct_r)
        blae4_1_destruct_bufchan_d <= blae4_1_destruct_d;
  Pointer_QTree_Int_t blae4_1_destruct_bufchan_buf;
  assign blae4_1_destruct_bufchan_r = (! blae4_1_destruct_bufchan_buf[0]);
  assign blae4_1_1_argbuf_d = (blae4_1_destruct_bufchan_buf[0] ? blae4_1_destruct_bufchan_buf :
                               blae4_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) blae4_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((blae4_1_1_argbuf_r && blae4_1_destruct_bufchan_buf[0]))
        blae4_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! blae4_1_1_argbuf_r) && (! blae4_1_destruct_bufchan_buf[0])))
        blae4_1_destruct_bufchan_buf <= blae4_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (blaec_destruct,Pointer_QTree_Int) > (blaec_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t blaec_destruct_bufchan_d;
  logic blaec_destruct_bufchan_r;
  assign blaec_destruct_r = ((! blaec_destruct_bufchan_d[0]) || blaec_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) blaec_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (blaec_destruct_r) blaec_destruct_bufchan_d <= blaec_destruct_d;
  Pointer_QTree_Int_t blaec_destruct_bufchan_buf;
  assign blaec_destruct_bufchan_r = (! blaec_destruct_bufchan_buf[0]);
  assign blaec_1_argbuf_d = (blaec_destruct_bufchan_buf[0] ? blaec_destruct_bufchan_buf :
                             blaec_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) blaec_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((blaec_1_argbuf_r && blaec_destruct_bufchan_buf[0]))
        blaec_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! blaec_1_argbuf_r) && (! blaec_destruct_bufchan_buf[0])))
        blaec_destruct_bufchan_buf <= blaec_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_4,Go),
                                                                             (boolConvert_1TupGo___Boolbool_3,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_4_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_3_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                              (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_3_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_4_d[0]} & {boolConvert_1TupGo___Boolbool_3_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_4_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool_3,Bool) > [(bool_3_1,Bool),
                                                           (bool_3_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_3_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_3_done;
  assign bool_3_1_d = {boolConvert_1TupGo___Boolbool_3_d[1:1],
                       (boolConvert_1TupGo___Boolbool_3_d[0] && (! boolConvert_1TupGo___Boolbool_3_emitted[0]))};
  assign bool_3_2_d = {boolConvert_1TupGo___Boolbool_3_d[1:1],
                       (boolConvert_1TupGo___Boolbool_3_d[0] && (! boolConvert_1TupGo___Boolbool_3_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_3_done = (boolConvert_1TupGo___Boolbool_3_emitted | ({bool_3_2_d[0],
                                                                                             bool_3_1_d[0]} & {bool_3_2_r,
                                                                                                               bool_3_1_r}));
  assign boolConvert_1TupGo___Boolbool_3_r = (& boolConvert_1TupGo___Boolbool_3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      boolConvert_1TupGo___Boolbool_3_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_3_emitted <= (boolConvert_1TupGo___Boolbool_3_r ? 2'd0 :
                                                  boolConvert_1TupGo___Boolbool_3_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet7_1,MyBool),
                                                    (lizzieLet7_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet7_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet7_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet7_2_d[0],
                                                                       lizzieLet7_1_d[0]} & {lizzieLet7_2_r,
                                                                                             lizzieLet7_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_2TupGo___Bool_1,TupGo___Bool) > [(boolConvert_2TupGo___Boolgo_3,Go),
                                                                             (boolConvert_2TupGo___Boolbool_2,Bool)] */
  logic [1:0] boolConvert_2TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_2TupGo___Bool_1_done;
  assign boolConvert_2TupGo___Boolgo_3_d = (boolConvert_2TupGo___Bool_1_d[0] && (! boolConvert_2TupGo___Bool_1_emitted[0]));
  assign boolConvert_2TupGo___Boolbool_2_d = {boolConvert_2TupGo___Bool_1_d[1:1],
                                              (boolConvert_2TupGo___Bool_1_d[0] && (! boolConvert_2TupGo___Bool_1_emitted[1]))};
  assign boolConvert_2TupGo___Bool_1_done = (boolConvert_2TupGo___Bool_1_emitted | ({boolConvert_2TupGo___Boolbool_2_d[0],
                                                                                     boolConvert_2TupGo___Boolgo_3_d[0]} & {boolConvert_2TupGo___Boolbool_2_r,
                                                                                                                            boolConvert_2TupGo___Boolgo_3_r}));
  assign boolConvert_2TupGo___Bool_1_r = (& boolConvert_2TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_2TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_2TupGo___Bool_1_emitted <= (boolConvert_2TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_2TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_2TupGo___Boolbool_2,Bool) > [(bool_2_1,Bool),
                                                           (bool_2_2,Bool)] */
  logic [1:0] boolConvert_2TupGo___Boolbool_2_emitted;
  logic [1:0] boolConvert_2TupGo___Boolbool_2_done;
  assign bool_2_1_d = {boolConvert_2TupGo___Boolbool_2_d[1:1],
                       (boolConvert_2TupGo___Boolbool_2_d[0] && (! boolConvert_2TupGo___Boolbool_2_emitted[0]))};
  assign bool_2_2_d = {boolConvert_2TupGo___Boolbool_2_d[1:1],
                       (boolConvert_2TupGo___Boolbool_2_d[0] && (! boolConvert_2TupGo___Boolbool_2_emitted[1]))};
  assign boolConvert_2TupGo___Boolbool_2_done = (boolConvert_2TupGo___Boolbool_2_emitted | ({bool_2_2_d[0],
                                                                                             bool_2_1_d[0]} & {bool_2_2_r,
                                                                                                               bool_2_1_r}));
  assign boolConvert_2TupGo___Boolbool_2_r = (& boolConvert_2TupGo___Boolbool_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      boolConvert_2TupGo___Boolbool_2_emitted <= 2'd0;
    else
      boolConvert_2TupGo___Boolbool_2_emitted <= (boolConvert_2TupGo___Boolbool_2_r ? 2'd0 :
                                                  boolConvert_2TupGo___Boolbool_2_done);
  
  /* fork (Ty MyBool) : (boolConvert_2_resbuf,MyBool) > [(lizzieLet17_1,MyBool),
                                                    (lizzieLet17_2,MyBool)] */
  logic [1:0] boolConvert_2_resbuf_emitted;
  logic [1:0] boolConvert_2_resbuf_done;
  assign lizzieLet17_1_d = {boolConvert_2_resbuf_d[1:1],
                            (boolConvert_2_resbuf_d[0] && (! boolConvert_2_resbuf_emitted[0]))};
  assign lizzieLet17_2_d = {boolConvert_2_resbuf_d[1:1],
                            (boolConvert_2_resbuf_d[0] && (! boolConvert_2_resbuf_emitted[1]))};
  assign boolConvert_2_resbuf_done = (boolConvert_2_resbuf_emitted | ({lizzieLet17_2_d[0],
                                                                       lizzieLet17_1_d[0]} & {lizzieLet17_2_r,
                                                                                              lizzieLet17_1_r}));
  assign boolConvert_2_resbuf_r = (& boolConvert_2_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_2_resbuf_emitted <= 2'd0;
    else
      boolConvert_2_resbuf_emitted <= (boolConvert_2_resbuf_r ? 2'd0 :
                                       boolConvert_2_resbuf_done);
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_3TupGo___Bool_1,TupGo___Bool) > [(boolConvert_3TupGo___Boolgo_2,Go),
                                                                             (boolConvert_3TupGo___Boolbool_1,Bool)] */
  logic [1:0] boolConvert_3TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_3TupGo___Bool_1_done;
  assign boolConvert_3TupGo___Boolgo_2_d = (boolConvert_3TupGo___Bool_1_d[0] && (! boolConvert_3TupGo___Bool_1_emitted[0]));
  assign boolConvert_3TupGo___Boolbool_1_d = {boolConvert_3TupGo___Bool_1_d[1:1],
                                              (boolConvert_3TupGo___Bool_1_d[0] && (! boolConvert_3TupGo___Bool_1_emitted[1]))};
  assign boolConvert_3TupGo___Bool_1_done = (boolConvert_3TupGo___Bool_1_emitted | ({boolConvert_3TupGo___Boolbool_1_d[0],
                                                                                     boolConvert_3TupGo___Boolgo_2_d[0]} & {boolConvert_3TupGo___Boolbool_1_r,
                                                                                                                            boolConvert_3TupGo___Boolgo_2_r}));
  assign boolConvert_3TupGo___Bool_1_r = (& boolConvert_3TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_3TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_3TupGo___Bool_1_emitted <= (boolConvert_3TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_3TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_3TupGo___Boolbool_1,Bool) > [(bool_1_1,Bool),
                                                           (bool_1_2,Bool)] */
  logic [1:0] boolConvert_3TupGo___Boolbool_1_emitted;
  logic [1:0] boolConvert_3TupGo___Boolbool_1_done;
  assign bool_1_1_d = {boolConvert_3TupGo___Boolbool_1_d[1:1],
                       (boolConvert_3TupGo___Boolbool_1_d[0] && (! boolConvert_3TupGo___Boolbool_1_emitted[0]))};
  assign bool_1_2_d = {boolConvert_3TupGo___Boolbool_1_d[1:1],
                       (boolConvert_3TupGo___Boolbool_1_d[0] && (! boolConvert_3TupGo___Boolbool_1_emitted[1]))};
  assign boolConvert_3TupGo___Boolbool_1_done = (boolConvert_3TupGo___Boolbool_1_emitted | ({bool_1_2_d[0],
                                                                                             bool_1_1_d[0]} & {bool_1_2_r,
                                                                                                               bool_1_1_r}));
  assign boolConvert_3TupGo___Boolbool_1_r = (& boolConvert_3TupGo___Boolbool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      boolConvert_3TupGo___Boolbool_1_emitted <= 2'd0;
    else
      boolConvert_3TupGo___Boolbool_1_emitted <= (boolConvert_3TupGo___Boolbool_1_r ? 2'd0 :
                                                  boolConvert_3TupGo___Boolbool_1_done);
  
  /* fork (Ty MyBool) : (boolConvert_3_resbuf,MyBool) > [(lizzieLet25_1,MyBool),
                                                    (lizzieLet25_2,MyBool)] */
  logic [1:0] boolConvert_3_resbuf_emitted;
  logic [1:0] boolConvert_3_resbuf_done;
  assign lizzieLet25_1_d = {boolConvert_3_resbuf_d[1:1],
                            (boolConvert_3_resbuf_d[0] && (! boolConvert_3_resbuf_emitted[0]))};
  assign lizzieLet25_2_d = {boolConvert_3_resbuf_d[1:1],
                            (boolConvert_3_resbuf_d[0] && (! boolConvert_3_resbuf_emitted[1]))};
  assign boolConvert_3_resbuf_done = (boolConvert_3_resbuf_emitted | ({lizzieLet25_2_d[0],
                                                                       lizzieLet25_1_d[0]} & {lizzieLet25_2_r,
                                                                                              lizzieLet25_1_r}));
  assign boolConvert_3_resbuf_r = (& boolConvert_3_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_3_resbuf_emitted <= 2'd0;
    else
      boolConvert_3_resbuf_emitted <= (boolConvert_3_resbuf_r ? 2'd0 :
                                       boolConvert_3_resbuf_done);
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_4TupGo___Bool_1,TupGo___Bool) > [(boolConvert_4TupGo___Boolgo_1,Go),
                                                                             (boolConvert_4TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_4TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_4TupGo___Bool_1_done;
  assign boolConvert_4TupGo___Boolgo_1_d = (boolConvert_4TupGo___Bool_1_d[0] && (! boolConvert_4TupGo___Bool_1_emitted[0]));
  assign boolConvert_4TupGo___Boolbool_d = {boolConvert_4TupGo___Bool_1_d[1:1],
                                            (boolConvert_4TupGo___Bool_1_d[0] && (! boolConvert_4TupGo___Bool_1_emitted[1]))};
  assign boolConvert_4TupGo___Bool_1_done = (boolConvert_4TupGo___Bool_1_emitted | ({boolConvert_4TupGo___Boolbool_d[0],
                                                                                     boolConvert_4TupGo___Boolgo_1_d[0]} & {boolConvert_4TupGo___Boolbool_r,
                                                                                                                            boolConvert_4TupGo___Boolgo_1_r}));
  assign boolConvert_4TupGo___Bool_1_r = (& boolConvert_4TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_4TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_4TupGo___Bool_1_emitted <= (boolConvert_4TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_4TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_4TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_4TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_4TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_4TupGo___Boolbool_d[1:1],
                     (boolConvert_4TupGo___Boolbool_d[0] && (! boolConvert_4TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_4TupGo___Boolbool_d[1:1],
                     (boolConvert_4TupGo___Boolbool_d[0] && (! boolConvert_4TupGo___Boolbool_emitted[1]))};
  assign boolConvert_4TupGo___Boolbool_done = (boolConvert_4TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_4TupGo___Boolbool_r = (& boolConvert_4TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_4TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_4TupGo___Boolbool_emitted <= (boolConvert_4TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_4TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_4_resbuf,MyBool) > [(lizzieLet30_1,MyBool),
                                                    (lizzieLet30_2,MyBool)] */
  logic [1:0] boolConvert_4_resbuf_emitted;
  logic [1:0] boolConvert_4_resbuf_done;
  assign lizzieLet30_1_d = {boolConvert_4_resbuf_d[1:1],
                            (boolConvert_4_resbuf_d[0] && (! boolConvert_4_resbuf_emitted[0]))};
  assign lizzieLet30_2_d = {boolConvert_4_resbuf_d[1:1],
                            (boolConvert_4_resbuf_d[0] && (! boolConvert_4_resbuf_emitted[1]))};
  assign boolConvert_4_resbuf_done = (boolConvert_4_resbuf_emitted | ({lizzieLet30_2_d[0],
                                                                       lizzieLet30_1_d[0]} & {lizzieLet30_2_r,
                                                                                              lizzieLet30_1_r}));
  assign boolConvert_4_resbuf_r = (& boolConvert_4_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_4_resbuf_emitted <= 2'd0;
    else
      boolConvert_4_resbuf_emitted <= (boolConvert_4_resbuf_r ? 2'd0 :
                                       boolConvert_4_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_4TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_4TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_4TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_4TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_4TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_4TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_4TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_4TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_4TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_4TupGo___Boolgo_1_r = (| (boolConvert_4TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_4TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_4_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_4_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_4_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_4_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1_1,Bool) (boolConvert_3TupGo___Boolgo_2,Go) > [(bool_1_1False,Go),
                                                                      (bool_1_1True,Go)] */
  logic [1:0] boolConvert_3TupGo___Boolgo_2_onehotd;
  always_comb
    if ((bool_1_1_d[0] && boolConvert_3TupGo___Boolgo_2_d[0]))
      unique case (bool_1_1_d[1:1])
        1'd0: boolConvert_3TupGo___Boolgo_2_onehotd = 2'd1;
        1'd1: boolConvert_3TupGo___Boolgo_2_onehotd = 2'd2;
        default: boolConvert_3TupGo___Boolgo_2_onehotd = 2'd0;
      endcase
    else boolConvert_3TupGo___Boolgo_2_onehotd = 2'd0;
  assign bool_1_1False_d = boolConvert_3TupGo___Boolgo_2_onehotd[0];
  assign bool_1_1True_d = boolConvert_3TupGo___Boolgo_2_onehotd[1];
  assign boolConvert_3TupGo___Boolgo_2_r = (| (boolConvert_3TupGo___Boolgo_2_onehotd & {bool_1_1True_r,
                                                                                        bool_1_1False_r}));
  assign bool_1_1_r = boolConvert_3TupGo___Boolgo_2_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1_1False,Go)] > (bool_1_1False_1MyFalse,MyBool) */
  assign bool_1_1False_1MyFalse_d = MyFalse_dc((& {bool_1_1False_d[0]}), bool_1_1False_d);
  assign {bool_1_1False_r} = {1 {(bool_1_1False_1MyFalse_r && bool_1_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux,MyBool) > (boolConvert_3_resbuf,MyBool) */
  MyBool_t bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d;
  logic bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_r;
  assign bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_r = ((! bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d[0]) || bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                                   1'd0};
    else
      if (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_r)
        bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d <= bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_d;
  MyBool_t bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_r = (! bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_3_resbuf_d = (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                     1'd0};
    else
      if ((boolConvert_3_resbuf_r && bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                       1'd0};
      else if (((! boolConvert_3_resbuf_r) && (! bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_buf <= bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1_1True,Go)] > (bool_1_1True_1MyTrue,MyBool) */
  assign bool_1_1True_1MyTrue_d = MyTrue_dc((& {bool_1_1True_d[0]}), bool_1_1True_d);
  assign {bool_1_1True_r} = {1 {(bool_1_1True_1MyTrue_r && bool_1_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_1_2,Bool) [(bool_1_1False_1MyFalse,MyBool),
                                   (bool_1_1True_1MyTrue,MyBool)] > (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_1_2_d[1:1])
      1'd0:
        {bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_onehot,
         bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux} = {2'd1,
                                                                bool_1_1False_1MyFalse_d};
      1'd1:
        {bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_onehot,
         bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux} = {2'd2,
                                                                bool_1_1True_1MyTrue_d};
      default:
        {bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_onehot,
         bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux} = {2'd0,
                                                                {1'd0, 1'd0}};
    endcase
  assign bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_d = {bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux[1:1],
                                                             (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_mux[0] && bool_1_2_d[0])};
  assign bool_1_2_r = (bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_d[0] && bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_r);
  assign {bool_1_1True_1MyTrue_r,
          bool_1_1False_1MyFalse_r} = (bool_1_2_r ? bool_1_1False_1MyFalsebool_1_1True_1MyTrue_mux_onehot :
                                       2'd0);
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_2_1,Bool) (boolConvert_2TupGo___Boolgo_3,Go) > [(bool_2_1False,Go),
                                                                      (bool_2_1True,Go)] */
  logic [1:0] boolConvert_2TupGo___Boolgo_3_onehotd;
  always_comb
    if ((bool_2_1_d[0] && boolConvert_2TupGo___Boolgo_3_d[0]))
      unique case (bool_2_1_d[1:1])
        1'd0: boolConvert_2TupGo___Boolgo_3_onehotd = 2'd1;
        1'd1: boolConvert_2TupGo___Boolgo_3_onehotd = 2'd2;
        default: boolConvert_2TupGo___Boolgo_3_onehotd = 2'd0;
      endcase
    else boolConvert_2TupGo___Boolgo_3_onehotd = 2'd0;
  assign bool_2_1False_d = boolConvert_2TupGo___Boolgo_3_onehotd[0];
  assign bool_2_1True_d = boolConvert_2TupGo___Boolgo_3_onehotd[1];
  assign boolConvert_2TupGo___Boolgo_3_r = (| (boolConvert_2TupGo___Boolgo_3_onehotd & {bool_2_1True_r,
                                                                                        bool_2_1False_r}));
  assign bool_2_1_r = boolConvert_2TupGo___Boolgo_3_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_2_1False,Go)] > (bool_2_1False_1MyFalse,MyBool) */
  assign bool_2_1False_1MyFalse_d = MyFalse_dc((& {bool_2_1False_d[0]}), bool_2_1False_d);
  assign {bool_2_1False_r} = {1 {(bool_2_1False_1MyFalse_r && bool_2_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux,MyBool) > (boolConvert_2_resbuf,MyBool) */
  MyBool_t bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d;
  logic bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_r;
  assign bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_r = ((! bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d[0]) || bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                                   1'd0};
    else
      if (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_r)
        bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d <= bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_d;
  MyBool_t bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf;
  assign bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_r = (! bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_2_resbuf_d = (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf[0] ? bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf :
                                   bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                     1'd0};
    else
      if ((boolConvert_2_resbuf_r && bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                       1'd0};
      else if (((! boolConvert_2_resbuf_r) && (! bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_buf <= bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_2_1True,Go)] > (bool_2_1True_1MyTrue,MyBool) */
  assign bool_2_1True_1MyTrue_d = MyTrue_dc((& {bool_2_1True_d[0]}), bool_2_1True_d);
  assign {bool_2_1True_r} = {1 {(bool_2_1True_1MyTrue_r && bool_2_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2_2,Bool) [(bool_2_1False_1MyFalse,MyBool),
                                   (bool_2_1True_1MyTrue,MyBool)] > (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux;
  logic [1:0] bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_2_d[1:1])
      1'd0:
        {bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_onehot,
         bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux} = {2'd1,
                                                                bool_2_1False_1MyFalse_d};
      1'd1:
        {bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_onehot,
         bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux} = {2'd2,
                                                                bool_2_1True_1MyTrue_d};
      default:
        {bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_onehot,
         bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux} = {2'd0,
                                                                {1'd0, 1'd0}};
    endcase
  assign bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_d = {bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux[1:1],
                                                             (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_mux[0] && bool_2_2_d[0])};
  assign bool_2_2_r = (bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_d[0] && bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_r);
  assign {bool_2_1True_1MyTrue_r,
          bool_2_1False_1MyFalse_r} = (bool_2_2_r ? bool_2_1False_1MyFalsebool_2_1True_1MyTrue_mux_onehot :
                                       2'd0);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_3_1,Bool) (boolConvert_1TupGo___Boolgo_4,Go) > [(bool_3_1False,Go),
                                                                      (bool_3_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_4_onehotd;
  always_comb
    if ((bool_3_1_d[0] && boolConvert_1TupGo___Boolgo_4_d[0]))
      unique case (bool_3_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_4_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_4_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_4_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_4_onehotd = 2'd0;
  assign bool_3_1False_d = boolConvert_1TupGo___Boolgo_4_onehotd[0];
  assign bool_3_1True_d = boolConvert_1TupGo___Boolgo_4_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_4_r = (| (boolConvert_1TupGo___Boolgo_4_onehotd & {bool_3_1True_r,
                                                                                        bool_3_1False_r}));
  assign bool_3_1_r = boolConvert_1TupGo___Boolgo_4_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_3_1False,Go)] > (bool_3_1False_1MyFalse,MyBool) */
  assign bool_3_1False_1MyFalse_d = MyFalse_dc((& {bool_3_1False_d[0]}), bool_3_1False_d);
  assign {bool_3_1False_r} = {1 {(bool_3_1False_1MyFalse_r && bool_3_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d;
  logic bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_r;
  assign bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_r = ((! bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d[0]) || bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                                   1'd0};
    else
      if (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_r)
        bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d <= bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_d;
  MyBool_t bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf;
  assign bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_r = (! bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf[0] ? bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf :
                                   bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                     1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                       1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_buf <= bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_3_1True,Go)] > (bool_3_1True_1MyTrue,MyBool) */
  assign bool_3_1True_1MyTrue_d = MyTrue_dc((& {bool_3_1True_d[0]}), bool_3_1True_d);
  assign {bool_3_1True_r} = {1 {(bool_3_1True_1MyTrue_r && bool_3_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_3_2,Bool) [(bool_3_1False_1MyFalse,MyBool),
                                   (bool_3_1True_1MyTrue,MyBool)] > (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux;
  logic [1:0] bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_3_2_d[1:1])
      1'd0:
        {bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_onehot,
         bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux} = {2'd1,
                                                                bool_3_1False_1MyFalse_d};
      1'd1:
        {bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_onehot,
         bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux} = {2'd2,
                                                                bool_3_1True_1MyTrue_d};
      default:
        {bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_onehot,
         bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux} = {2'd0,
                                                                {1'd0, 1'd0}};
    endcase
  assign bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_d = {bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux[1:1],
                                                             (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_mux[0] && bool_3_2_d[0])};
  assign bool_3_2_r = (bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_d[0] && bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_r);
  assign {bool_3_1True_1MyTrue_r,
          bool_3_1False_1MyFalse_r} = (bool_3_2_r ? bool_3_1False_1MyFalsebool_3_1True_1MyTrue_mux_onehot :
                                       2'd0);
  
  /* buf (Ty Pointer_QTree_Int) : (brae5_destruct,Pointer_QTree_Int) > (brae5_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t brae5_destruct_bufchan_d;
  logic brae5_destruct_bufchan_r;
  assign brae5_destruct_r = ((! brae5_destruct_bufchan_d[0]) || brae5_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) brae5_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (brae5_destruct_r) brae5_destruct_bufchan_d <= brae5_destruct_d;
  Pointer_QTree_Int_t brae5_destruct_bufchan_buf;
  assign brae5_destruct_bufchan_r = (! brae5_destruct_bufchan_buf[0]);
  assign brae5_1_argbuf_d = (brae5_destruct_bufchan_buf[0] ? brae5_destruct_bufchan_buf :
                             brae5_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) brae5_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((brae5_1_argbuf_r && brae5_destruct_bufchan_buf[0]))
        brae5_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! brae5_1_argbuf_r) && (! brae5_destruct_bufchan_buf[0])))
        brae5_destruct_bufchan_buf <= brae5_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (braed_destruct,Pointer_QTree_Int) > (braed_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t braed_destruct_bufchan_d;
  logic braed_destruct_bufchan_r;
  assign braed_destruct_r = ((! braed_destruct_bufchan_d[0]) || braed_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) braed_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (braed_destruct_r) braed_destruct_bufchan_d <= braed_destruct_d;
  Pointer_QTree_Int_t braed_destruct_bufchan_buf;
  assign braed_destruct_bufchan_r = (! braed_destruct_bufchan_buf[0]);
  assign braed_1_argbuf_d = (braed_destruct_bufchan_buf[0] ? braed_destruct_bufchan_buf :
                             braed_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) braed_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((braed_1_argbuf_r && braed_destruct_bufchan_buf[0]))
        braed_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! braed_1_argbuf_r) && (! braed_destruct_bufchan_buf[0])))
        braed_destruct_bufchan_buf <= braed_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) : (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) > [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13,Go),
                                                                                                                                                                          (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1,Pointer_QTree_Bool),
                                                                                                                                                                          (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] */
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted;
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done;
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d = (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[0]));
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[16:1],
                                                                           (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[1]))};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[32:17],
                                                                         (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[2]))};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done = (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted | ({call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d[0],
                                                                                                                                               call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d[0],
                                                                                                                                               call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d[0]} & {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_r,
                                                                                                                                                                                                                    call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_r,
                                                                                                                                                                                                                    call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_r}));
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r = (& call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted <= 3'd0;
    else
      call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted <= (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r ? 3'd0 :
                                                                           call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_goConst,Go) > (call_$wnnz_initBufi,Go) */
  Go_t call_$wnnz_goConst_buf;
  assign call_$wnnz_goConst_r = (! call_$wnnz_goConst_buf[0]);
  assign call_$wnnz_initBufi_d = (call_$wnnz_goConst_buf[0] ? call_$wnnz_goConst_buf :
                                  call_$wnnz_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_initBufi_r && call_$wnnz_goConst_buf[0]))
        call_$wnnz_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_initBufi_r) && (! call_$wnnz_goConst_buf[0])))
        call_$wnnz_goConst_buf <= call_$wnnz_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_goMux1,Go),
                           (lizzieLet44_3Lcall_$wnnz3_1_argbuf,Go),
                           (lizzieLet44_3Lcall_$wnnz2_1_argbuf,Go),
                           (lizzieLet44_3Lcall_$wnnz1_1_argbuf,Go),
                           (lizzieLet1_3QNode_Bool_1_argbuf,Go)] > (go_13_goMux_choice,C5) (go_13_goMux_data,Go) */
  logic [4:0] call_$wnnz_goMux1_select_d;
  assign call_$wnnz_goMux1_select_d = ((| call_$wnnz_goMux1_select_q) ? call_$wnnz_goMux1_select_q :
                                       (call_$wnnz_goMux1_d[0] ? 5'd1 :
                                        (lizzieLet44_3Lcall_$wnnz3_1_argbuf_d[0] ? 5'd2 :
                                         (lizzieLet44_3Lcall_$wnnz2_1_argbuf_d[0] ? 5'd4 :
                                          (lizzieLet44_3Lcall_$wnnz1_1_argbuf_d[0] ? 5'd8 :
                                           (lizzieLet1_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                            5'd0))))));
  logic [4:0] call_$wnnz_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_goMux1_select_q <= (call_$wnnz_goMux1_done ? 5'd0 :
                                     call_$wnnz_goMux1_select_d);
  logic [1:0] call_$wnnz_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_goMux1_emit_q <= (call_$wnnz_goMux1_done ? 2'd0 :
                                   call_$wnnz_goMux1_emit_d);
  logic [1:0] call_$wnnz_goMux1_emit_d;
  assign call_$wnnz_goMux1_emit_d = (call_$wnnz_goMux1_emit_q | ({go_13_goMux_choice_d[0],
                                                                  go_13_goMux_data_d[0]} & {go_13_goMux_choice_r,
                                                                                            go_13_goMux_data_r}));
  logic call_$wnnz_goMux1_done;
  assign call_$wnnz_goMux1_done = (& call_$wnnz_goMux1_emit_d);
  assign {lizzieLet1_3QNode_Bool_1_argbuf_r,
          lizzieLet44_3Lcall_$wnnz1_1_argbuf_r,
          lizzieLet44_3Lcall_$wnnz2_1_argbuf_r,
          lizzieLet44_3Lcall_$wnnz3_1_argbuf_r,
          call_$wnnz_goMux1_r} = (call_$wnnz_goMux1_done ? call_$wnnz_goMux1_select_d :
                                  5'd0);
  assign go_13_goMux_data_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[0])) ? call_$wnnz_goMux1_d :
                               ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_$wnnz3_1_argbuf_d :
                                ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_$wnnz2_1_argbuf_d :
                                 ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet44_3Lcall_$wnnz1_1_argbuf_d :
                                  ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet1_3QNode_Bool_1_argbuf_d :
                                   1'd0)))));
  assign go_13_goMux_choice_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_initBuf,Go) > [(call_$wnnz_unlockFork1,Go),
                                          (call_$wnnz_unlockFork2,Go),
                                          (call_$wnnz_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_initBuf_emitted;
  logic [2:0] call_$wnnz_initBuf_done;
  assign call_$wnnz_unlockFork1_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[0]));
  assign call_$wnnz_unlockFork2_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[1]));
  assign call_$wnnz_unlockFork3_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[2]));
  assign call_$wnnz_initBuf_done = (call_$wnnz_initBuf_emitted | ({call_$wnnz_unlockFork3_d[0],
                                                                   call_$wnnz_unlockFork2_d[0],
                                                                   call_$wnnz_unlockFork1_d[0]} & {call_$wnnz_unlockFork3_r,
                                                                                                   call_$wnnz_unlockFork2_r,
                                                                                                   call_$wnnz_unlockFork1_r}));
  assign call_$wnnz_initBuf_r = (& call_$wnnz_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_initBuf_emitted <= (call_$wnnz_initBuf_r ? 3'd0 :
                                     call_$wnnz_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_initBufi,Go) > (call_$wnnz_initBuf,Go) */
  assign call_$wnnz_initBufi_r = ((! call_$wnnz_initBuf_d[0]) || call_$wnnz_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_initBufi_r)
        call_$wnnz_initBuf_d <= call_$wnnz_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_unlockFork1,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13,Go)] > (call_$wnnz_goMux1,Go) */
  assign call_$wnnz_goMux1_d = (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d[0]);
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d[0]));
  assign call_$wnnz_unlockFork1_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_13_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_$wnnz_unlockFork2,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1,Pointer_QTree_Bool)] > (call_$wnnz_goMux2,Pointer_QTree_Bool) */
  assign call_$wnnz_goMux2_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d[16:1],
                                (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d[0]));
  assign call_$wnnz_unlockFork2_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwspF_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz) : (call_$wnnz_unlockFork3,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0,Pointer_CT$wnnz)] > (call_$wnnz_goMux3,Pointer_CT$wnnz) */
  assign call_$wnnz_goMux3_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d[16:1],
                                (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d[0]));
  assign call_$wnnz_unlockFork3_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''',
          Dcon TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''') : (call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1,TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''') > [(call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14,Go),
                                                                                                                                                                                                                               (call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u,Pointer_QTree_Int),
                                                                                                                                                                                                                               (call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1,Pointer_CTf''''''''_f'''''''')] */
  logic [2:0] \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted ;
  logic [2:0] \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_done ;
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d  = (\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [0] && (! \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted [0]));
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d  = {\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [16:1],
                                                                                                       (\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [0] && (! \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted [1]))};
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d  = {\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [32:17],
                                                                                                        (\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [0] && (! \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted [2]))};
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_done  = (\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted  | ({\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d [0],
                                                                                                                                                                                                         \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d [0],
                                                                                                                                                                                                         \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d [0]} & {\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_r ,
                                                                                                                                                                                                                                                                                                           \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_r ,
                                                                                                                                                                                                                                                                                                           \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_r }));
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_r  = (& \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted  <= 3'd0;
    else
      \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_emitted  <= (\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_r  ? 3'd0 :
                                                                                                        \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_done );
  
  /* rbuf (Ty Go) : (call_f''''''''_f''''''''_goConst,Go) > (call_f''''''''_f''''''''_initBufi,Go) */
  Go_t \call_f''''''''_f''''''''_goConst_buf ;
  assign \call_f''''''''_f''''''''_goConst_r  = (! \call_f''''''''_f''''''''_goConst_buf [0]);
  assign \call_f''''''''_f''''''''_initBufi_d  = (\call_f''''''''_f''''''''_goConst_buf [0] ? \call_f''''''''_f''''''''_goConst_buf  :
                                                  \call_f''''''''_f''''''''_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_goConst_buf  <= 1'd0;
    else
      if ((\call_f''''''''_f''''''''_initBufi_r  && \call_f''''''''_f''''''''_goConst_buf [0]))
        \call_f''''''''_f''''''''_goConst_buf  <= 1'd0;
      else if (((! \call_f''''''''_f''''''''_initBufi_r ) && (! \call_f''''''''_f''''''''_goConst_buf [0])))
        \call_f''''''''_f''''''''_goConst_buf  <= \call_f''''''''_f''''''''_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f''''''''_f''''''''_goMux1,Go),
                           (lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf,Go),
                           (lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf,Go),
                           (lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf,Go),
                           (lizzieLet3_3QNode_Int_1_argbuf,Go)] > (go_14_goMux_choice,C5) (go_14_goMux_data,Go) */
  logic [4:0] \call_f''''''''_f''''''''_goMux1_select_d ;
  assign \call_f''''''''_f''''''''_goMux1_select_d  = ((| \call_f''''''''_f''''''''_goMux1_select_q ) ? \call_f''''''''_f''''''''_goMux1_select_q  :
                                                       (\call_f''''''''_f''''''''_goMux1_d [0] ? 5'd1 :
                                                        (\lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_d [0] ? 5'd2 :
                                                         (\lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_d [0] ? 5'd4 :
                                                          (\lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_d [0] ? 5'd8 :
                                                           (lizzieLet3_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                            5'd0))))));
  logic [4:0] \call_f''''''''_f''''''''_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_goMux1_select_q  <= 5'd0;
    else
      \call_f''''''''_f''''''''_goMux1_select_q  <= (\call_f''''''''_f''''''''_goMux1_done  ? 5'd0 :
                                                     \call_f''''''''_f''''''''_goMux1_select_d );
  logic [1:0] \call_f''''''''_f''''''''_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_goMux1_emit_q  <= 2'd0;
    else
      \call_f''''''''_f''''''''_goMux1_emit_q  <= (\call_f''''''''_f''''''''_goMux1_done  ? 2'd0 :
                                                   \call_f''''''''_f''''''''_goMux1_emit_d );
  logic [1:0] \call_f''''''''_f''''''''_goMux1_emit_d ;
  assign \call_f''''''''_f''''''''_goMux1_emit_d  = (\call_f''''''''_f''''''''_goMux1_emit_q  | ({go_14_goMux_choice_d[0],
                                                                                                  go_14_goMux_data_d[0]} & {go_14_goMux_choice_r,
                                                                                                                            go_14_goMux_data_r}));
  logic \call_f''''''''_f''''''''_goMux1_done ;
  assign \call_f''''''''_f''''''''_goMux1_done  = (& \call_f''''''''_f''''''''_goMux1_emit_d );
  assign {lizzieLet3_3QNode_Int_1_argbuf_r,
          \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_r ,
          \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_r ,
          \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_r ,
          \call_f''''''''_f''''''''_goMux1_r } = (\call_f''''''''_f''''''''_goMux1_done  ? \call_f''''''''_f''''''''_goMux1_select_d  :
                                                  5'd0);
  assign go_14_goMux_data_d = ((\call_f''''''''_f''''''''_goMux1_select_d [0] && (! \call_f''''''''_f''''''''_goMux1_emit_q [0])) ? \call_f''''''''_f''''''''_goMux1_d  :
                               ((\call_f''''''''_f''''''''_goMux1_select_d [1] && (! \call_f''''''''_f''''''''_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_d  :
                                ((\call_f''''''''_f''''''''_goMux1_select_d [2] && (! \call_f''''''''_f''''''''_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_d  :
                                 ((\call_f''''''''_f''''''''_goMux1_select_d [3] && (! \call_f''''''''_f''''''''_goMux1_emit_q [0])) ? \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_d  :
                                  ((\call_f''''''''_f''''''''_goMux1_select_d [4] && (! \call_f''''''''_f''''''''_goMux1_emit_q [0])) ? lizzieLet3_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_14_goMux_choice_d = ((\call_f''''''''_f''''''''_goMux1_select_d [0] && (! \call_f''''''''_f''''''''_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_f''''''''_f''''''''_goMux1_select_d [1] && (! \call_f''''''''_f''''''''_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_f''''''''_f''''''''_goMux1_select_d [2] && (! \call_f''''''''_f''''''''_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_f''''''''_f''''''''_goMux1_select_d [3] && (! \call_f''''''''_f''''''''_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_f''''''''_f''''''''_goMux1_select_d [4] && (! \call_f''''''''_f''''''''_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f''''''''_f''''''''_initBuf,Go) > [(call_f''''''''_f''''''''_unlockFork1,Go),
                                                        (call_f''''''''_f''''''''_unlockFork2,Go),
                                                        (call_f''''''''_f''''''''_unlockFork3,Go)] */
  logic [2:0] \call_f''''''''_f''''''''_initBuf_emitted ;
  logic [2:0] \call_f''''''''_f''''''''_initBuf_done ;
  assign \call_f''''''''_f''''''''_unlockFork1_d  = (\call_f''''''''_f''''''''_initBuf_d [0] && (! \call_f''''''''_f''''''''_initBuf_emitted [0]));
  assign \call_f''''''''_f''''''''_unlockFork2_d  = (\call_f''''''''_f''''''''_initBuf_d [0] && (! \call_f''''''''_f''''''''_initBuf_emitted [1]));
  assign \call_f''''''''_f''''''''_unlockFork3_d  = (\call_f''''''''_f''''''''_initBuf_d [0] && (! \call_f''''''''_f''''''''_initBuf_emitted [2]));
  assign \call_f''''''''_f''''''''_initBuf_done  = (\call_f''''''''_f''''''''_initBuf_emitted  | ({\call_f''''''''_f''''''''_unlockFork3_d [0],
                                                                                                   \call_f''''''''_f''''''''_unlockFork2_d [0],
                                                                                                   \call_f''''''''_f''''''''_unlockFork1_d [0]} & {\call_f''''''''_f''''''''_unlockFork3_r ,
                                                                                                                                                   \call_f''''''''_f''''''''_unlockFork2_r ,
                                                                                                                                                   \call_f''''''''_f''''''''_unlockFork1_r }));
  assign \call_f''''''''_f''''''''_initBuf_r  = (& \call_f''''''''_f''''''''_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_initBuf_emitted  <= 3'd0;
    else
      \call_f''''''''_f''''''''_initBuf_emitted  <= (\call_f''''''''_f''''''''_initBuf_r  ? 3'd0 :
                                                     \call_f''''''''_f''''''''_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f''''''''_f''''''''_initBufi,Go) > (call_f''''''''_f''''''''_initBuf,Go) */
  assign \call_f''''''''_f''''''''_initBufi_r  = ((! \call_f''''''''_f''''''''_initBuf_d [0]) || \call_f''''''''_f''''''''_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f''''''''_f''''''''_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f''''''''_f''''''''_initBufi_r )
        \call_f''''''''_f''''''''_initBuf_d  <= \call_f''''''''_f''''''''_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f''''''''_f''''''''_unlockFork1,Go) [(call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14,Go)] > (call_f''''''''_f''''''''_goMux1,Go) */
  assign \call_f''''''''_f''''''''_goMux1_d  = (\call_f''''''''_f''''''''_unlockFork1_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d [0]);
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_r  = (\call_f''''''''_f''''''''_goMux1_r  && (\call_f''''''''_f''''''''_unlockFork1_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d [0]));
  assign \call_f''''''''_f''''''''_unlockFork1_r  = (\call_f''''''''_f''''''''_goMux1_r  && (\call_f''''''''_f''''''''_unlockFork1_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''go_14_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f''''''''_f''''''''_unlockFork2,Go) [(call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u,Pointer_QTree_Int)] > (call_f''''''''_f''''''''_goMux2,Pointer_QTree_Int) */
  assign \call_f''''''''_f''''''''_goMux2_d  = {\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d [16:1],
                                                (\call_f''''''''_f''''''''_unlockFork2_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d [0])};
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_r  = (\call_f''''''''_f''''''''_goMux2_r  && (\call_f''''''''_f''''''''_unlockFork2_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d [0]));
  assign \call_f''''''''_f''''''''_unlockFork2_r  = (\call_f''''''''_f''''''''_goMux2_r  && (\call_f''''''''_f''''''''_unlockFork2_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''q4a8u_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf''''''''_f'''''''') : (call_f''''''''_f''''''''_unlockFork3,Go) [(call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1,Pointer_CTf''''''''_f'''''''')] > (call_f''''''''_f''''''''_goMux3,Pointer_CTf''''''''_f'''''''') */
  assign \call_f''''''''_f''''''''_goMux3_d  = {\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d [16:1],
                                                (\call_f''''''''_f''''''''_unlockFork3_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d [0])};
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_r  = (\call_f''''''''_f''''''''_goMux3_r  && (\call_f''''''''_f''''''''_unlockFork3_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d [0]));
  assign \call_f''''''''_f''''''''_unlockFork3_r  = (\call_f''''''''_f''''''''_goMux3_r  && (\call_f''''''''_f''''''''_unlockFork3_d [0] && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''sc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f) : (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f) > [(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15,Go),
                                                                                                                                                                                                                           (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6,Pointer_QTree_Int),
                                                                                                                                                                                                                           (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7,Pointer_QTree_Int),
                                                                                                                                                                                                                           (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2,Pointer_CTf_f)] */
  logic [3:0] call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted;
  logic [3:0] call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_done;
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d = (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[0] && (! call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted[0]));
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[16:1],
                                                                                         (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[0] && (! call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted[1]))};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[32:17],
                                                                                         (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[0] && (! call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted[2]))};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[48:33],
                                                                                          (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[0] && (! call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted[3]))};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_done = (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted | ({call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d[0],
                                                                                                                                                                             call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d[0],
                                                                                                                                                                             call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d[0],
                                                                                                                                                                             call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d[0]} & {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_r,
                                                                                                                                                                                                                                                                 call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_r,
                                                                                                                                                                                                                                                                 call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_r,
                                                                                                                                                                                                                                                                 call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_r}));
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_r = (& call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted <= 4'd0;
    else
      call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_emitted <= (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_r ? 4'd0 :
                                                                                          call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_done);
  
  /* rbuf (Ty Go) : (call_f_f_goConst,Go) > (call_f_f_initBufi,Go) */
  Go_t call_f_f_goConst_buf;
  assign call_f_f_goConst_r = (! call_f_f_goConst_buf[0]);
  assign call_f_f_initBufi_d = (call_f_f_goConst_buf[0] ? call_f_f_goConst_buf :
                                call_f_f_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_goConst_buf <= 1'd0;
    else
      if ((call_f_f_initBufi_r && call_f_f_goConst_buf[0]))
        call_f_f_goConst_buf <= 1'd0;
      else if (((! call_f_f_initBufi_r) && (! call_f_f_goConst_buf[0])))
        call_f_f_goConst_buf <= call_f_f_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_f_goMux1,Go),
                           (lizzieLet53_3Lcall_f_f3_1_argbuf,Go),
                           (lizzieLet53_3Lcall_f_f2_1_argbuf,Go),
                           (lizzieLet53_3Lcall_f_f1_1_argbuf,Go),
                           (lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_15_goMux_choice,C5) (go_15_goMux_data,Go) */
  logic [4:0] call_f_f_goMux1_select_d;
  assign call_f_f_goMux1_select_d = ((| call_f_f_goMux1_select_q) ? call_f_f_goMux1_select_q :
                                     (call_f_f_goMux1_d[0] ? 5'd1 :
                                      (lizzieLet53_3Lcall_f_f3_1_argbuf_d[0] ? 5'd2 :
                                       (lizzieLet53_3Lcall_f_f2_1_argbuf_d[0] ? 5'd4 :
                                        (lizzieLet53_3Lcall_f_f1_1_argbuf_d[0] ? 5'd8 :
                                         (lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                          5'd0))))));
  logic [4:0] call_f_f_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_goMux1_select_q <= 5'd0;
    else
      call_f_f_goMux1_select_q <= (call_f_f_goMux1_done ? 5'd0 :
                                   call_f_f_goMux1_select_d);
  logic [1:0] call_f_f_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_goMux1_emit_q <= 2'd0;
    else
      call_f_f_goMux1_emit_q <= (call_f_f_goMux1_done ? 2'd0 :
                                 call_f_f_goMux1_emit_d);
  logic [1:0] call_f_f_goMux1_emit_d;
  assign call_f_f_goMux1_emit_d = (call_f_f_goMux1_emit_q | ({go_15_goMux_choice_d[0],
                                                              go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                        go_15_goMux_data_r}));
  logic call_f_f_goMux1_done;
  assign call_f_f_goMux1_done = (& call_f_f_goMux1_emit_d);
  assign {lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_r,
          lizzieLet53_3Lcall_f_f1_1_argbuf_r,
          lizzieLet53_3Lcall_f_f2_1_argbuf_r,
          lizzieLet53_3Lcall_f_f3_1_argbuf_r,
          call_f_f_goMux1_r} = (call_f_f_goMux1_done ? call_f_f_goMux1_select_d :
                                5'd0);
  assign go_15_goMux_data_d = ((call_f_f_goMux1_select_d[0] && (! call_f_f_goMux1_emit_q[0])) ? call_f_f_goMux1_d :
                               ((call_f_f_goMux1_select_d[1] && (! call_f_f_goMux1_emit_q[0])) ? lizzieLet53_3Lcall_f_f3_1_argbuf_d :
                                ((call_f_f_goMux1_select_d[2] && (! call_f_f_goMux1_emit_q[0])) ? lizzieLet53_3Lcall_f_f2_1_argbuf_d :
                                 ((call_f_f_goMux1_select_d[3] && (! call_f_f_goMux1_emit_q[0])) ? lizzieLet53_3Lcall_f_f1_1_argbuf_d :
                                  ((call_f_f_goMux1_select_d[4] && (! call_f_f_goMux1_emit_q[0])) ? lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_15_goMux_choice_d = ((call_f_f_goMux1_select_d[0] && (! call_f_f_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_f_f_goMux1_select_d[1] && (! call_f_f_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_f_f_goMux1_select_d[2] && (! call_f_f_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_f_f_goMux1_select_d[3] && (! call_f_f_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_f_f_goMux1_select_d[4] && (! call_f_f_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_f_initBuf,Go) > [(call_f_f_unlockFork1,Go),
                                        (call_f_f_unlockFork2,Go),
                                        (call_f_f_unlockFork3,Go),
                                        (call_f_f_unlockFork4,Go)] */
  logic [3:0] call_f_f_initBuf_emitted;
  logic [3:0] call_f_f_initBuf_done;
  assign call_f_f_unlockFork1_d = (call_f_f_initBuf_d[0] && (! call_f_f_initBuf_emitted[0]));
  assign call_f_f_unlockFork2_d = (call_f_f_initBuf_d[0] && (! call_f_f_initBuf_emitted[1]));
  assign call_f_f_unlockFork3_d = (call_f_f_initBuf_d[0] && (! call_f_f_initBuf_emitted[2]));
  assign call_f_f_unlockFork4_d = (call_f_f_initBuf_d[0] && (! call_f_f_initBuf_emitted[3]));
  assign call_f_f_initBuf_done = (call_f_f_initBuf_emitted | ({call_f_f_unlockFork4_d[0],
                                                               call_f_f_unlockFork3_d[0],
                                                               call_f_f_unlockFork2_d[0],
                                                               call_f_f_unlockFork1_d[0]} & {call_f_f_unlockFork4_r,
                                                                                             call_f_f_unlockFork3_r,
                                                                                             call_f_f_unlockFork2_r,
                                                                                             call_f_f_unlockFork1_r}));
  assign call_f_f_initBuf_r = (& call_f_f_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_initBuf_emitted <= 4'd0;
    else
      call_f_f_initBuf_emitted <= (call_f_f_initBuf_r ? 4'd0 :
                                   call_f_f_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_f_initBufi,Go) > (call_f_f_initBuf,Go) */
  assign call_f_f_initBufi_r = ((! call_f_f_initBuf_d[0]) || call_f_f_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_initBuf_d <= Go_dc(1'd1);
    else
      if (call_f_f_initBufi_r) call_f_f_initBuf_d <= call_f_f_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_f_unlockFork1,Go) [(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15,Go)] > (call_f_f_goMux1,Go) */
  assign call_f_f_goMux1_d = (call_f_f_unlockFork1_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d[0]);
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_r = (call_f_f_goMux1_r && (call_f_f_unlockFork1_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d[0]));
  assign call_f_f_unlockFork1_r = (call_f_f_goMux1_r && (call_f_f_unlockFork1_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fgo_15_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_unlockFork2,Go) [(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6,Pointer_QTree_Int)] > (call_f_f_goMux2,Pointer_QTree_Int) */
  assign call_f_f_goMux2_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d[16:1],
                              (call_f_f_unlockFork2_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d[0])};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_r = (call_f_f_goMux2_r && (call_f_f_unlockFork2_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d[0]));
  assign call_f_f_unlockFork2_r = (call_f_f_goMux2_r && (call_f_f_unlockFork2_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm1ae6_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_unlockFork3,Go) [(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7,Pointer_QTree_Int)] > (call_f_f_goMux3,Pointer_QTree_Int) */
  assign call_f_f_goMux3_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d[16:1],
                              (call_f_f_unlockFork3_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d[0])};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_r = (call_f_f_goMux3_r && (call_f_f_unlockFork3_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d[0]));
  assign call_f_f_unlockFork3_r = (call_f_f_goMux3_r && (call_f_f_unlockFork3_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fm2ae7_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf_f) : (call_f_f_unlockFork4,Go) [(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2,Pointer_CTf_f)] > (call_f_f_goMux4,Pointer_CTf_f) */
  assign call_f_f_goMux4_d = {call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d[16:1],
                              (call_f_f_unlockFork4_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d[0])};
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_r = (call_f_f_goMux4_r && (call_f_f_unlockFork4_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d[0]));
  assign call_f_f_unlockFork4_r = (call_f_f_goMux4_r && (call_f_f_unlockFork4_d[0] && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_fsc_0_2_d[0]));
  
  /* buf (Ty QTree_Bool) : (es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) > (lizzieLet20_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  logic es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_r;
  assign es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_r = ((! es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d[0]) || es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_r)
        es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d <= es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_d;
  QTree_Bool_t es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf;
  assign es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_r = (! es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_1_argbuf_d = (es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0] ? es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf :
                                     es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                             1'd0};
    else
      if ((lizzieLet20_1_1_argbuf_r && es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0]))
        es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                               1'd0};
      else if (((! lizzieLet20_1_1_argbuf_r) && (! es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf[0])))
        es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_buf <= es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_bufchan_d;
  
  /* sink (Ty Int) : (es_1_1I#,Int) > */
  assign {\es_1_1I#_r , \es_1_1I#_dout } = {\es_1_1I#_rout ,
                                            \es_1_1I#_d };
  
  /* buf (Ty Int#) : (es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d;
  logic es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_r;
  assign es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_r = ((! es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d[0]) || es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d <= {32'd0,
                                                              1'd0};
    else
      if (es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_r)
        es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d <= es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_d;
  \Int#_t  es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf;
  assign es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_r = (! es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf[0] ? es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf :
                                 es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]))
        es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                  1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf[0])))
        es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_buf <= es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (es_5_1es_6_1es_7_1es_8_1QNode_Bool,QTree_Bool) > (lizzieLet36_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d;
  logic es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_r;
  assign es_5_1es_6_1es_7_1es_8_1QNode_Bool_r = ((! es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d[0]) || es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_5_1es_6_1es_7_1es_8_1QNode_Bool_r)
        es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d <= es_5_1es_6_1es_7_1es_8_1QNode_Bool_d;
  QTree_Bool_t es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf;
  assign es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_r = (! es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf[0] ? es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf :
                                   es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf[0]))
        es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf[0])))
        es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_buf <= es_5_1es_6_1es_7_1es_8_1QNode_Bool_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_1_1ww2Xqu_1_1_Add32,Int#) (lizzieLet44_4Lcall_$wnnz0,Int#) > (es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32,Int#) */
  assign es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_d = {(es_6_1_1ww2Xqu_1_1_Add32_d[32:1] + lizzieLet44_4Lcall_$wnnz0_d[32:1]),
                                                        (es_6_1_1ww2Xqu_1_1_Add32_d[0] && lizzieLet44_4Lcall_$wnnz0_d[0])};
  assign {es_6_1_1ww2Xqu_1_1_Add32_r,
          lizzieLet44_4Lcall_$wnnz0_r} = {2 {(es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_r && es_4_1_1lizzieLet44_4Lcall_$wnnz0_1_Add32_d[0])}};
  
  /* mergectrl (Ty C4,Ty TupGo) : [(f''''''''1TupGo_1,TupGo),
                              (f''''''''1TupGo2,TupGo),
                              (f''''''''1TupGo3,TupGo),
                              (f''''''''1TupGo4,TupGo)] > (f''''''''1_choice,C4) (f''''''''1_data,TupGo) */
  logic [3:0] \f''''''''1TupGo_1_select_d ;
  assign \f''''''''1TupGo_1_select_d  = ((| \f''''''''1TupGo_1_select_q ) ? \f''''''''1TupGo_1_select_q  :
                                         (\f''''''''1TupGo_1_d [0] ? 4'd1 :
                                          (\f''''''''1TupGo2_d [0] ? 4'd2 :
                                           (\f''''''''1TupGo3_d [0] ? 4'd4 :
                                            (\f''''''''1TupGo4_d [0] ? 4'd8 :
                                             4'd0)))));
  logic [3:0] \f''''''''1TupGo_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1TupGo_1_select_q  <= 4'd0;
    else
      \f''''''''1TupGo_1_select_q  <= (\f''''''''1TupGo_1_done  ? 4'd0 :
                                       \f''''''''1TupGo_1_select_d );
  logic [1:0] \f''''''''1TupGo_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1TupGo_1_emit_q  <= 2'd0;
    else
      \f''''''''1TupGo_1_emit_q  <= (\f''''''''1TupGo_1_done  ? 2'd0 :
                                     \f''''''''1TupGo_1_emit_d );
  logic [1:0] \f''''''''1TupGo_1_emit_d ;
  assign \f''''''''1TupGo_1_emit_d  = (\f''''''''1TupGo_1_emit_q  | ({\f''''''''1_choice_d [0],
                                                                      \f''''''''1_data_d [0]} & {\f''''''''1_choice_r ,
                                                                                                 \f''''''''1_data_r }));
  logic \f''''''''1TupGo_1_done ;
  assign \f''''''''1TupGo_1_done  = (& \f''''''''1TupGo_1_emit_d );
  assign {\f''''''''1TupGo4_r ,
          \f''''''''1TupGo3_r ,
          \f''''''''1TupGo2_r ,
          \f''''''''1TupGo_1_r } = (\f''''''''1TupGo_1_done  ? \f''''''''1TupGo_1_select_d  :
                                    4'd0);
  assign \f''''''''1_data_d  = ((\f''''''''1TupGo_1_select_d [0] && (! \f''''''''1TupGo_1_emit_q [0])) ? \f''''''''1TupGo_1_d  :
                                ((\f''''''''1TupGo_1_select_d [1] && (! \f''''''''1TupGo_1_emit_q [0])) ? \f''''''''1TupGo2_d  :
                                 ((\f''''''''1TupGo_1_select_d [2] && (! \f''''''''1TupGo_1_emit_q [0])) ? \f''''''''1TupGo3_d  :
                                  ((\f''''''''1TupGo_1_select_d [3] && (! \f''''''''1TupGo_1_emit_q [0])) ? \f''''''''1TupGo4_d  :
                                   1'd0))));
  assign \f''''''''1_choice_d  = ((\f''''''''1TupGo_1_select_d [0] && (! \f''''''''1TupGo_1_emit_q [1])) ? C1_4_dc(1'd1) :
                                  ((\f''''''''1TupGo_1_select_d [1] && (! \f''''''''1TupGo_1_emit_q [1])) ? C2_4_dc(1'd1) :
                                   ((\f''''''''1TupGo_1_select_d [2] && (! \f''''''''1TupGo_1_emit_q [1])) ? C3_4_dc(1'd1) :
                                    ((\f''''''''1TupGo_1_select_d [3] && (! \f''''''''1TupGo_1_emit_q [1])) ? C4_4_dc(1'd1) :
                                     {2'd0, 1'd0}))));
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(f''''''''1TupGogo_16,Go)] > (go_16_1MyTrue,MyBool) */
  assign go_16_1MyTrue_d = MyTrue_dc((& {\f''''''''1TupGogo_16_d [0]}), \f''''''''1TupGogo_16_d );
  assign {\f''''''''1TupGogo_16_r } = {1 {(go_16_1MyTrue_r && go_16_1MyTrue_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_1,Pointer_QTree_Bool) > (f''''''''1_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_1_bufchan_d ;
  logic \f''''''''1_1_bufchan_r ;
  assign \f''''''''1_1_r  = ((! \f''''''''1_1_bufchan_d [0]) || \f''''''''1_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_1_r ) \f''''''''1_1_bufchan_d  <= \f''''''''1_1_d ;
  Pointer_QTree_Bool_t \f''''''''1_1_bufchan_buf ;
  assign \f''''''''1_1_bufchan_r  = (! \f''''''''1_1_bufchan_buf [0]);
  assign \f''''''''1_resbuf_d  = (\f''''''''1_1_bufchan_buf [0] ? \f''''''''1_1_bufchan_buf  :
                                  \f''''''''1_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''1_resbuf_r  && \f''''''''1_1_bufchan_buf [0]))
        \f''''''''1_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''1_resbuf_r ) && (! \f''''''''1_1_bufchan_buf [0])))
        \f''''''''1_1_bufchan_buf  <= \f''''''''1_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_2,Pointer_QTree_Bool) > (f''''''''1_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_2_bufchan_d ;
  logic \f''''''''1_2_bufchan_r ;
  assign \f''''''''1_2_r  = ((! \f''''''''1_2_bufchan_d [0]) || \f''''''''1_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_2_r ) \f''''''''1_2_bufchan_d  <= \f''''''''1_2_d ;
  Pointer_QTree_Bool_t \f''''''''1_2_bufchan_buf ;
  assign \f''''''''1_2_bufchan_r  = (! \f''''''''1_2_bufchan_buf [0]);
  assign \f''''''''1_2_argbuf_d  = (\f''''''''1_2_bufchan_buf [0] ? \f''''''''1_2_bufchan_buf  :
                                    \f''''''''1_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''1_2_argbuf_r  && \f''''''''1_2_bufchan_buf [0]))
        \f''''''''1_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''1_2_argbuf_r ) && (! \f''''''''1_2_bufchan_buf [0])))
        \f''''''''1_2_bufchan_buf  <= \f''''''''1_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_2_argbuf,Pointer_QTree_Bool) > (lizzieLet8_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_2_argbuf_bufchan_d ;
  logic \f''''''''1_2_argbuf_bufchan_r ;
  assign \f''''''''1_2_argbuf_r  = ((! \f''''''''1_2_argbuf_bufchan_d [0]) || \f''''''''1_2_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_2_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_2_argbuf_r )
        \f''''''''1_2_argbuf_bufchan_d  <= \f''''''''1_2_argbuf_d ;
  Pointer_QTree_Bool_t \f''''''''1_2_argbuf_bufchan_buf ;
  assign \f''''''''1_2_argbuf_bufchan_r  = (! \f''''''''1_2_argbuf_bufchan_buf [0]);
  assign lizzieLet8_1_argbuf_d = (\f''''''''1_2_argbuf_bufchan_buf [0] ? \f''''''''1_2_argbuf_bufchan_buf  :
                                  \f''''''''1_2_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && \f''''''''1_2_argbuf_bufchan_buf [0]))
        \f''''''''1_2_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! \f''''''''1_2_argbuf_bufchan_buf [0])))
        \f''''''''1_2_argbuf_bufchan_buf  <= \f''''''''1_2_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_3,Pointer_QTree_Bool) > (f''''''''1_3_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_3_bufchan_d ;
  logic \f''''''''1_3_bufchan_r ;
  assign \f''''''''1_3_r  = ((! \f''''''''1_3_bufchan_d [0]) || \f''''''''1_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_3_r ) \f''''''''1_3_bufchan_d  <= \f''''''''1_3_d ;
  Pointer_QTree_Bool_t \f''''''''1_3_bufchan_buf ;
  assign \f''''''''1_3_bufchan_r  = (! \f''''''''1_3_bufchan_buf [0]);
  assign \f''''''''1_3_argbuf_d  = (\f''''''''1_3_bufchan_buf [0] ? \f''''''''1_3_bufchan_buf  :
                                    \f''''''''1_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''1_3_argbuf_r  && \f''''''''1_3_bufchan_buf [0]))
        \f''''''''1_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''1_3_argbuf_r ) && (! \f''''''''1_3_bufchan_buf [0])))
        \f''''''''1_3_bufchan_buf  <= \f''''''''1_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_3_argbuf,Pointer_QTree_Bool) > (lizzieLet26_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_3_argbuf_bufchan_d ;
  logic \f''''''''1_3_argbuf_bufchan_r ;
  assign \f''''''''1_3_argbuf_r  = ((! \f''''''''1_3_argbuf_bufchan_d [0]) || \f''''''''1_3_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_3_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_3_argbuf_r )
        \f''''''''1_3_argbuf_bufchan_d  <= \f''''''''1_3_argbuf_d ;
  Pointer_QTree_Bool_t \f''''''''1_3_argbuf_bufchan_buf ;
  assign \f''''''''1_3_argbuf_bufchan_r  = (! \f''''''''1_3_argbuf_bufchan_buf [0]);
  assign lizzieLet26_1_argbuf_d = (\f''''''''1_3_argbuf_bufchan_buf [0] ? \f''''''''1_3_argbuf_bufchan_buf  :
                                   \f''''''''1_3_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_3_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && \f''''''''1_3_argbuf_bufchan_buf [0]))
        \f''''''''1_3_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! \f''''''''1_3_argbuf_bufchan_buf [0])))
        \f''''''''1_3_argbuf_bufchan_buf  <= \f''''''''1_3_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_4,Pointer_QTree_Bool) > (f''''''''1_4_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_4_bufchan_d ;
  logic \f''''''''1_4_bufchan_r ;
  assign \f''''''''1_4_r  = ((! \f''''''''1_4_bufchan_d [0]) || \f''''''''1_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_4_r ) \f''''''''1_4_bufchan_d  <= \f''''''''1_4_d ;
  Pointer_QTree_Bool_t \f''''''''1_4_bufchan_buf ;
  assign \f''''''''1_4_bufchan_r  = (! \f''''''''1_4_bufchan_buf [0]);
  assign \f''''''''1_4_argbuf_d  = (\f''''''''1_4_bufchan_buf [0] ? \f''''''''1_4_bufchan_buf  :
                                    \f''''''''1_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''1_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''1_4_argbuf_r  && \f''''''''1_4_bufchan_buf [0]))
        \f''''''''1_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''1_4_argbuf_r ) && (! \f''''''''1_4_bufchan_buf [0])))
        \f''''''''1_4_bufchan_buf  <= \f''''''''1_4_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_4_argbuf,Pointer_QTree_Bool) > (lizzieLet31_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_4_argbuf_bufchan_d ;
  logic \f''''''''1_4_argbuf_bufchan_r ;
  assign \f''''''''1_4_argbuf_r  = ((! \f''''''''1_4_argbuf_bufchan_d [0]) || \f''''''''1_4_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_4_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_4_argbuf_r )
        \f''''''''1_4_argbuf_bufchan_d  <= \f''''''''1_4_argbuf_d ;
  Pointer_QTree_Bool_t \f''''''''1_4_argbuf_bufchan_buf ;
  assign \f''''''''1_4_argbuf_bufchan_r  = (! \f''''''''1_4_argbuf_bufchan_buf [0]);
  assign lizzieLet31_1_argbuf_d = (\f''''''''1_4_argbuf_bufchan_buf [0] ? \f''''''''1_4_argbuf_bufchan_buf  :
                                   \f''''''''1_4_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_4_argbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && \f''''''''1_4_argbuf_bufchan_buf [0]))
        \f''''''''1_4_argbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! \f''''''''1_4_argbuf_bufchan_buf [0])))
        \f''''''''1_4_argbuf_bufchan_buf  <= \f''''''''1_4_argbuf_bufchan_d ;
  
  /* demux (Ty C4,
       Ty Pointer_QTree_Bool) : (f''''''''1_choice,C4) (writeQTree_BoollizzieLet41_1_argbuf_rwb,Pointer_QTree_Bool) > [(f''''''''1_1,Pointer_QTree_Bool),
                                                                                                                       (f''''''''1_2,Pointer_QTree_Bool),
                                                                                                                       (f''''''''1_3,Pointer_QTree_Bool),
                                                                                                                       (f''''''''1_4,Pointer_QTree_Bool)] */
  logic [3:0] writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd;
  always_comb
    if ((\f''''''''1_choice_d [0] && writeQTree_BoollizzieLet41_1_argbuf_rwb_d[0]))
      unique case (\f''''''''1_choice_d [2:1])
        2'd0: writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd8;
        default: writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd = 4'd0;
  assign \f''''''''1_1_d  = {writeQTree_BoollizzieLet41_1_argbuf_rwb_d[16:1],
                             writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd[0]};
  assign \f''''''''1_2_d  = {writeQTree_BoollizzieLet41_1_argbuf_rwb_d[16:1],
                             writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd[1]};
  assign \f''''''''1_3_d  = {writeQTree_BoollizzieLet41_1_argbuf_rwb_d[16:1],
                             writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd[2]};
  assign \f''''''''1_4_d  = {writeQTree_BoollizzieLet41_1_argbuf_rwb_d[16:1],
                             writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd[3]};
  assign writeQTree_BoollizzieLet41_1_argbuf_rwb_r = (| (writeQTree_BoollizzieLet41_1_argbuf_rwb_onehotd & {\f''''''''1_4_r ,
                                                                                                            \f''''''''1_3_r ,
                                                                                                            \f''''''''1_2_r ,
                                                                                                            \f''''''''1_1_r }));
  assign \f''''''''1_choice_r  = writeQTree_BoollizzieLet41_1_argbuf_rwb_r;
  
  /* destruct (Ty TupGo,
          Dcon TupGo) : (f''''''''1_data,TupGo) > [(f''''''''1TupGogo_16,Go)] */
  assign \f''''''''1TupGogo_16_d  = \f''''''''1_data_d [0];
  assign \f''''''''1_data_r  = \f''''''''1TupGogo_16_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''1_resbuf,Pointer_QTree_Bool) > (lizzieLet18_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''1_resbuf_bufchan_d ;
  logic \f''''''''1_resbuf_bufchan_r ;
  assign \f''''''''1_resbuf_r  = ((! \f''''''''1_resbuf_bufchan_d [0]) || \f''''''''1_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''1_resbuf_r )
        \f''''''''1_resbuf_bufchan_d  <= \f''''''''1_resbuf_d ;
  Pointer_QTree_Bool_t \f''''''''1_resbuf_bufchan_buf ;
  assign \f''''''''1_resbuf_bufchan_r  = (! \f''''''''1_resbuf_bufchan_buf [0]);
  assign lizzieLet18_2_1_argbuf_d = (\f''''''''1_resbuf_bufchan_buf [0] ? \f''''''''1_resbuf_bufchan_buf  :
                                     \f''''''''1_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''1_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet18_2_1_argbuf_r && \f''''''''1_resbuf_bufchan_buf [0]))
        \f''''''''1_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet18_2_1_argbuf_r) && (! \f''''''''1_resbuf_bufchan_buf [0])))
        \f''''''''1_resbuf_bufchan_buf  <= \f''''''''1_resbuf_bufchan_d ;
  
  /* mergectrl (Ty C8,
           Ty TupGo___Pointer_QTree_Int) : [(f''''''''_f''''''''TupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int2,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int3,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int4,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int5,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int6,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int7,TupGo___Pointer_QTree_Int),
                                            (f''''''''_f''''''''TupGo___Pointer_QTree_Int8,TupGo___Pointer_QTree_Int)] > (f''''''''_f''''''''_choice,C8) (f''''''''_f''''''''_data,TupGo___Pointer_QTree_Int) */
  logic [7:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d  = ((| \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_q ) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_q  :
                                                                      (\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_d [0] ? 8'd1 :
                                                                       (\f''''''''_f''''''''TupGo___Pointer_QTree_Int2_d [0] ? 8'd2 :
                                                                        (\f''''''''_f''''''''TupGo___Pointer_QTree_Int3_d [0] ? 8'd4 :
                                                                         (\f''''''''_f''''''''TupGo___Pointer_QTree_Int4_d [0] ? 8'd8 :
                                                                          (\f''''''''_f''''''''TupGo___Pointer_QTree_Int5_d [0] ? 8'd16 :
                                                                           (\f''''''''_f''''''''TupGo___Pointer_QTree_Int6_d [0] ? 8'd32 :
                                                                            (\f''''''''_f''''''''TupGo___Pointer_QTree_Int7_d [0] ? 8'd64 :
                                                                             (\f''''''''_f''''''''TupGo___Pointer_QTree_Int8_d [0] ? 8'd128 :
                                                                              8'd0)))))))));
  logic [7:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_q  <= 8'd0;
    else
      \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_q  <= (\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_done  ? 8'd0 :
                                                                    \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d );
  logic [1:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q  <= 2'd0;
    else
      \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q  <= (\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_done  ? 2'd0 :
                                                                  \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_d );
  logic [1:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_d ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_d  = (\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q  | ({\f''''''''_f''''''''_choice_d [0],
                                                                                                                                \f''''''''_f''''''''_data_d [0]} & {\f''''''''_f''''''''_choice_r ,
                                                                                                                                                                    \f''''''''_f''''''''_data_r }));
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_done ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_done  = (& \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_d );
  assign {\f''''''''_f''''''''TupGo___Pointer_QTree_Int8_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_r ,
          \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_r } = (\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_done  ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d  :
                                                                 8'd0);
  assign \f''''''''_f''''''''_data_d  = ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [0] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_d  :
                                         ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [1] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_d  :
                                          ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [2] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_d  :
                                           ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [3] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_d  :
                                            ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [4] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_d  :
                                             ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [5] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_d  :
                                              ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [6] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_d  :
                                               ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [7] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [0])) ? \f''''''''_f''''''''TupGo___Pointer_QTree_Int8_d  :
                                                {16'd0, 1'd0}))))))));
  assign \f''''''''_f''''''''_choice_d  = ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [0] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C1_8_dc(1'd1) :
                                           ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [1] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C2_8_dc(1'd1) :
                                            ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [2] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C3_8_dc(1'd1) :
                                             ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [3] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C4_8_dc(1'd1) :
                                              ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [4] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C5_8_dc(1'd1) :
                                               ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [5] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C6_8_dc(1'd1) :
                                                ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [6] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C7_8_dc(1'd1) :
                                                 ((\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_select_d [7] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_emit_q [1])) ? C8_8_dc(1'd1) :
                                                  {3'd0, 1'd0}))))))));
  
  /* fork (Ty Go) : (f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17,Go) > [(go_17_1,Go),
                                                                         (go_17_2,Go)] */
  logic [1:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted ;
  logic [1:0] \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_done ;
  assign go_17_1_d = (\f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_d [0] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted [0]));
  assign go_17_2_d = (\f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_d [0] && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted [1]));
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_done  = (\f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted  | ({go_17_2_d[0],
                                                                                                                                     go_17_1_d[0]} & {go_17_2_r,
                                                                                                                                                      go_17_1_r}));
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_r  = (& \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted  <= 2'd0;
    else
      \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_emitted  <= (\f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_r  ? 2'd0 :
                                                                      \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_done );
  
  /* buf (Ty Pointer_QTree_Int) : (f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1,Pointer_QTree_Int) > (q4a8u_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d ;
  logic \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_r ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_r  = ((! \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d [0]) || \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d  <= {16'd0,
                                                                          1'd0};
    else
      if (\f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_r )
        \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d  <= \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_d ;
  Pointer_QTree_Int_t \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_r  = (! \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf [0]);
  assign q4a8u_1_1_argbuf_d = (\f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf [0] ? \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf  :
                               \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf  <= {16'd0,
                                                                            1'd0};
    else
      if ((q4a8u_1_1_argbuf_r && \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf [0]))
        \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf  <= {16'd0,
                                                                              1'd0};
      else if (((! q4a8u_1_1_argbuf_r) && (! \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf [0])))
        \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_buf  <= \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_1,Pointer_QTree_Bool) > (f''''''''_f''''''''_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_1_bufchan_d ;
  logic \f''''''''_f''''''''_1_bufchan_r ;
  assign \f''''''''_f''''''''_1_r  = ((! \f''''''''_f''''''''_1_bufchan_d [0]) || \f''''''''_f''''''''_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_1_r )
        \f''''''''_f''''''''_1_bufchan_d  <= \f''''''''_f''''''''_1_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_1_bufchan_buf ;
  assign \f''''''''_f''''''''_1_bufchan_r  = (! \f''''''''_f''''''''_1_bufchan_buf [0]);
  assign \f''''''''_f''''''''_resbuf_d  = (\f''''''''_f''''''''_1_bufchan_buf [0] ? \f''''''''_f''''''''_1_bufchan_buf  :
                                           \f''''''''_f''''''''_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_resbuf_r  && \f''''''''_f''''''''_1_bufchan_buf [0]))
        \f''''''''_f''''''''_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_resbuf_r ) && (! \f''''''''_f''''''''_1_bufchan_buf [0])))
        \f''''''''_f''''''''_1_bufchan_buf  <= \f''''''''_f''''''''_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_2,Pointer_QTree_Bool) > (f''''''''_f''''''''_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_2_bufchan_d ;
  logic \f''''''''_f''''''''_2_bufchan_r ;
  assign \f''''''''_f''''''''_2_r  = ((! \f''''''''_f''''''''_2_bufchan_d [0]) || \f''''''''_f''''''''_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_2_r )
        \f''''''''_f''''''''_2_bufchan_d  <= \f''''''''_f''''''''_2_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_2_bufchan_buf ;
  assign \f''''''''_f''''''''_2_bufchan_r  = (! \f''''''''_f''''''''_2_bufchan_buf [0]);
  assign \f''''''''_f''''''''_2_argbuf_d  = (\f''''''''_f''''''''_2_bufchan_buf [0] ? \f''''''''_f''''''''_2_bufchan_buf  :
                                             \f''''''''_f''''''''_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_2_argbuf_r  && \f''''''''_f''''''''_2_bufchan_buf [0]))
        \f''''''''_f''''''''_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_2_argbuf_r ) && (! \f''''''''_f''''''''_2_bufchan_buf [0])))
        \f''''''''_f''''''''_2_bufchan_buf  <= \f''''''''_f''''''''_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_3,Pointer_QTree_Bool) > (f''''''''_f''''''''_3_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_3_bufchan_d ;
  logic \f''''''''_f''''''''_3_bufchan_r ;
  assign \f''''''''_f''''''''_3_r  = ((! \f''''''''_f''''''''_3_bufchan_d [0]) || \f''''''''_f''''''''_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_3_r )
        \f''''''''_f''''''''_3_bufchan_d  <= \f''''''''_f''''''''_3_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_3_bufchan_buf ;
  assign \f''''''''_f''''''''_3_bufchan_r  = (! \f''''''''_f''''''''_3_bufchan_buf [0]);
  assign \f''''''''_f''''''''_3_argbuf_d  = (\f''''''''_f''''''''_3_bufchan_buf [0] ? \f''''''''_f''''''''_3_bufchan_buf  :
                                             \f''''''''_f''''''''_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_3_argbuf_r  && \f''''''''_f''''''''_3_bufchan_buf [0]))
        \f''''''''_f''''''''_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_3_argbuf_r ) && (! \f''''''''_f''''''''_3_bufchan_buf [0])))
        \f''''''''_f''''''''_3_bufchan_buf  <= \f''''''''_f''''''''_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_4,Pointer_QTree_Bool) > (f''''''''_f''''''''_4_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_4_bufchan_d ;
  logic \f''''''''_f''''''''_4_bufchan_r ;
  assign \f''''''''_f''''''''_4_r  = ((! \f''''''''_f''''''''_4_bufchan_d [0]) || \f''''''''_f''''''''_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_4_r )
        \f''''''''_f''''''''_4_bufchan_d  <= \f''''''''_f''''''''_4_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_4_bufchan_buf ;
  assign \f''''''''_f''''''''_4_bufchan_r  = (! \f''''''''_f''''''''_4_bufchan_buf [0]);
  assign \f''''''''_f''''''''_4_argbuf_d  = (\f''''''''_f''''''''_4_bufchan_buf [0] ? \f''''''''_f''''''''_4_bufchan_buf  :
                                             \f''''''''_f''''''''_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_4_argbuf_r  && \f''''''''_f''''''''_4_bufchan_buf [0]))
        \f''''''''_f''''''''_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_4_argbuf_r ) && (! \f''''''''_f''''''''_4_bufchan_buf [0])))
        \f''''''''_f''''''''_4_bufchan_buf  <= \f''''''''_f''''''''_4_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f''''''''_f''''''''_4_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_3_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_2_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_resbuf,Pointer_QTree_Bool)] > (es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool,QTree_Bool) */
  assign es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_d = QNode_Bool_dc((& {\f''''''''_f''''''''_4_argbuf_d [0],
                                                                      \f''''''''_f''''''''_3_argbuf_d [0],
                                                                      \f''''''''_f''''''''_2_argbuf_d [0],
                                                                      \f''''''''_f''''''''_resbuf_d [0]}), \f''''''''_f''''''''_4_argbuf_d , \f''''''''_f''''''''_3_argbuf_d , \f''''''''_f''''''''_2_argbuf_d , \f''''''''_f''''''''_resbuf_d );
  assign {\f''''''''_f''''''''_4_argbuf_r ,
          \f''''''''_f''''''''_3_argbuf_r ,
          \f''''''''_f''''''''_2_argbuf_r ,
          \f''''''''_f''''''''_resbuf_r } = {4 {(es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_r && es_0_1_1es_1_1_1es_2_1es_3_1QNode_Bool_d[0])}};
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_5,Pointer_QTree_Bool) > (f''''''''_f''''''''_5_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_5_bufchan_d ;
  logic \f''''''''_f''''''''_5_bufchan_r ;
  assign \f''''''''_f''''''''_5_r  = ((! \f''''''''_f''''''''_5_bufchan_d [0]) || \f''''''''_f''''''''_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_5_r )
        \f''''''''_f''''''''_5_bufchan_d  <= \f''''''''_f''''''''_5_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_5_bufchan_buf ;
  assign \f''''''''_f''''''''_5_bufchan_r  = (! \f''''''''_f''''''''_5_bufchan_buf [0]);
  assign \f''''''''_f''''''''_5_argbuf_d  = (\f''''''''_f''''''''_5_bufchan_buf [0] ? \f''''''''_f''''''''_5_bufchan_buf  :
                                             \f''''''''_f''''''''_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_5_argbuf_r  && \f''''''''_f''''''''_5_bufchan_buf [0]))
        \f''''''''_f''''''''_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_5_argbuf_r ) && (! \f''''''''_f''''''''_5_bufchan_buf [0])))
        \f''''''''_f''''''''_5_bufchan_buf  <= \f''''''''_f''''''''_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_6,Pointer_QTree_Bool) > (f''''''''_f''''''''_6_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_6_bufchan_d ;
  logic \f''''''''_f''''''''_6_bufchan_r ;
  assign \f''''''''_f''''''''_6_r  = ((! \f''''''''_f''''''''_6_bufchan_d [0]) || \f''''''''_f''''''''_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_6_r )
        \f''''''''_f''''''''_6_bufchan_d  <= \f''''''''_f''''''''_6_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_6_bufchan_buf ;
  assign \f''''''''_f''''''''_6_bufchan_r  = (! \f''''''''_f''''''''_6_bufchan_buf [0]);
  assign \f''''''''_f''''''''_6_argbuf_d  = (\f''''''''_f''''''''_6_bufchan_buf [0] ? \f''''''''_f''''''''_6_bufchan_buf  :
                                             \f''''''''_f''''''''_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_6_argbuf_r  && \f''''''''_f''''''''_6_bufchan_buf [0]))
        \f''''''''_f''''''''_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_6_argbuf_r ) && (! \f''''''''_f''''''''_6_bufchan_buf [0])))
        \f''''''''_f''''''''_6_bufchan_buf  <= \f''''''''_f''''''''_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_7,Pointer_QTree_Bool) > (f''''''''_f''''''''_7_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_7_bufchan_d ;
  logic \f''''''''_f''''''''_7_bufchan_r ;
  assign \f''''''''_f''''''''_7_r  = ((! \f''''''''_f''''''''_7_bufchan_d [0]) || \f''''''''_f''''''''_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_7_r )
        \f''''''''_f''''''''_7_bufchan_d  <= \f''''''''_f''''''''_7_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_7_bufchan_buf ;
  assign \f''''''''_f''''''''_7_bufchan_r  = (! \f''''''''_f''''''''_7_bufchan_buf [0]);
  assign \f''''''''_f''''''''_7_argbuf_d  = (\f''''''''_f''''''''_7_bufchan_buf [0] ? \f''''''''_f''''''''_7_bufchan_buf  :
                                             \f''''''''_f''''''''_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_7_argbuf_r  && \f''''''''_f''''''''_7_bufchan_buf [0]))
        \f''''''''_f''''''''_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_7_argbuf_r ) && (! \f''''''''_f''''''''_7_bufchan_buf [0])))
        \f''''''''_f''''''''_7_bufchan_buf  <= \f''''''''_f''''''''_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_8,Pointer_QTree_Bool) > (f''''''''_f''''''''_8_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \f''''''''_f''''''''_8_bufchan_d ;
  logic \f''''''''_f''''''''_8_bufchan_r ;
  assign \f''''''''_f''''''''_8_r  = ((! \f''''''''_f''''''''_8_bufchan_d [0]) || \f''''''''_f''''''''_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f''''''''_f''''''''_8_r )
        \f''''''''_f''''''''_8_bufchan_d  <= \f''''''''_f''''''''_8_d ;
  Pointer_QTree_Bool_t \f''''''''_f''''''''_8_bufchan_buf ;
  assign \f''''''''_f''''''''_8_bufchan_r  = (! \f''''''''_f''''''''_8_bufchan_buf [0]);
  assign \f''''''''_f''''''''_8_argbuf_d  = (\f''''''''_f''''''''_8_bufchan_buf [0] ? \f''''''''_f''''''''_8_bufchan_buf  :
                                             \f''''''''_f''''''''_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f''''''''_f''''''''_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f''''''''_f''''''''_8_argbuf_r  && \f''''''''_f''''''''_8_bufchan_buf [0]))
        \f''''''''_f''''''''_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f''''''''_f''''''''_8_argbuf_r ) && (! \f''''''''_f''''''''_8_bufchan_buf [0])))
        \f''''''''_f''''''''_8_bufchan_buf  <= \f''''''''_f''''''''_8_bufchan_d ;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(f''''''''_f''''''''_8_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_7_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_6_argbuf,Pointer_QTree_Bool),
                          (f''''''''_f''''''''_5_argbuf,Pointer_QTree_Bool)] > (es_5_1es_6_1es_7_1es_8_1QNode_Bool,QTree_Bool) */
  assign es_5_1es_6_1es_7_1es_8_1QNode_Bool_d = QNode_Bool_dc((& {\f''''''''_f''''''''_8_argbuf_d [0],
                                                                  \f''''''''_f''''''''_7_argbuf_d [0],
                                                                  \f''''''''_f''''''''_6_argbuf_d [0],
                                                                  \f''''''''_f''''''''_5_argbuf_d [0]}), \f''''''''_f''''''''_8_argbuf_d , \f''''''''_f''''''''_7_argbuf_d , \f''''''''_f''''''''_6_argbuf_d , \f''''''''_f''''''''_5_argbuf_d );
  assign {\f''''''''_f''''''''_8_argbuf_r ,
          \f''''''''_f''''''''_7_argbuf_r ,
          \f''''''''_f''''''''_6_argbuf_r ,
          \f''''''''_f''''''''_5_argbuf_r } = {4 {(es_5_1es_6_1es_7_1es_8_1QNode_Bool_r && es_5_1es_6_1es_7_1es_8_1QNode_Bool_d[0])}};
  
  /* demux (Ty C8,
       Ty Pointer_QTree_Bool) : (f''''''''_f''''''''_choice,C8) (lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > [(f''''''''_f''''''''_1,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_2,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_3,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_4,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_5,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_6,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_7,Pointer_QTree_Bool),
                                                                                                                                                   (f''''''''_f''''''''_8,Pointer_QTree_Bool)] */
  logic [7:0] \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f''''''''_f''''''''_choice_d [0] && \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [0]))
      unique case (\f''''''''_f''''''''_choice_d [3:1])
        3'd0:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd1;
        3'd1:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd2;
        3'd2:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd4;
        3'd3:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd8;
        3'd4:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd16;
        3'd5:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd32;
        3'd6:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd64;
        3'd7:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd128;
        default:
          \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd0;
      endcase
    else
      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  = 8'd0;
  assign \f''''''''_f''''''''_1_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f''''''''_f''''''''_2_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f''''''''_f''''''''_3_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f''''''''_f''''''''_4_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f''''''''_f''''''''_5_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f''''''''_f''''''''_6_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f''''''''_f''''''''_7_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f''''''''_f''''''''_8_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [16:1],
                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd [7]};
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_r  = (| (\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_onehotd  & {\f''''''''_f''''''''_8_r ,
                                                                                                                                                      \f''''''''_f''''''''_7_r ,
                                                                                                                                                      \f''''''''_f''''''''_6_r ,
                                                                                                                                                      \f''''''''_f''''''''_5_r ,
                                                                                                                                                      \f''''''''_f''''''''_4_r ,
                                                                                                                                                      \f''''''''_f''''''''_3_r ,
                                                                                                                                                      \f''''''''_f''''''''_2_r ,
                                                                                                                                                      \f''''''''_f''''''''_1_r }));
  assign \f''''''''_f''''''''_choice_r  = \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : (f''''''''_f''''''''_data,TupGo___Pointer_QTree_Int) > [(f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17,Go),
                                                                                                    (f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1,Pointer_QTree_Int)] */
  logic [1:0] \f''''''''_f''''''''_data_emitted ;
  logic [1:0] \f''''''''_f''''''''_data_done ;
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_d  = (\f''''''''_f''''''''_data_d [0] && (! \f''''''''_f''''''''_data_emitted [0]));
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_d  = {\f''''''''_f''''''''_data_d [16:1],
                                                                    (\f''''''''_f''''''''_data_d [0] && (! \f''''''''_f''''''''_data_emitted [1]))};
  assign \f''''''''_f''''''''_data_done  = (\f''''''''_f''''''''_data_emitted  | ({\f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_d [0],
                                                                                   \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_d [0]} & {\f''''''''_f''''''''TupGo___Pointer_QTree_Intq4a8u_1_r ,
                                                                                                                                                \f''''''''_f''''''''TupGo___Pointer_QTree_Intgo_17_r }));
  assign \f''''''''_f''''''''_data_r  = (& \f''''''''_f''''''''_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f''''''''_f''''''''_data_emitted  <= 2'd0;
    else
      \f''''''''_f''''''''_data_emitted  <= (\f''''''''_f''''''''_data_r  ? 2'd0 :
                                             \f''''''''_f''''''''_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) > [(f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18,Go),
                                                                                                                                                                      (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1,Pointer_QTree_Int),
                                                                                                                                                                      (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1,Pointer_QTree_Int)] */
  logic [2:0] f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted;
  logic [2:0] f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done;
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_d = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[0]));
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_d = {f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[16:1],
                                                                      (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[1]))};
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_d = {f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[32:17],
                                                                      (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0] && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted[2]))};
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted | ({f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_d[0],
                                                                                                                                   f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_d[0],
                                                                                                                                   f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_d[0]} & {f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_r,
                                                                                                                                                                                                  f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_r,
                                                                                                                                                                                                  f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_r}));
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r = (& f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= 3'd0;
    else
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted <= (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r ? 3'd0 :
                                                                     f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done);
  
  /* fork (Ty Go) : (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18,Go) > [(go_18_1,Go),
                                                                             (go_18_2,Go)] */
  logic [1:0] f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted;
  logic [1:0] f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_done;
  assign go_18_1_d = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_d[0] && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted[0]));
  assign go_18_2_d = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_d[0] && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted[1]));
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_done = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted | ({go_18_2_d[0],
                                                                                                                                         go_18_1_d[0]} & {go_18_2_r,
                                                                                                                                                          go_18_1_r}));
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_r = (& f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted <= 2'd0;
    else
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_emitted <= (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_r ? 2'd0 :
                                                                        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_18_done);
  
  /* buf (Ty Pointer_QTree_Int) : (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1,Pointer_QTree_Int) > (m1ae6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_r;
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_r = ((! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d[0]) || f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_r)
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d <= f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_d;
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf;
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_r = (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf[0]);
  assign m1ae6_1_1_argbuf_d = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf[0] ? f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf :
                               f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((m1ae6_1_1_argbuf_r && f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf[0]))
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! m1ae6_1_1_argbuf_r) && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf[0])))
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_buf <= f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm1ae6_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1,Pointer_QTree_Int) > (m2ae7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d;
  logic f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_r;
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_r = ((! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d[0]) || f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_r)
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d <= f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_d;
  Pointer_QTree_Int_t f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf;
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_r = (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf[0]);
  assign m2ae7_1_1_argbuf_d = (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf[0] ? f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf :
                               f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((m2ae7_1_1_argbuf_r && f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf[0]))
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! m2ae7_1_1_argbuf_r) && (! f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf[0])))
        f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_buf <= f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Intm2ae7_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (f_f_resbuf,Pointer_QTree_Bool) > (es_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t f_f_resbuf_bufchan_d;
  logic f_f_resbuf_bufchan_r;
  assign f_f_resbuf_r = ((! f_f_resbuf_bufchan_d[0]) || f_f_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_resbuf_bufchan_d <= {16'd0, 1'd0};
    else if (f_f_resbuf_r) f_f_resbuf_bufchan_d <= f_f_resbuf_d;
  Pointer_QTree_Bool_t f_f_resbuf_bufchan_buf;
  assign f_f_resbuf_bufchan_r = (! f_f_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (f_f_resbuf_bufchan_buf[0] ? f_f_resbuf_bufchan_buf :
                            f_f_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && f_f_resbuf_bufchan_buf[0]))
        f_f_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! f_f_resbuf_bufchan_buf[0])))
        f_f_resbuf_bufchan_buf <= f_f_resbuf_bufchan_d;
  
  /* buf (Ty Go) : (go_1,Go) > (go_1_argbuf,Go) */
  Go_t go_1_bufchan_d;
  logic go_1_bufchan_r;
  assign go_1_r = ((! go_1_bufchan_d[0]) || go_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1_bufchan_d <= 1'd0;
    else if (go_1_r) go_1_bufchan_d <= go_1_d;
  Go_t go_1_bufchan_buf;
  assign go_1_bufchan_r = (! go_1_bufchan_buf[0]);
  assign go_1_argbuf_d = (go_1_bufchan_buf[0] ? go_1_bufchan_buf :
                          go_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1_bufchan_buf <= 1'd0;
    else
      if ((go_1_argbuf_r && go_1_bufchan_buf[0]))
        go_1_bufchan_buf <= 1'd0;
      else if (((! go_1_argbuf_r) && (! go_1_bufchan_buf[0])))
        go_1_bufchan_buf <= go_1_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon L$wnnzsbos) : [(go_12_1,Go)] > (go_12_1L$wnnzsbos,CT$wnnz) */
  assign go_12_1L$wnnzsbos_d = L$wnnzsbos_dc((& {go_12_1_d[0]}), go_12_1_d);
  assign {go_12_1_r} = {1 {(go_12_1L$wnnzsbos_r && go_12_1L$wnnzsbos_d[0])}};
  
  /* buf (Ty CT$wnnz) : (go_12_1L$wnnzsbos,CT$wnnz) > (lizzieLet0_1_argbuf,CT$wnnz) */
  CT$wnnz_t go_12_1L$wnnzsbos_bufchan_d;
  logic go_12_1L$wnnzsbos_bufchan_r;
  assign go_12_1L$wnnzsbos_r = ((! go_12_1L$wnnzsbos_bufchan_d[0]) || go_12_1L$wnnzsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_1L$wnnzsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_12_1L$wnnzsbos_r)
        go_12_1L$wnnzsbos_bufchan_d <= go_12_1L$wnnzsbos_d;
  CT$wnnz_t go_12_1L$wnnzsbos_bufchan_buf;
  assign go_12_1L$wnnzsbos_bufchan_r = (! go_12_1L$wnnzsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_12_1L$wnnzsbos_bufchan_buf[0] ? go_12_1L$wnnzsbos_bufchan_buf :
                                  go_12_1L$wnnzsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_12_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_12_1L$wnnzsbos_bufchan_buf[0]))
        go_12_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_12_1L$wnnzsbos_bufchan_buf[0])))
        go_12_1L$wnnzsbos_bufchan_buf <= go_12_1L$wnnzsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_12_2,Go) > (go_12_2_argbuf,Go) */
  Go_t go_12_2_bufchan_d;
  logic go_12_2_bufchan_r;
  assign go_12_2_r = ((! go_12_2_bufchan_d[0]) || go_12_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_d <= 1'd0;
    else if (go_12_2_r) go_12_2_bufchan_d <= go_12_2_d;
  Go_t go_12_2_bufchan_buf;
  assign go_12_2_bufchan_r = (! go_12_2_bufchan_buf[0]);
  assign go_12_2_argbuf_d = (go_12_2_bufchan_buf[0] ? go_12_2_bufchan_buf :
                             go_12_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_buf <= 1'd0;
    else
      if ((go_12_2_argbuf_r && go_12_2_bufchan_buf[0]))
        go_12_2_bufchan_buf <= 1'd0;
      else if (((! go_12_2_argbuf_r) && (! go_12_2_bufchan_buf[0])))
        go_12_2_bufchan_buf <= go_12_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) : [(go_12_2_argbuf,Go),
                                                            (wspF_1_argbuf,Pointer_QTree_Bool),
                                                            (lizzieLet20_1_argbuf,Pointer_CT$wnnz)] > (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) */
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d = TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_dc((& {go_12_2_argbuf_d[0],
                                                                                                                          wspF_1_argbuf_d[0],
                                                                                                                          lizzieLet20_1_argbuf_d[0]}), go_12_2_argbuf_d, wspF_1_argbuf_d, lizzieLet20_1_argbuf_d);
  assign {go_12_2_argbuf_r,
          wspF_1_argbuf_r,
          lizzieLet20_1_argbuf_r} = {3 {(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0])}};
  
  /* fork (Ty C5) : (go_13_goMux_choice,C5) > [(go_13_goMux_choice_1,C5),
                                          (go_13_goMux_choice_2,C5)] */
  logic [1:0] go_13_goMux_choice_emitted;
  logic [1:0] go_13_goMux_choice_done;
  assign go_13_goMux_choice_1_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[0]))};
  assign go_13_goMux_choice_2_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[1]))};
  assign go_13_goMux_choice_done = (go_13_goMux_choice_emitted | ({go_13_goMux_choice_2_d[0],
                                                                   go_13_goMux_choice_1_d[0]} & {go_13_goMux_choice_2_r,
                                                                                                 go_13_goMux_choice_1_r}));
  assign go_13_goMux_choice_r = (& go_13_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_goMux_choice_emitted <= 2'd0;
    else
      go_13_goMux_choice_emitted <= (go_13_goMux_choice_r ? 2'd0 :
                                     go_13_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_13_goMux_choice_1,C5) [(call_$wnnz_goMux2,Pointer_QTree_Bool),
                                                         (q2a85_1_1_argbuf,Pointer_QTree_Bool),
                                                         (q3a86_2_1_argbuf,Pointer_QTree_Bool),
                                                         (q4a87_3_1_argbuf,Pointer_QTree_Bool),
                                                         (q1a84_1_argbuf,Pointer_QTree_Bool)] > (wspF_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] wspF_1_goMux_mux_mux;
  logic [4:0] wspF_1_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_1_d[3:1])
      3'd0:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_goMux2_d};
      3'd1:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd2,
                                                           q2a85_1_1_argbuf_d};
      3'd2:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd4,
                                                           q3a86_2_1_argbuf_d};
      3'd3:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd8,
                                                           q4a87_3_1_argbuf_d};
      3'd4:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd16,
                                                           q1a84_1_argbuf_d};
      default:
        {wspF_1_goMux_mux_onehot, wspF_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wspF_1_goMux_mux_d = {wspF_1_goMux_mux_mux[16:1],
                               (wspF_1_goMux_mux_mux[0] && go_13_goMux_choice_1_d[0])};
  assign go_13_goMux_choice_1_r = (wspF_1_goMux_mux_d[0] && wspF_1_goMux_mux_r);
  assign {q1a84_1_argbuf_r,
          q4a87_3_1_argbuf_r,
          q3a86_2_1_argbuf_r,
          q2a85_1_1_argbuf_r,
          call_$wnnz_goMux2_r} = (go_13_goMux_choice_1_r ? wspF_1_goMux_mux_onehot :
                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz) : (go_13_goMux_choice_2,C5) [(call_$wnnz_goMux3,Pointer_CT$wnnz),
                                                      (sca2_1_argbuf,Pointer_CT$wnnz),
                                                      (sca1_1_argbuf,Pointer_CT$wnnz),
                                                      (sca0_1_argbuf,Pointer_CT$wnnz),
                                                      (sca3_1_argbuf,Pointer_CT$wnnz)] > (sc_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_13_goMux_choice_2_d[0])};
  assign go_13_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_goMux3_r} = (go_13_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                  5'd0);
  
  /* fork (Ty C5) : (go_14_goMux_choice,C5) > [(go_14_goMux_choice_1,C5),
                                          (go_14_goMux_choice_2,C5)] */
  logic [1:0] go_14_goMux_choice_emitted;
  logic [1:0] go_14_goMux_choice_done;
  assign go_14_goMux_choice_1_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[0]))};
  assign go_14_goMux_choice_2_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[1]))};
  assign go_14_goMux_choice_done = (go_14_goMux_choice_emitted | ({go_14_goMux_choice_2_d[0],
                                                                   go_14_goMux_choice_1_d[0]} & {go_14_goMux_choice_2_r,
                                                                                                 go_14_goMux_choice_1_r}));
  assign go_14_goMux_choice_r = (& go_14_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_goMux_choice_emitted <= 2'd0;
    else
      go_14_goMux_choice_emitted <= (go_14_goMux_choice_r ? 2'd0 :
                                     go_14_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_14_goMux_choice_1,C5) [(call_f''''''''_f''''''''_goMux2,Pointer_QTree_Int),
                                                        (blae4_1_1_argbuf,Pointer_QTree_Int),
                                                        (trae3_2_1_argbuf,Pointer_QTree_Int),
                                                        (tlae2_3_1_argbuf,Pointer_QTree_Int),
                                                        (brae5_1_argbuf,Pointer_QTree_Int)] > (q4a8u_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] q4a8u_goMux_mux_mux;
  logic [4:0] q4a8u_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_1_d[3:1])
      3'd0:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd1,
                                                         \call_f''''''''_f''''''''_goMux2_d };
      3'd1:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd2,
                                                         blae4_1_1_argbuf_d};
      3'd2:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd4,
                                                         trae3_2_1_argbuf_d};
      3'd3:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd8,
                                                         tlae2_3_1_argbuf_d};
      3'd4:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd16,
                                                         brae5_1_argbuf_d};
      default:
        {q4a8u_goMux_mux_onehot, q4a8u_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4a8u_goMux_mux_d = {q4a8u_goMux_mux_mux[16:1],
                              (q4a8u_goMux_mux_mux[0] && go_14_goMux_choice_1_d[0])};
  assign go_14_goMux_choice_1_r = (q4a8u_goMux_mux_d[0] && q4a8u_goMux_mux_r);
  assign {brae5_1_argbuf_r,
          tlae2_3_1_argbuf_r,
          trae3_2_1_argbuf_r,
          blae4_1_1_argbuf_r,
          \call_f''''''''_f''''''''_goMux2_r } = (go_14_goMux_choice_1_r ? q4a8u_goMux_mux_onehot :
                                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf''''''''_f'''''''') : (go_14_goMux_choice_2,C5) [(call_f''''''''_f''''''''_goMux3,Pointer_CTf''''''''_f''''''''),
                                                                    (sca2_1_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (sca1_1_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (sca0_1_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (sca3_1_1_argbuf,Pointer_CTf''''''''_f'''''''')] > (sc_0_1_goMux_mux,Pointer_CTf''''''''_f'''''''') */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f''''''''_f''''''''_goMux3_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_14_goMux_choice_2_d[0])};
  assign go_14_goMux_choice_2_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f''''''''_f''''''''_goMux3_r } = (go_14_goMux_choice_2_r ? sc_0_1_goMux_mux_onehot :
                                                  5'd0);
  
  /* fork (Ty C5) : (go_15_goMux_choice,C5) > [(go_15_goMux_choice_1,C5),
                                          (go_15_goMux_choice_2,C5),
                                          (go_15_goMux_choice_3,C5)] */
  logic [2:0] go_15_goMux_choice_emitted;
  logic [2:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[3:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[3:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_3_d = {go_15_goMux_choice_d[3:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[2]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_3_d[0],
                                                                   go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_3_r,
                                                                                                 go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 3'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 3'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_15_goMux_choice_1,C5) [(call_f_f_goMux2,Pointer_QTree_Int),
                                                        (q3aep_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2aeo_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1aen_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m1ae6_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1ae6_goMux_mux_mux;
  logic [4:0] m1ae6_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[3:1])
      3'd0:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd1,
                                                         call_f_f_goMux2_d};
      3'd1:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd2,
                                                         q3aep_1_1_argbuf_d};
      3'd2:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd4,
                                                         q2aeo_2_1_argbuf_d};
      3'd3:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd8,
                                                         q1aen_3_1_argbuf_d};
      3'd4:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd16,
                                                         lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_d};
      default:
        {m1ae6_goMux_mux_onehot, m1ae6_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1ae6_goMux_mux_d = {m1ae6_goMux_mux_mux[16:1],
                              (m1ae6_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (m1ae6_goMux_mux_d[0] && m1ae6_goMux_mux_r);
  assign {lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_r,
          q1aen_3_1_argbuf_r,
          q2aeo_2_1_argbuf_r,
          q3aep_1_1_argbuf_r,
          call_f_f_goMux2_r} = (go_15_goMux_choice_1_r ? m1ae6_goMux_mux_onehot :
                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_15_goMux_choice_2,C5) [(call_f_f_goMux3,Pointer_QTree_Int),
                                                        (t3aeu_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2aet_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1aes_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4aev_1_argbuf,Pointer_QTree_Int)] > (m2ae7_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2ae7_goMux_mux_mux;
  logic [4:0] m2ae7_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[3:1])
      3'd0:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd1,
                                                         call_f_f_goMux3_d};
      3'd1:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd2,
                                                         t3aeu_1_1_argbuf_d};
      3'd2:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd4,
                                                         t2aet_2_1_argbuf_d};
      3'd3:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd8,
                                                         t1aes_3_1_argbuf_d};
      3'd4:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd16,
                                                         t4aev_1_argbuf_d};
      default:
        {m2ae7_goMux_mux_onehot, m2ae7_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ae7_goMux_mux_d = {m2ae7_goMux_mux_mux[16:1],
                              (m2ae7_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (m2ae7_goMux_mux_d[0] && m2ae7_goMux_mux_r);
  assign {t4aev_1_argbuf_r,
          t1aes_3_1_argbuf_r,
          t2aet_2_1_argbuf_r,
          t3aeu_1_1_argbuf_r,
          call_f_f_goMux3_r} = (go_15_goMux_choice_2_r ? m2ae7_goMux_mux_onehot :
                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf_f) : (go_15_goMux_choice_3,C5) [(call_f_f_goMux4,Pointer_CTf_f),
                                                    (sca2_2_1_argbuf,Pointer_CTf_f),
                                                    (sca1_2_1_argbuf,Pointer_CTf_f),
                                                    (sca0_2_1_argbuf,Pointer_CTf_f),
                                                    (sca3_2_1_argbuf,Pointer_CTf_f)] > (sc_0_2_goMux_mux,Pointer_CTf_f) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_f_f_goMux4_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_15_goMux_choice_3_d[0])};
  assign go_15_goMux_choice_3_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_f_f_goMux4_r} = (go_15_goMux_choice_3_r ? sc_0_2_goMux_mux_onehot :
                                5'd0);
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(go_16_1MyTrue,MyBool)] > (lizzieLet0_1_1QVal_Bool,QTree_Bool) */
  assign lizzieLet0_1_1QVal_Bool_d = QVal_Bool_dc((& {go_16_1MyTrue_d[0]}), go_16_1MyTrue_d);
  assign {go_16_1MyTrue_r} = {1 {(lizzieLet0_1_1QVal_Bool_r && lizzieLet0_1_1QVal_Bool_d[0])}};
  
  /* dcon (Ty CTf''''''''_f'''''''',
      Dcon Lf''''''''_f''''''''sbos) : [(go_17_1,Go)] > (go_17_1Lf''''''''_f''''''''sbos,CTf''''''''_f'''''''') */
  assign \go_17_1Lf''''''''_f''''''''sbos_d  = \Lf''''''''_f''''''''sbos_dc ((& {go_17_1_d[0]}), go_17_1_d);
  assign {go_17_1_r} = {1 {(\go_17_1Lf''''''''_f''''''''sbos_r  && \go_17_1Lf''''''''_f''''''''sbos_d [0])}};
  
  /* buf (Ty CTf''''''''_f'''''''') : (go_17_1Lf''''''''_f''''''''sbos,CTf''''''''_f'''''''') > (lizzieLet42_1_argbuf,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \go_17_1Lf''''''''_f''''''''sbos_bufchan_d ;
  logic \go_17_1Lf''''''''_f''''''''sbos_bufchan_r ;
  assign \go_17_1Lf''''''''_f''''''''sbos_r  = ((! \go_17_1Lf''''''''_f''''''''sbos_bufchan_d [0]) || \go_17_1Lf''''''''_f''''''''sbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_17_1Lf''''''''_f''''''''sbos_bufchan_d  <= {67'd0, 1'd0};
    else
      if (\go_17_1Lf''''''''_f''''''''sbos_r )
        \go_17_1Lf''''''''_f''''''''sbos_bufchan_d  <= \go_17_1Lf''''''''_f''''''''sbos_d ;
  \CTf''''''''_f''''''''_t  \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf ;
  assign \go_17_1Lf''''''''_f''''''''sbos_bufchan_r  = (! \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf [0]);
  assign lizzieLet42_1_argbuf_d = (\go_17_1Lf''''''''_f''''''''sbos_bufchan_buf [0] ? \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf  :
                                   \go_17_1Lf''''''''_f''''''''sbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf  <= {67'd0, 1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf [0]))
        \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf  <= {67'd0, 1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf [0])))
        \go_17_1Lf''''''''_f''''''''sbos_bufchan_buf  <= \go_17_1Lf''''''''_f''''''''sbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_17_2,Go) > (go_17_2_argbuf,Go) */
  Go_t go_17_2_bufchan_d;
  logic go_17_2_bufchan_r;
  assign go_17_2_r = ((! go_17_2_bufchan_d[0]) || go_17_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_2_bufchan_d <= 1'd0;
    else if (go_17_2_r) go_17_2_bufchan_d <= go_17_2_d;
  Go_t go_17_2_bufchan_buf;
  assign go_17_2_bufchan_r = (! go_17_2_bufchan_buf[0]);
  assign go_17_2_argbuf_d = (go_17_2_bufchan_buf[0] ? go_17_2_bufchan_buf :
                             go_17_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_2_bufchan_buf <= 1'd0;
    else
      if ((go_17_2_argbuf_r && go_17_2_bufchan_buf[0]))
        go_17_2_bufchan_buf <= 1'd0;
      else if (((! go_17_2_argbuf_r) && (! go_17_2_bufchan_buf[0])))
        go_17_2_bufchan_buf <= go_17_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''',
      Dcon TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''') : [(go_17_2_argbuf,Go),
                                                                         (q4a8u_1_1_argbuf,Pointer_QTree_Int),
                                                                         (lizzieLet4_1_1_argbuf,Pointer_CTf''''''''_f'''''''')] > (call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1,TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f'''''''') */
  assign \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d  = \TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_dc ((& {go_17_2_argbuf_d[0],
                                                                                                                                                                      q4a8u_1_1_argbuf_d[0],
                                                                                                                                                                      lizzieLet4_1_1_argbuf_d[0]}), go_17_2_argbuf_d, q4a8u_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_17_2_argbuf_r,
          q4a8u_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {3 {(\call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_r  && \call_f''''''''_f''''''''TupGo___Pointer_QTree_Int___Pointer_CTf''''''''_f''''''''_1_d [0])}};
  
  /* dcon (Ty CTf_f,
      Dcon Lf_fsbos) : [(go_18_1,Go)] > (go_18_1Lf_fsbos,CTf_f) */
  assign go_18_1Lf_fsbos_d = Lf_fsbos_dc((& {go_18_1_d[0]}), go_18_1_d);
  assign {go_18_1_r} = {1 {(go_18_1Lf_fsbos_r && go_18_1Lf_fsbos_d[0])}};
  
  /* buf (Ty CTf_f) : (go_18_1Lf_fsbos,CTf_f) > (lizzieLet43_1_argbuf,CTf_f) */
  CTf_f_t go_18_1Lf_fsbos_bufchan_d;
  logic go_18_1Lf_fsbos_bufchan_r;
  assign go_18_1Lf_fsbos_r = ((! go_18_1Lf_fsbos_bufchan_d[0]) || go_18_1Lf_fsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_1Lf_fsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_18_1Lf_fsbos_r)
        go_18_1Lf_fsbos_bufchan_d <= go_18_1Lf_fsbos_d;
  CTf_f_t go_18_1Lf_fsbos_bufchan_buf;
  assign go_18_1Lf_fsbos_bufchan_r = (! go_18_1Lf_fsbos_bufchan_buf[0]);
  assign lizzieLet43_1_argbuf_d = (go_18_1Lf_fsbos_bufchan_buf[0] ? go_18_1Lf_fsbos_bufchan_buf :
                                   go_18_1Lf_fsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_1Lf_fsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && go_18_1Lf_fsbos_bufchan_buf[0]))
        go_18_1Lf_fsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! go_18_1Lf_fsbos_bufchan_buf[0])))
        go_18_1Lf_fsbos_bufchan_buf <= go_18_1Lf_fsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_18_2,Go) > (go_18_2_argbuf,Go) */
  Go_t go_18_2_bufchan_d;
  logic go_18_2_bufchan_r;
  assign go_18_2_r = ((! go_18_2_bufchan_d[0]) || go_18_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_2_bufchan_d <= 1'd0;
    else if (go_18_2_r) go_18_2_bufchan_d <= go_18_2_d;
  Go_t go_18_2_bufchan_buf;
  assign go_18_2_bufchan_r = (! go_18_2_bufchan_buf[0]);
  assign go_18_2_argbuf_d = (go_18_2_bufchan_buf[0] ? go_18_2_bufchan_buf :
                             go_18_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_2_bufchan_buf <= 1'd0;
    else
      if ((go_18_2_argbuf_r && go_18_2_bufchan_buf[0]))
        go_18_2_bufchan_buf <= 1'd0;
      else if (((! go_18_2_argbuf_r) && (! go_18_2_bufchan_buf[0])))
        go_18_2_bufchan_buf <= go_18_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f) : [(go_18_2_argbuf,Go),
                                                                             (m1ae6_1_1_argbuf,Pointer_QTree_Int),
                                                                             (m2ae7_1_1_argbuf,Pointer_QTree_Int),
                                                                             (lizzieLet17_1_1_argbuf,Pointer_CTf_f)] > (call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f) */
  assign call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_dc((& {go_18_2_argbuf_d[0],
                                                                                                                                                          m1ae6_1_1_argbuf_d[0],
                                                                                                                                                          m2ae7_1_1_argbuf_d[0],
                                                                                                                                                          lizzieLet17_1_1_argbuf_d[0]}), go_18_2_argbuf_d, m1ae6_1_1_argbuf_d, m2ae7_1_1_argbuf_d, lizzieLet17_1_1_argbuf_d);
  assign {go_18_2_argbuf_r,
          m1ae6_1_1_argbuf_r,
          m2ae7_1_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r} = {4 {(call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_r && call_f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CTf_f_1_d[0])}};
  
  /* fork (Ty C4) : (go_19_goMux_choice,C4) > [(go_19_goMux_choice_1,C4),
                                          (go_19_goMux_choice_2,C4)] */
  logic [1:0] go_19_goMux_choice_emitted;
  logic [1:0] go_19_goMux_choice_done;
  assign go_19_goMux_choice_1_d = {go_19_goMux_choice_d[2:1],
                                   (go_19_goMux_choice_d[0] && (! go_19_goMux_choice_emitted[0]))};
  assign go_19_goMux_choice_2_d = {go_19_goMux_choice_d[2:1],
                                   (go_19_goMux_choice_d[0] && (! go_19_goMux_choice_emitted[1]))};
  assign go_19_goMux_choice_done = (go_19_goMux_choice_emitted | ({go_19_goMux_choice_2_d[0],
                                                                   go_19_goMux_choice_1_d[0]} & {go_19_goMux_choice_2_r,
                                                                                                 go_19_goMux_choice_1_r}));
  assign go_19_goMux_choice_r = (& go_19_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_19_goMux_choice_emitted <= 2'd0;
    else
      go_19_goMux_choice_emitted <= (go_19_goMux_choice_r ? 2'd0 :
                                     go_19_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_19_goMux_choice_1,C4) [(lizzieLet18_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet19_1_argbuf,Int#),
                                           (lizzieLet18_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_19_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet18_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet19_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet18_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_19_goMux_choice_1_d[0])};
  assign go_19_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet18_1_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet18_1_argbuf_r} = (go_19_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz) : (go_19_goMux_choice_2,C4) [(lizzieLet1_4QNone_Bool_1_argbuf,Pointer_CT$wnnz),
                                                      (sc_0_6_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet1_4QVal_Bool_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet1_4QError_Bool_1_argbuf,Pointer_CT$wnnz)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_19_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet1_4QNone_Bool_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet1_4QVal_Bool_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet1_4QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_19_goMux_choice_2_d[0])};
  assign go_19_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet1_4QError_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet1_4QNone_Bool_1_argbuf_r} = (go_19_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                                4'd0);
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_1_argbuf,Go),
                                                             (m1aex_0,Pointer_QTree_Int),
                                                             (m2aey_1,Pointer_QTree_Int)] > (f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_1_argbuf_d[0],
                                                                                                                     m1aex_0_d[0],
                                                                                                                     m2aey_1_d[0]}), go_1_argbuf_d, m1aex_0_d, m2aey_1_d);
  assign {go_1_argbuf_r,
          m1aex_0_r,
          m2aey_1_r} = {3 {(f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r && f_fTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_2,Go) > (go_2_argbuf,Go) */
  Go_t go_2_bufchan_d;
  logic go_2_bufchan_r;
  assign go_2_r = ((! go_2_bufchan_d[0]) || go_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_d <= 1'd0;
    else if (go_2_r) go_2_bufchan_d <= go_2_d;
  Go_t go_2_bufchan_buf;
  assign go_2_bufchan_r = (! go_2_bufchan_buf[0]);
  assign go_2_argbuf_d = (go_2_bufchan_buf[0] ? go_2_bufchan_buf :
                          go_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_buf <= 1'd0;
    else
      if ((go_2_argbuf_r && go_2_bufchan_buf[0]))
        go_2_bufchan_buf <= 1'd0;
      else if (((! go_2_argbuf_r) && (! go_2_bufchan_buf[0])))
        go_2_bufchan_buf <= go_2_bufchan_d;
  
  /* fork (Ty C5) : (go_20_goMux_choice,C5) > [(go_20_goMux_choice_1,C5),
                                          (go_20_goMux_choice_2,C5)] */
  logic [1:0] go_20_goMux_choice_emitted;
  logic [1:0] go_20_goMux_choice_done;
  assign go_20_goMux_choice_1_d = {go_20_goMux_choice_d[3:1],
                                   (go_20_goMux_choice_d[0] && (! go_20_goMux_choice_emitted[0]))};
  assign go_20_goMux_choice_2_d = {go_20_goMux_choice_d[3:1],
                                   (go_20_goMux_choice_d[0] && (! go_20_goMux_choice_emitted[1]))};
  assign go_20_goMux_choice_done = (go_20_goMux_choice_emitted | ({go_20_goMux_choice_2_d[0],
                                                                   go_20_goMux_choice_1_d[0]} & {go_20_goMux_choice_2_r,
                                                                                                 go_20_goMux_choice_1_r}));
  assign go_20_goMux_choice_r = (& go_20_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_20_goMux_choice_emitted <= 2'd0;
    else
      go_20_goMux_choice_emitted <= (go_20_goMux_choice_r ? 2'd0 :
                                     go_20_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_20_goMux_choice_1,C5) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet8_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [4:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_20_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet8_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_20_goMux_choice_1_d[0])};
  assign go_20_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_20_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf''''''''_f'''''''') : (go_20_goMux_choice_2,C5) [(lizzieLet3_4QNone_Int_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (sc_0_10_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (lizzieLet7_2MyFalse_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (lizzieLet7_2MyTrue_1_argbuf,Pointer_CTf''''''''_f''''''''),
                                                                    (lizzieLet3_4QError_Int_1_argbuf,Pointer_CTf''''''''_f'''''''')] > (scfarg_0_1_goMux_mux,Pointer_CTf''''''''_f'''''''') */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [4:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_20_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet3_4QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   sc_0_10_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet7_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet7_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet3_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_20_goMux_choice_2_d[0])};
  assign go_20_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet3_4QError_Int_1_argbuf_r,
          lizzieLet7_2MyTrue_1_argbuf_r,
          lizzieLet7_2MyFalse_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet3_4QNone_Int_1_argbuf_r} = (go_20_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               5'd0);
  
  /* fork (Ty C16) : (go_21_goMux_choice,C16) > [(go_21_goMux_choice_1,C16),
                                            (go_21_goMux_choice_2,C16)] */
  logic [1:0] go_21_goMux_choice_emitted;
  logic [1:0] go_21_goMux_choice_done;
  assign go_21_goMux_choice_1_d = {go_21_goMux_choice_d[4:1],
                                   (go_21_goMux_choice_d[0] && (! go_21_goMux_choice_emitted[0]))};
  assign go_21_goMux_choice_2_d = {go_21_goMux_choice_d[4:1],
                                   (go_21_goMux_choice_d[0] && (! go_21_goMux_choice_emitted[1]))};
  assign go_21_goMux_choice_done = (go_21_goMux_choice_emitted | ({go_21_goMux_choice_2_d[0],
                                                                   go_21_goMux_choice_1_d[0]} & {go_21_goMux_choice_2_r,
                                                                                                 go_21_goMux_choice_1_r}));
  assign go_21_goMux_choice_r = (& go_21_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_21_goMux_choice_emitted <= 2'd0;
    else
      go_21_goMux_choice_emitted <= (go_21_goMux_choice_r ? 2'd0 :
                                     go_21_goMux_choice_done);
  
  /* mux (Ty C16,
     Ty Pointer_QTree_Bool) : (go_21_goMux_choice_1,C16) [(lizzieLet5_1_1_argbuf,Pointer_QTree_Bool),
                                                          (contRet_0_2_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet18_2_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet26_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet9_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet31_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet10_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet11_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet12_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet13_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet14_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet15_1_1_argbuf,Pointer_QTree_Bool),
                                                          (lizzieLet16_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [15:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_21_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd1,
                                                                   lizzieLet5_1_1_argbuf_d};
      4'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd2,
                                                                   contRet_0_2_1_argbuf_d};
      4'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd4,
                                                                   lizzieLet18_2_1_argbuf_d};
      4'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd8,
                                                                   lizzieLet6_1_1_argbuf_d};
      4'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd16,
                                                                   lizzieLet7_1_1_argbuf_d};
      4'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd32,
                                                                   lizzieLet8_1_1_argbuf_d};
      4'd6:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd64,
                                                                   lizzieLet26_1_argbuf_d};
      4'd7:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd128,
                                                                   lizzieLet9_1_1_argbuf_d};
      4'd8:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd256,
                                                                   lizzieLet31_1_argbuf_d};
      4'd9:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd512,
                                                                   lizzieLet10_1_1_argbuf_d};
      4'd10:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd1024, lizzieLet11_1_1_argbuf_d};
      4'd11:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd2048, lizzieLet12_1_1_argbuf_d};
      4'd12:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd4096, lizzieLet13_1_1_argbuf_d};
      4'd13:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd8192, lizzieLet14_1_1_argbuf_d};
      4'd14:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd16384, lizzieLet15_1_1_argbuf_d};
      4'd15:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {16'd32768, lizzieLet16_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {16'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_21_goMux_choice_1_d[0])};
  assign go_21_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet16_1_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          lizzieLet18_2_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = (go_21_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      16'd0);
  
  /* mux (Ty C16,
     Ty Pointer_CTf_f) : (go_21_goMux_choice_2,C16) [(lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf,Pointer_CTf_f),
                                                     (sc_0_14_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet17_2MyFalse_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet17_2MyTrue_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QNone_Int_4QError_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet25_2MyFalse_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet25_2MyTrue_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet30_2MyFalse_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet30_2MyTrue_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_4QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f),
                                                     (lizzieLet12_5QError_Int_1_argbuf,Pointer_CTf_f)] > (scfarg_0_2_goMux_mux,Pointer_CTf_f) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [15:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_21_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd1,
                                                                   lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_d};
      4'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd2,
                                                                   sc_0_14_1_argbuf_d};
      4'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd4,
                                                                   lizzieLet17_2MyFalse_1_argbuf_d};
      4'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd8,
                                                                   lizzieLet17_2MyTrue_1_argbuf_d};
      4'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd16,
                                                                   lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_d};
      4'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd32,
                                                                   lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd64,
                                                                   lizzieLet25_2MyFalse_1_argbuf_d};
      4'd7:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd128,
                                                                   lizzieLet25_2MyTrue_1_argbuf_d};
      4'd8:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd256,
                                                                   lizzieLet30_2MyFalse_1_argbuf_d};
      4'd9:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd512,
                                                                   lizzieLet30_2MyTrue_1_argbuf_d};
      4'd10:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd1024,
                                      lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_d};
      4'd11:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd2048,
                                      lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_d};
      4'd12:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd4096,
                                      lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_d};
      4'd13:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd8192,
                                      lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_d};
      4'd14:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd16384,
                                      lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_d};
      4'd15:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {16'd32768,
                                      lizzieLet12_5QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {16'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_21_goMux_choice_2_d[0])};
  assign go_21_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet12_5QError_Int_1_argbuf_r,
          lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_r,
          lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_r,
          lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_r,
          lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_r,
          lizzieLet30_2MyTrue_1_argbuf_r,
          lizzieLet30_2MyFalse_1_argbuf_r,
          lizzieLet25_2MyTrue_1_argbuf_r,
          lizzieLet25_2MyFalse_1_argbuf_r,
          lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_r,
          lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_r,
          lizzieLet17_2MyTrue_1_argbuf_r,
          lizzieLet17_2MyFalse_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_r} = (go_21_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                           16'd0);
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool) : [(go_2_argbuf,Go),
                                          (es_0_1_argbuf,Pointer_QTree_Bool)] > ($wnnzTupGo___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool) */
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_d  = TupGo___Pointer_QTree_Bool_dc((& {go_2_argbuf_d[0],
                                                                                   es_0_1_argbuf_d[0]}), go_2_argbuf_d, es_0_1_argbuf_d);
  assign {go_2_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnzTupGo___Pointer_QTree_Bool_1_r  && \$wnnzTupGo___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet0_1_1QVal_Bool,QTree_Bool) > (lizzieLet41_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_d;
  logic lizzieLet0_1_1QVal_Bool_bufchan_r;
  assign lizzieLet0_1_1QVal_Bool_r = ((! lizzieLet0_1_1QVal_Bool_bufchan_d[0]) || lizzieLet0_1_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet0_1_1QVal_Bool_r)
        lizzieLet0_1_1QVal_Bool_bufchan_d <= lizzieLet0_1_1QVal_Bool_d;
  QTree_Bool_t lizzieLet0_1_1QVal_Bool_bufchan_buf;
  assign lizzieLet0_1_1QVal_Bool_bufchan_r = (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet41_1_argbuf_d = (lizzieLet0_1_1QVal_Bool_bufchan_buf[0] ? lizzieLet0_1_1QVal_Bool_bufchan_buf :
                                   lizzieLet0_1_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && lizzieLet0_1_1QVal_Bool_bufchan_buf[0]))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! lizzieLet0_1_1QVal_Bool_bufchan_buf[0])))
        lizzieLet0_1_1QVal_Bool_bufchan_buf <= lizzieLet0_1_1QVal_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_1QNode_Int,QTree_Int) > [(q1aen_destruct,Pointer_QTree_Int),
                                                                  (q2aeo_destruct,Pointer_QTree_Int),
                                                                  (q3aep_destruct,Pointer_QTree_Int),
                                                                  (q4aeq_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_1QNode_Int_done;
  assign q1aen_destruct_d = {lizzieLet12_1QNode_Int_d[18:3],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[0]))};
  assign q2aeo_destruct_d = {lizzieLet12_1QNode_Int_d[34:19],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[1]))};
  assign q3aep_destruct_d = {lizzieLet12_1QNode_Int_d[50:35],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[2]))};
  assign q4aeq_destruct_d = {lizzieLet12_1QNode_Int_d[66:51],
                             (lizzieLet12_1QNode_Int_d[0] && (! lizzieLet12_1QNode_Int_emitted[3]))};
  assign lizzieLet12_1QNode_Int_done = (lizzieLet12_1QNode_Int_emitted | ({q4aeq_destruct_d[0],
                                                                           q3aep_destruct_d[0],
                                                                           q2aeo_destruct_d[0],
                                                                           q1aen_destruct_d[0]} & {q4aeq_destruct_r,
                                                                                                   q3aep_destruct_r,
                                                                                                   q2aeo_destruct_r,
                                                                                                   q1aen_destruct_r}));
  assign lizzieLet12_1QNode_Int_r = (& lizzieLet12_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_1QNode_Int_emitted <= (lizzieLet12_1QNode_Int_r ? 4'd0 :
                                         lizzieLet12_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_1QVal_Int,QTree_Int) > [(v1aee_destruct,Int)] */
  assign v1aee_destruct_d = {lizzieLet12_1QVal_Int_d[34:3],
                             lizzieLet12_1QVal_Int_d[0]};
  assign lizzieLet12_1QVal_Int_r = v1aee_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_2,QTree_Int) (lizzieLet12_1,QTree_Int) > [(_31,QTree_Int),
                                                                              (lizzieLet12_1QVal_Int,QTree_Int),
                                                                              (lizzieLet12_1QNode_Int,QTree_Int),
                                                                              (_30,QTree_Int)] */
  logic [3:0] lizzieLet12_1_onehotd;
  always_comb
    if ((lizzieLet12_2_d[0] && lizzieLet12_1_d[0]))
      unique case (lizzieLet12_2_d[2:1])
        2'd0: lizzieLet12_1_onehotd = 4'd1;
        2'd1: lizzieLet12_1_onehotd = 4'd2;
        2'd2: lizzieLet12_1_onehotd = 4'd4;
        2'd3: lizzieLet12_1_onehotd = 4'd8;
        default: lizzieLet12_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_1_onehotd = 4'd0;
  assign _31_d = {lizzieLet12_1_d[66:1], lizzieLet12_1_onehotd[0]};
  assign lizzieLet12_1QVal_Int_d = {lizzieLet12_1_d[66:1],
                                    lizzieLet12_1_onehotd[1]};
  assign lizzieLet12_1QNode_Int_d = {lizzieLet12_1_d[66:1],
                                     lizzieLet12_1_onehotd[2]};
  assign _30_d = {lizzieLet12_1_d[66:1], lizzieLet12_1_onehotd[3]};
  assign lizzieLet12_1_r = (| (lizzieLet12_1_onehotd & {_30_r,
                                                        lizzieLet12_1QNode_Int_r,
                                                        lizzieLet12_1QVal_Int_r,
                                                        _31_r}));
  assign lizzieLet12_2_r = lizzieLet12_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_3,QTree_Int) (go_15_goMux_data,Go) > [(lizzieLet12_3QNone_Int,Go),
                                                                   (lizzieLet12_3QVal_Int,Go),
                                                                   (lizzieLet12_3QNode_Int,Go),
                                                                   (lizzieLet12_3QError_Int,Go)] */
  logic [3:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet12_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet12_3_d[2:1])
        2'd0: go_15_goMux_data_onehotd = 4'd1;
        2'd1: go_15_goMux_data_onehotd = 4'd2;
        2'd2: go_15_goMux_data_onehotd = 4'd4;
        2'd3: go_15_goMux_data_onehotd = 4'd8;
        default: go_15_goMux_data_onehotd = 4'd0;
      endcase
    else go_15_goMux_data_onehotd = 4'd0;
  assign lizzieLet12_3QNone_Int_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet12_3QVal_Int_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet12_3QNode_Int_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet12_3QError_Int_d = go_15_goMux_data_onehotd[3];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet12_3QError_Int_r,
                                                              lizzieLet12_3QNode_Int_r,
                                                              lizzieLet12_3QVal_Int_r,
                                                              lizzieLet12_3QNone_Int_r}));
  assign lizzieLet12_3_r = go_15_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet12_3QError_Int,Go) > [(lizzieLet12_3QError_Int_1,Go),
                                               (lizzieLet12_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_3QError_Int_emitted;
  logic [1:0] lizzieLet12_3QError_Int_done;
  assign lizzieLet12_3QError_Int_1_d = (lizzieLet12_3QError_Int_d[0] && (! lizzieLet12_3QError_Int_emitted[0]));
  assign lizzieLet12_3QError_Int_2_d = (lizzieLet12_3QError_Int_d[0] && (! lizzieLet12_3QError_Int_emitted[1]));
  assign lizzieLet12_3QError_Int_done = (lizzieLet12_3QError_Int_emitted | ({lizzieLet12_3QError_Int_2_d[0],
                                                                             lizzieLet12_3QError_Int_1_d[0]} & {lizzieLet12_3QError_Int_2_r,
                                                                                                                lizzieLet12_3QError_Int_1_r}));
  assign lizzieLet12_3QError_Int_r = (& lizzieLet12_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_3QError_Int_emitted <= (lizzieLet12_3QError_Int_r ? 2'd0 :
                                          lizzieLet12_3QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_3QError_Int_1,Go)] > (lizzieLet12_3QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_3QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_3QError_Int_1_d[0]}), lizzieLet12_3QError_Int_1_d);
  assign {lizzieLet12_3QError_Int_1_r} = {1 {(lizzieLet12_3QError_Int_1QError_Bool_r && lizzieLet12_3QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_3QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet40_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_3QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_3QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_3QError_Int_1QError_Bool_r = ((! lizzieLet12_3QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_3QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_3QError_Int_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet12_3QError_Int_1QError_Bool_r)
        lizzieLet12_3QError_Int_1QError_Bool_bufchan_d <= lizzieLet12_3QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_3QError_Int_1QError_Bool_bufchan_r = (! lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet40_1_argbuf_d = (lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_3QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_3QError_Int_1QError_Bool_bufchan_buf <= lizzieLet12_3QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_3QError_Int_2,Go) > (lizzieLet12_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_3QError_Int_2_bufchan_d;
  logic lizzieLet12_3QError_Int_2_bufchan_r;
  assign lizzieLet12_3QError_Int_2_r = ((! lizzieLet12_3QError_Int_2_bufchan_d[0]) || lizzieLet12_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_3QError_Int_2_r)
        lizzieLet12_3QError_Int_2_bufchan_d <= lizzieLet12_3QError_Int_2_d;
  Go_t lizzieLet12_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_3QError_Int_2_bufchan_r = (! lizzieLet12_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_3QError_Int_2_argbuf_d = (lizzieLet12_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_3QError_Int_2_bufchan_buf :
                                               lizzieLet12_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_3QError_Int_2_argbuf_r && lizzieLet12_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_3QError_Int_2_argbuf_r) && (! lizzieLet12_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_3QError_Int_2_bufchan_buf <= lizzieLet12_3QError_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_4,QTree_Int) (readPointer_QTree_Intm2ae7_1_argbuf_rwb,QTree_Int) > [(lizzieLet12_4QNone_Int,QTree_Int),
                                                                                                        (lizzieLet12_4QVal_Int,QTree_Int),
                                                                                                        (lizzieLet12_4QNode_Int,QTree_Int),
                                                                                                        (_29,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet12_4_d[0] && readPointer_QTree_Intm2ae7_1_argbuf_rwb_d[0]))
      unique case (lizzieLet12_4_d[2:1])
        2'd0: readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd = 4'd0;
  assign lizzieLet12_4QNone_Int_d = {readPointer_QTree_Intm2ae7_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet12_4QVal_Int_d = {readPointer_QTree_Intm2ae7_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet12_4QNode_Int_d = {readPointer_QTree_Intm2ae7_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd[2]};
  assign _29_d = {readPointer_QTree_Intm2ae7_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intm2ae7_1_argbuf_rwb_r = (| (readPointer_QTree_Intm2ae7_1_argbuf_rwb_onehotd & {_29_r,
                                                                                                            lizzieLet12_4QNode_Int_r,
                                                                                                            lizzieLet12_4QVal_Int_r,
                                                                                                            lizzieLet12_4QNone_Int_r}));
  assign lizzieLet12_4_r = readPointer_QTree_Intm2ae7_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_4QNode_Int,QTree_Int) > [(lizzieLet12_4QNode_Int_1,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_2,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_3,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_4,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_5,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_6,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_7,QTree_Int),
                                                            (lizzieLet12_4QNode_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet12_4QNode_Int_emitted;
  logic [7:0] lizzieLet12_4QNode_Int_done;
  assign lizzieLet12_4QNode_Int_1_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[0]))};
  assign lizzieLet12_4QNode_Int_2_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[1]))};
  assign lizzieLet12_4QNode_Int_3_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[2]))};
  assign lizzieLet12_4QNode_Int_4_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[3]))};
  assign lizzieLet12_4QNode_Int_5_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[4]))};
  assign lizzieLet12_4QNode_Int_6_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[5]))};
  assign lizzieLet12_4QNode_Int_7_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[6]))};
  assign lizzieLet12_4QNode_Int_8_d = {lizzieLet12_4QNode_Int_d[66:1],
                                       (lizzieLet12_4QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_emitted[7]))};
  assign lizzieLet12_4QNode_Int_done = (lizzieLet12_4QNode_Int_emitted | ({lizzieLet12_4QNode_Int_8_d[0],
                                                                           lizzieLet12_4QNode_Int_7_d[0],
                                                                           lizzieLet12_4QNode_Int_6_d[0],
                                                                           lizzieLet12_4QNode_Int_5_d[0],
                                                                           lizzieLet12_4QNode_Int_4_d[0],
                                                                           lizzieLet12_4QNode_Int_3_d[0],
                                                                           lizzieLet12_4QNode_Int_2_d[0],
                                                                           lizzieLet12_4QNode_Int_1_d[0]} & {lizzieLet12_4QNode_Int_8_r,
                                                                                                             lizzieLet12_4QNode_Int_7_r,
                                                                                                             lizzieLet12_4QNode_Int_6_r,
                                                                                                             lizzieLet12_4QNode_Int_5_r,
                                                                                                             lizzieLet12_4QNode_Int_4_r,
                                                                                                             lizzieLet12_4QNode_Int_3_r,
                                                                                                             lizzieLet12_4QNode_Int_2_r,
                                                                                                             lizzieLet12_4QNode_Int_1_r}));
  assign lizzieLet12_4QNode_Int_r = (& lizzieLet12_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_4QNode_Int_emitted <= 8'd0;
    else
      lizzieLet12_4QNode_Int_emitted <= (lizzieLet12_4QNode_Int_r ? 8'd0 :
                                         lizzieLet12_4QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_4QNode_Int_1QNode_Int,QTree_Int) > [(t1aes_destruct,Pointer_QTree_Int),
                                                                             (t2aet_destruct,Pointer_QTree_Int),
                                                                             (t3aeu_destruct,Pointer_QTree_Int),
                                                                             (t4aev_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_4QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_4QNode_Int_1QNode_Int_done;
  assign t1aes_destruct_d = {lizzieLet12_4QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet12_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_1QNode_Int_emitted[0]))};
  assign t2aet_destruct_d = {lizzieLet12_4QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet12_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_1QNode_Int_emitted[1]))};
  assign t3aeu_destruct_d = {lizzieLet12_4QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet12_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_1QNode_Int_emitted[2]))};
  assign t4aev_destruct_d = {lizzieLet12_4QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet12_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet12_4QNode_Int_1QNode_Int_done = (lizzieLet12_4QNode_Int_1QNode_Int_emitted | ({t4aev_destruct_d[0],
                                                                                                 t3aeu_destruct_d[0],
                                                                                                 t2aet_destruct_d[0],
                                                                                                 t1aes_destruct_d[0]} & {t4aev_destruct_r,
                                                                                                                         t3aeu_destruct_r,
                                                                                                                         t2aet_destruct_r,
                                                                                                                         t1aes_destruct_r}));
  assign lizzieLet12_4QNode_Int_1QNode_Int_r = (& lizzieLet12_4QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_4QNode_Int_1QNode_Int_emitted <= (lizzieLet12_4QNode_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_4QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_4QNode_Int_2,QTree_Int) (lizzieLet12_4QNode_Int_1,QTree_Int) > [(_28,QTree_Int),
                                                                                                    (_27,QTree_Int),
                                                                                                    (lizzieLet12_4QNode_Int_1QNode_Int,QTree_Int),
                                                                                                    (_26,QTree_Int)] */
  logic [3:0] lizzieLet12_4QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_2_d[0] && lizzieLet12_4QNode_Int_1_d[0]))
      unique case (lizzieLet12_4QNode_Int_2_d[2:1])
        2'd0: lizzieLet12_4QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_4QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_4QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_4QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet12_4QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_4QNode_Int_1_onehotd = 4'd0;
  assign _28_d = {lizzieLet12_4QNode_Int_1_d[66:1],
                  lizzieLet12_4QNode_Int_1_onehotd[0]};
  assign _27_d = {lizzieLet12_4QNode_Int_1_d[66:1],
                  lizzieLet12_4QNode_Int_1_onehotd[1]};
  assign lizzieLet12_4QNode_Int_1QNode_Int_d = {lizzieLet12_4QNode_Int_1_d[66:1],
                                                lizzieLet12_4QNode_Int_1_onehotd[2]};
  assign _26_d = {lizzieLet12_4QNode_Int_1_d[66:1],
                  lizzieLet12_4QNode_Int_1_onehotd[3]};
  assign lizzieLet12_4QNode_Int_1_r = (| (lizzieLet12_4QNode_Int_1_onehotd & {_26_r,
                                                                              lizzieLet12_4QNode_Int_1QNode_Int_r,
                                                                              _27_r,
                                                                              _28_r}));
  assign lizzieLet12_4QNode_Int_2_r = lizzieLet12_4QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_4QNode_Int_3,QTree_Int) (lizzieLet12_3QNode_Int,Go) > [(lizzieLet12_4QNode_Int_3QNone_Int,Go),
                                                                                    (lizzieLet12_4QNode_Int_3QVal_Int,Go),
                                                                                    (lizzieLet12_4QNode_Int_3QNode_Int,Go),
                                                                                    (lizzieLet12_4QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_3_d[0] && lizzieLet12_3QNode_Int_d[0]))
      unique case (lizzieLet12_4QNode_Int_3_d[2:1])
        2'd0: lizzieLet12_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_3QNone_Int_d = lizzieLet12_3QNode_Int_onehotd[0];
  assign lizzieLet12_4QNode_Int_3QVal_Int_d = lizzieLet12_3QNode_Int_onehotd[1];
  assign lizzieLet12_4QNode_Int_3QNode_Int_d = lizzieLet12_3QNode_Int_onehotd[2];
  assign lizzieLet12_4QNode_Int_3QError_Int_d = lizzieLet12_3QNode_Int_onehotd[3];
  assign lizzieLet12_3QNode_Int_r = (| (lizzieLet12_3QNode_Int_onehotd & {lizzieLet12_4QNode_Int_3QError_Int_r,
                                                                          lizzieLet12_4QNode_Int_3QNode_Int_r,
                                                                          lizzieLet12_4QNode_Int_3QVal_Int_r,
                                                                          lizzieLet12_4QNode_Int_3QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_3_r = lizzieLet12_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_4QNode_Int_3QError_Int,Go) > [(lizzieLet12_4QNode_Int_3QError_Int_1,Go),
                                                          (lizzieLet12_4QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_4QNode_Int_3QError_Int_done;
  assign lizzieLet12_4QNode_Int_3QError_Int_1_d = (lizzieLet12_4QNode_Int_3QError_Int_d[0] && (! lizzieLet12_4QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_4QNode_Int_3QError_Int_2_d = (lizzieLet12_4QNode_Int_3QError_Int_d[0] && (! lizzieLet12_4QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_4QNode_Int_3QError_Int_done = (lizzieLet12_4QNode_Int_3QError_Int_emitted | ({lizzieLet12_4QNode_Int_3QError_Int_2_d[0],
                                                                                                   lizzieLet12_4QNode_Int_3QError_Int_1_d[0]} & {lizzieLet12_4QNode_Int_3QError_Int_2_r,
                                                                                                                                                 lizzieLet12_4QNode_Int_3QError_Int_1_r}));
  assign lizzieLet12_4QNode_Int_3QError_Int_r = (& lizzieLet12_4QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QNode_Int_3QError_Int_emitted <= (lizzieLet12_4QNode_Int_3QError_Int_r ? 2'd0 :
                                                     lizzieLet12_4QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_4QNode_Int_3QError_Int_1,Go)] > (lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_4QNode_Int_3QError_Int_1_d[0]}), lizzieLet12_4QNode_Int_3QError_Int_1_d);
  assign {lizzieLet12_4QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_r && lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet39_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_r = ((! lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_r)
        lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d <= lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_r = (! lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_buf <= lizzieLet12_4QNode_Int_3QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QError_Int_2,Go) > (lizzieLet12_4QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QError_Int_2_r = ((! lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QError_Int_2_r)
        lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet12_4QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf :
                                                          lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_r && lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_4QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNode_Int,Go) > (lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNode_Int_r = ((! lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNode_Int_r)
        lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d <= lizzieLet12_4QNode_Int_3QNode_Int_d;
  Go_t lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet12_4QNode_Int_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int,Go) > [(lizzieLet12_4QNode_Int_3QNone_Int_1,Go),
                                                         (lizzieLet12_4QNode_Int_3QNone_Int_2,Go),
                                                         (lizzieLet12_4QNode_Int_3QNone_Int_3,Go),
                                                         (lizzieLet12_4QNode_Int_3QNone_Int_4,Go),
                                                         (lizzieLet12_4QNode_Int_3QNone_Int_5,Go)] */
  logic [4:0] lizzieLet12_4QNode_Int_3QNone_Int_emitted;
  logic [4:0] lizzieLet12_4QNode_Int_3QNone_Int_done;
  assign lizzieLet12_4QNode_Int_3QNone_Int_1_d = (lizzieLet12_4QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNode_Int_3QNone_Int_emitted[0]));
  assign lizzieLet12_4QNode_Int_3QNone_Int_2_d = (lizzieLet12_4QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNode_Int_3QNone_Int_emitted[1]));
  assign lizzieLet12_4QNode_Int_3QNone_Int_3_d = (lizzieLet12_4QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNode_Int_3QNone_Int_emitted[2]));
  assign lizzieLet12_4QNode_Int_3QNone_Int_4_d = (lizzieLet12_4QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNode_Int_3QNone_Int_emitted[3]));
  assign lizzieLet12_4QNode_Int_3QNone_Int_5_d = (lizzieLet12_4QNode_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNode_Int_3QNone_Int_emitted[4]));
  assign lizzieLet12_4QNode_Int_3QNone_Int_done = (lizzieLet12_4QNode_Int_3QNone_Int_emitted | ({lizzieLet12_4QNode_Int_3QNone_Int_5_d[0],
                                                                                                 lizzieLet12_4QNode_Int_3QNone_Int_4_d[0],
                                                                                                 lizzieLet12_4QNode_Int_3QNone_Int_3_d[0],
                                                                                                 lizzieLet12_4QNode_Int_3QNone_Int_2_d[0],
                                                                                                 lizzieLet12_4QNode_Int_3QNone_Int_1_d[0]} & {lizzieLet12_4QNode_Int_3QNone_Int_5_r,
                                                                                                                                              lizzieLet12_4QNode_Int_3QNone_Int_4_r,
                                                                                                                                              lizzieLet12_4QNode_Int_3QNone_Int_3_r,
                                                                                                                                              lizzieLet12_4QNode_Int_3QNone_Int_2_r,
                                                                                                                                              lizzieLet12_4QNode_Int_3QNone_Int_1_r}));
  assign lizzieLet12_4QNode_Int_3QNone_Int_r = (& lizzieLet12_4QNode_Int_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_emitted <= 5'd0;
    else
      lizzieLet12_4QNode_Int_3QNone_Int_emitted <= (lizzieLet12_4QNode_Int_3QNone_Int_r ? 5'd0 :
                                                    lizzieLet12_4QNode_Int_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int_1,Go) > (lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNone_Int_1_r = ((! lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNone_Int_1_r)
        lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d <= lizzieLet12_4QNode_Int_3QNone_Int_1_d;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_r = (! lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_buf <= lizzieLet12_4QNode_Int_3QNone_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf,Go),
                                         (lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int5,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_d[0],
                                                                                              lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_d[0]}), lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_d, lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_d);
  assign {lizzieLet12_4QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int5_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int_2,Go) > (lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNone_Int_2_r = ((! lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNone_Int_2_r)
        lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d <= lizzieLet12_4QNode_Int_3QNone_Int_2_d;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_r = (! lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_d = (lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_r && lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_buf <= lizzieLet12_4QNode_Int_3QNone_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf,Go),
                                         (lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int6,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_d[0],
                                                                                              lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_d[0]}), lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_d, lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_d);
  assign {lizzieLet12_4QNode_Int_3QNone_Int_2_argbuf_r,
          lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int6_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int_3,Go) > (lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNone_Int_3_r = ((! lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNone_Int_3_r)
        lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d <= lizzieLet12_4QNode_Int_3QNone_Int_3_d;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_r = (! lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_d = (lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_r && lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_buf <= lizzieLet12_4QNode_Int_3QNone_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf,Go),
                                         (lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int7,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_d[0],
                                                                                              lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_d[0]}), lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_d, lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_d);
  assign {lizzieLet12_4QNode_Int_3QNone_Int_3_argbuf_r,
          lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int7_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int_4,Go) > (lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNone_Int_4_r = ((! lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNone_Int_4_r)
        lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d <= lizzieLet12_4QNode_Int_3QNone_Int_4_d;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_r = (! lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_d = (lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_r && lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_buf <= lizzieLet12_4QNode_Int_3QNone_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf,Go),
                                         (lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int8,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int8_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_d[0],
                                                                                              lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_d[0]}), lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_d, lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_d);
  assign {lizzieLet12_4QNode_Int_3QNone_Int_4_argbuf_r,
          lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int8_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QNone_Int_5,Go) > (lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QNone_Int_5_r = ((! lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QNone_Int_5_r)
        lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d <= lizzieLet12_4QNode_Int_3QNone_Int_5_d;
  Go_t lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_r = (! lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_d = (lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_r && lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_r) && (! lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_buf <= lizzieLet12_4QNode_Int_3QNone_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_4QNode_Int_3QVal_Int,Go) > [(lizzieLet12_4QNode_Int_3QVal_Int_1,Go),
                                                        (lizzieLet12_4QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet12_4QNode_Int_3QVal_Int_done;
  assign lizzieLet12_4QNode_Int_3QVal_Int_1_d = (lizzieLet12_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet12_4QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet12_4QNode_Int_3QVal_Int_2_d = (lizzieLet12_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet12_4QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet12_4QNode_Int_3QVal_Int_done = (lizzieLet12_4QNode_Int_3QVal_Int_emitted | ({lizzieLet12_4QNode_Int_3QVal_Int_2_d[0],
                                                                                               lizzieLet12_4QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet12_4QNode_Int_3QVal_Int_2_r,
                                                                                                                                           lizzieLet12_4QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet12_4QNode_Int_3QVal_Int_r = (& lizzieLet12_4QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QNode_Int_3QVal_Int_emitted <= (lizzieLet12_4QNode_Int_3QVal_Int_r ? 2'd0 :
                                                   lizzieLet12_4QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_4QNode_Int_3QVal_Int_1,Go)] > (lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_4QNode_Int_3QVal_Int_1_d[0]}), lizzieLet12_4QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet12_4QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_r && lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool,QTree_Bool) > (lizzieLet37_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_r = ((! lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_r)
        lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d <= lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_r = (! lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet37_1_argbuf_d = (lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_buf <= lizzieLet12_4QNode_Int_3QVal_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QNode_Int_3QVal_Int_2,Go) > (lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet12_4QNode_Int_3QVal_Int_2_r = ((! lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNode_Int_3QVal_Int_2_r)
        lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet12_4QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf :
                                                        lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet12_4QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QNode_Int_4,QTree_Int) (lizzieLet12_5QNode_Int,Pointer_CTf_f) > [(lizzieLet12_4QNode_Int_4QNone_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNode_Int_4QVal_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNode_Int_4QNode_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNode_Int_4QError_Int,Pointer_CTf_f)] */
  logic [3:0] lizzieLet12_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_4_d[0] && lizzieLet12_5QNode_Int_d[0]))
      unique case (lizzieLet12_4QNode_Int_4_d[2:1])
        2'd0: lizzieLet12_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet12_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_4QNone_Int_d = {lizzieLet12_5QNode_Int_d[16:1],
                                                lizzieLet12_5QNode_Int_onehotd[0]};
  assign lizzieLet12_4QNode_Int_4QVal_Int_d = {lizzieLet12_5QNode_Int_d[16:1],
                                               lizzieLet12_5QNode_Int_onehotd[1]};
  assign lizzieLet12_4QNode_Int_4QNode_Int_d = {lizzieLet12_5QNode_Int_d[16:1],
                                                lizzieLet12_5QNode_Int_onehotd[2]};
  assign lizzieLet12_4QNode_Int_4QError_Int_d = {lizzieLet12_5QNode_Int_d[16:1],
                                                 lizzieLet12_5QNode_Int_onehotd[3]};
  assign lizzieLet12_5QNode_Int_r = (| (lizzieLet12_5QNode_Int_onehotd & {lizzieLet12_4QNode_Int_4QError_Int_r,
                                                                          lizzieLet12_4QNode_Int_4QNode_Int_r,
                                                                          lizzieLet12_4QNode_Int_4QVal_Int_r,
                                                                          lizzieLet12_4QNode_Int_4QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_4_r = lizzieLet12_5QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNode_Int_4QError_Int,Pointer_CTf_f) > (lizzieLet12_4QNode_Int_4QError_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QError_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_4QError_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_4QError_Int_r = ((! lizzieLet12_4QNode_Int_4QError_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_4QError_Int_r)
        lizzieLet12_4QNode_Int_4QError_Int_bufchan_d <= lizzieLet12_4QNode_Int_4QError_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_4QError_Int_bufchan_r = (! lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf :
                                                          lizzieLet12_4QNode_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_r && lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_4QError_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_4QError_Int_bufchan_buf <= lizzieLet12_4QNode_Int_4QError_Int_bufchan_d;
  
  /* dcon (Ty CTf_f,
      Dcon Lcall_f_f3) : [(lizzieLet12_4QNode_Int_4QNode_Int,Pointer_CTf_f),
                          (lizzieLet12_4QNode_Int_5QNode_Int,Pointer_QTree_Int),
                          (t1aes_destruct,Pointer_QTree_Int),
                          (lizzieLet12_4QNode_Int_6QNode_Int,Pointer_QTree_Int),
                          (t2aet_destruct,Pointer_QTree_Int),
                          (lizzieLet12_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                          (t3aeu_destruct,Pointer_QTree_Int)] > (lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3,CTf_f) */
  assign lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_d = Lcall_f_f3_dc((& {lizzieLet12_4QNode_Int_4QNode_Int_d[0],
                                                                                                                                                                                                           lizzieLet12_4QNode_Int_5QNode_Int_d[0],
                                                                                                                                                                                                           t1aes_destruct_d[0],
                                                                                                                                                                                                           lizzieLet12_4QNode_Int_6QNode_Int_d[0],
                                                                                                                                                                                                           t2aet_destruct_d[0],
                                                                                                                                                                                                           lizzieLet12_4QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                           t3aeu_destruct_d[0]}), lizzieLet12_4QNode_Int_4QNode_Int_d, lizzieLet12_4QNode_Int_5QNode_Int_d, t1aes_destruct_d, lizzieLet12_4QNode_Int_6QNode_Int_d, t2aet_destruct_d, lizzieLet12_4QNode_Int_7QNode_Int_d, t3aeu_destruct_d);
  assign {lizzieLet12_4QNode_Int_4QNode_Int_r,
          lizzieLet12_4QNode_Int_5QNode_Int_r,
          t1aes_destruct_r,
          lizzieLet12_4QNode_Int_6QNode_Int_r,
          t2aet_destruct_r,
          lizzieLet12_4QNode_Int_7QNode_Int_r,
          t3aeu_destruct_r} = {7 {(lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_r && lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_d[0])}};
  
  /* buf (Ty CTf_f) : (lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3,CTf_f) > (lizzieLet38_1_argbuf,CTf_f) */
  CTf_f_t lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d;
  logic lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_r;
  assign lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_r = ((! lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d[0]) || lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d <= {115'd0,
                                                                                                                                                                                                1'd0};
    else
      if (lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_r)
        lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d <= lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_d;
  CTf_f_t lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf;
  assign lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_r = (! lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf[0] ? lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf :
                                   lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                  1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                    1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_buf <= lizzieLet12_4QNode_Int_4QNode_Int_1lizzieLet12_4QNode_Int_5QNode_Int_1t1aes_1lizzieLet12_4QNode_Int_6QNode_Int_1t2aet_1lizzieLet12_4QNode_Int_7QNode_Int_1t3aeu_1Lcall_f_f3_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNode_Int_4QNone_Int,Pointer_CTf_f) > (lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_4QNone_Int_r = ((! lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_4QNone_Int_r)
        lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d <= lizzieLet12_4QNode_Int_4QNone_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet12_4QNode_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNode_Int_4QVal_Int,Pointer_CTf_f) > (lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_4QVal_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_4QVal_Int_r = ((! lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_4QVal_Int_r)
        lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d <= lizzieLet12_4QNode_Int_4QVal_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_4QVal_Int_bufchan_r = (! lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf :
                                                        lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_r && lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_4QVal_Int_bufchan_buf <= lizzieLet12_4QNode_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_5,QTree_Int) (q1aen_destruct,Pointer_QTree_Int) > [(lizzieLet12_4QNode_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                          (_25,Pointer_QTree_Int),
                                                                                                          (lizzieLet12_4QNode_Int_5QNode_Int,Pointer_QTree_Int),
                                                                                                          (_24,Pointer_QTree_Int)] */
  logic [3:0] q1aen_destruct_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_5_d[0] && q1aen_destruct_d[0]))
      unique case (lizzieLet12_4QNode_Int_5_d[2:1])
        2'd0: q1aen_destruct_onehotd = 4'd1;
        2'd1: q1aen_destruct_onehotd = 4'd2;
        2'd2: q1aen_destruct_onehotd = 4'd4;
        2'd3: q1aen_destruct_onehotd = 4'd8;
        default: q1aen_destruct_onehotd = 4'd0;
      endcase
    else q1aen_destruct_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_5QNone_Int_d = {q1aen_destruct_d[16:1],
                                                q1aen_destruct_onehotd[0]};
  assign _25_d = {q1aen_destruct_d[16:1], q1aen_destruct_onehotd[1]};
  assign lizzieLet12_4QNode_Int_5QNode_Int_d = {q1aen_destruct_d[16:1],
                                                q1aen_destruct_onehotd[2]};
  assign _24_d = {q1aen_destruct_d[16:1], q1aen_destruct_onehotd[3]};
  assign q1aen_destruct_r = (| (q1aen_destruct_onehotd & {_24_r,
                                                          lizzieLet12_4QNode_Int_5QNode_Int_r,
                                                          _25_r,
                                                          lizzieLet12_4QNode_Int_5QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_5_r = q1aen_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_5QNone_Int_r = ((! lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_5QNone_Int_r)
        lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d <= lizzieLet12_4QNode_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet12_4QNode_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_6,QTree_Int) (q2aeo_destruct,Pointer_QTree_Int) > [(lizzieLet12_4QNode_Int_6QNone_Int,Pointer_QTree_Int),
                                                                                                          (_23,Pointer_QTree_Int),
                                                                                                          (lizzieLet12_4QNode_Int_6QNode_Int,Pointer_QTree_Int),
                                                                                                          (_22,Pointer_QTree_Int)] */
  logic [3:0] q2aeo_destruct_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_6_d[0] && q2aeo_destruct_d[0]))
      unique case (lizzieLet12_4QNode_Int_6_d[2:1])
        2'd0: q2aeo_destruct_onehotd = 4'd1;
        2'd1: q2aeo_destruct_onehotd = 4'd2;
        2'd2: q2aeo_destruct_onehotd = 4'd4;
        2'd3: q2aeo_destruct_onehotd = 4'd8;
        default: q2aeo_destruct_onehotd = 4'd0;
      endcase
    else q2aeo_destruct_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_6QNone_Int_d = {q2aeo_destruct_d[16:1],
                                                q2aeo_destruct_onehotd[0]};
  assign _23_d = {q2aeo_destruct_d[16:1], q2aeo_destruct_onehotd[1]};
  assign lizzieLet12_4QNode_Int_6QNode_Int_d = {q2aeo_destruct_d[16:1],
                                                q2aeo_destruct_onehotd[2]};
  assign _22_d = {q2aeo_destruct_d[16:1], q2aeo_destruct_onehotd[3]};
  assign q2aeo_destruct_r = (| (q2aeo_destruct_onehotd & {_22_r,
                                                          lizzieLet12_4QNode_Int_6QNode_Int_r,
                                                          _23_r,
                                                          lizzieLet12_4QNode_Int_6QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_6_r = q2aeo_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_6QNone_Int,Pointer_QTree_Int) > (lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_6QNone_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_6QNone_Int_r = ((! lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_6QNone_Int_r)
        lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d <= lizzieLet12_4QNode_Int_6QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_6QNone_Int_bufchan_r = (! lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_6QNone_Int_bufchan_buf <= lizzieLet12_4QNode_Int_6QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_7,QTree_Int) (q3aep_destruct,Pointer_QTree_Int) > [(lizzieLet12_4QNode_Int_7QNone_Int,Pointer_QTree_Int),
                                                                                                          (_21,Pointer_QTree_Int),
                                                                                                          (lizzieLet12_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                                                                                                          (_20,Pointer_QTree_Int)] */
  logic [3:0] q3aep_destruct_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_7_d[0] && q3aep_destruct_d[0]))
      unique case (lizzieLet12_4QNode_Int_7_d[2:1])
        2'd0: q3aep_destruct_onehotd = 4'd1;
        2'd1: q3aep_destruct_onehotd = 4'd2;
        2'd2: q3aep_destruct_onehotd = 4'd4;
        2'd3: q3aep_destruct_onehotd = 4'd8;
        default: q3aep_destruct_onehotd = 4'd0;
      endcase
    else q3aep_destruct_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_7QNone_Int_d = {q3aep_destruct_d[16:1],
                                                q3aep_destruct_onehotd[0]};
  assign _21_d = {q3aep_destruct_d[16:1], q3aep_destruct_onehotd[1]};
  assign lizzieLet12_4QNode_Int_7QNode_Int_d = {q3aep_destruct_d[16:1],
                                                q3aep_destruct_onehotd[2]};
  assign _20_d = {q3aep_destruct_d[16:1], q3aep_destruct_onehotd[3]};
  assign q3aep_destruct_r = (| (q3aep_destruct_onehotd & {_20_r,
                                                          lizzieLet12_4QNode_Int_7QNode_Int_r,
                                                          _21_r,
                                                          lizzieLet12_4QNode_Int_7QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_7_r = q3aep_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_7QNone_Int,Pointer_QTree_Int) > (lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_7QNone_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_7QNone_Int_r = ((! lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_7QNone_Int_r)
        lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d <= lizzieLet12_4QNode_Int_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_7QNone_Int_bufchan_r = (! lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_7QNone_Int_bufchan_buf <= lizzieLet12_4QNode_Int_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_8,QTree_Int) (q4aeq_destruct,Pointer_QTree_Int) > [(lizzieLet12_4QNode_Int_8QNone_Int,Pointer_QTree_Int),
                                                                                                          (_19,Pointer_QTree_Int),
                                                                                                          (lizzieLet12_4QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                          (_18,Pointer_QTree_Int)] */
  logic [3:0] q4aeq_destruct_onehotd;
  always_comb
    if ((lizzieLet12_4QNode_Int_8_d[0] && q4aeq_destruct_d[0]))
      unique case (lizzieLet12_4QNode_Int_8_d[2:1])
        2'd0: q4aeq_destruct_onehotd = 4'd1;
        2'd1: q4aeq_destruct_onehotd = 4'd2;
        2'd2: q4aeq_destruct_onehotd = 4'd4;
        2'd3: q4aeq_destruct_onehotd = 4'd8;
        default: q4aeq_destruct_onehotd = 4'd0;
      endcase
    else q4aeq_destruct_onehotd = 4'd0;
  assign lizzieLet12_4QNode_Int_8QNone_Int_d = {q4aeq_destruct_d[16:1],
                                                q4aeq_destruct_onehotd[0]};
  assign _19_d = {q4aeq_destruct_d[16:1], q4aeq_destruct_onehotd[1]};
  assign lizzieLet12_4QNode_Int_8QNode_Int_d = {q4aeq_destruct_d[16:1],
                                                q4aeq_destruct_onehotd[2]};
  assign _18_d = {q4aeq_destruct_d[16:1], q4aeq_destruct_onehotd[3]};
  assign q4aeq_destruct_r = (| (q4aeq_destruct_onehotd & {_18_r,
                                                          lizzieLet12_4QNode_Int_8QNode_Int_r,
                                                          _19_r,
                                                          lizzieLet12_4QNode_Int_8QNone_Int_r}));
  assign lizzieLet12_4QNode_Int_8_r = q4aeq_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_8QNode_Int,Pointer_QTree_Int) > (lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_8QNode_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_8QNode_Int_r = ((! lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_8QNode_Int_r)
        lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d <= lizzieLet12_4QNode_Int_8QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_8QNode_Int_bufchan_r = (! lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_r && lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_8QNode_Int_bufchan_buf <= lizzieLet12_4QNode_Int_8QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet12_4QNode_Int_8QNone_Int,Pointer_QTree_Int) > (lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d;
  logic lizzieLet12_4QNode_Int_8QNone_Int_bufchan_r;
  assign lizzieLet12_4QNode_Int_8QNone_Int_r = ((! lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d[0]) || lizzieLet12_4QNode_Int_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNode_Int_8QNone_Int_r)
        lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d <= lizzieLet12_4QNode_Int_8QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNode_Int_8QNone_Int_bufchan_r = (! lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_d = (lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_r && lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNode_Int_8QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNode_Int_8QNone_Int_bufchan_buf <= lizzieLet12_4QNode_Int_8QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_4QNone_Int,QTree_Int) > [(lizzieLet12_4QNone_Int_1,QTree_Int),
                                                            (lizzieLet12_4QNone_Int_2,QTree_Int),
                                                            (lizzieLet12_4QNone_Int_3,QTree_Int),
                                                            (lizzieLet12_4QNone_Int_4,QTree_Int)] */
  logic [3:0] lizzieLet12_4QNone_Int_emitted;
  logic [3:0] lizzieLet12_4QNone_Int_done;
  assign lizzieLet12_4QNone_Int_1_d = {lizzieLet12_4QNone_Int_d[66:1],
                                       (lizzieLet12_4QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_emitted[0]))};
  assign lizzieLet12_4QNone_Int_2_d = {lizzieLet12_4QNone_Int_d[66:1],
                                       (lizzieLet12_4QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_emitted[1]))};
  assign lizzieLet12_4QNone_Int_3_d = {lizzieLet12_4QNone_Int_d[66:1],
                                       (lizzieLet12_4QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_emitted[2]))};
  assign lizzieLet12_4QNone_Int_4_d = {lizzieLet12_4QNone_Int_d[66:1],
                                       (lizzieLet12_4QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_emitted[3]))};
  assign lizzieLet12_4QNone_Int_done = (lizzieLet12_4QNone_Int_emitted | ({lizzieLet12_4QNone_Int_4_d[0],
                                                                           lizzieLet12_4QNone_Int_3_d[0],
                                                                           lizzieLet12_4QNone_Int_2_d[0],
                                                                           lizzieLet12_4QNone_Int_1_d[0]} & {lizzieLet12_4QNone_Int_4_r,
                                                                                                             lizzieLet12_4QNone_Int_3_r,
                                                                                                             lizzieLet12_4QNone_Int_2_r,
                                                                                                             lizzieLet12_4QNone_Int_1_r}));
  assign lizzieLet12_4QNone_Int_r = (& lizzieLet12_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_4QNone_Int_emitted <= 4'd0;
    else
      lizzieLet12_4QNone_Int_emitted <= (lizzieLet12_4QNone_Int_r ? 4'd0 :
                                         lizzieLet12_4QNone_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet12_4QNone_Int_1QNode_Int,QTree_Int) > [(tlaea_destruct,Pointer_QTree_Int),
                                                                             (traeb_destruct,Pointer_QTree_Int),
                                                                             (blaec_destruct,Pointer_QTree_Int),
                                                                             (braed_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet12_4QNone_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet12_4QNone_Int_1QNode_Int_done;
  assign tlaea_destruct_d = {lizzieLet12_4QNone_Int_1QNode_Int_d[18:3],
                             (lizzieLet12_4QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_1QNode_Int_emitted[0]))};
  assign traeb_destruct_d = {lizzieLet12_4QNone_Int_1QNode_Int_d[34:19],
                             (lizzieLet12_4QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_1QNode_Int_emitted[1]))};
  assign blaec_destruct_d = {lizzieLet12_4QNone_Int_1QNode_Int_d[50:35],
                             (lizzieLet12_4QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_1QNode_Int_emitted[2]))};
  assign braed_destruct_d = {lizzieLet12_4QNone_Int_1QNode_Int_d[66:51],
                             (lizzieLet12_4QNone_Int_1QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet12_4QNone_Int_1QNode_Int_done = (lizzieLet12_4QNone_Int_1QNode_Int_emitted | ({braed_destruct_d[0],
                                                                                                 blaec_destruct_d[0],
                                                                                                 traeb_destruct_d[0],
                                                                                                 tlaea_destruct_d[0]} & {braed_destruct_r,
                                                                                                                         blaec_destruct_r,
                                                                                                                         traeb_destruct_r,
                                                                                                                         tlaea_destruct_r}));
  assign lizzieLet12_4QNone_Int_1QNode_Int_r = (& lizzieLet12_4QNone_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet12_4QNone_Int_1QNode_Int_emitted <= (lizzieLet12_4QNone_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet12_4QNone_Int_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_4QNone_Int_1QVal_Int,QTree_Int) > [(vae8_destruct,Int)] */
  assign vae8_destruct_d = {lizzieLet12_4QNone_Int_1QVal_Int_d[34:3],
                            lizzieLet12_4QNone_Int_1QVal_Int_d[0]};
  assign lizzieLet12_4QNone_Int_1QVal_Int_r = vae8_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_4QNone_Int_2,QTree_Int) (lizzieLet12_4QNone_Int_1,QTree_Int) > [(_17,QTree_Int),
                                                                                                    (lizzieLet12_4QNone_Int_1QVal_Int,QTree_Int),
                                                                                                    (lizzieLet12_4QNone_Int_1QNode_Int,QTree_Int),
                                                                                                    (_16,QTree_Int)] */
  logic [3:0] lizzieLet12_4QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_4QNone_Int_2_d[0] && lizzieLet12_4QNone_Int_1_d[0]))
      unique case (lizzieLet12_4QNone_Int_2_d[2:1])
        2'd0: lizzieLet12_4QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_4QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_4QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_4QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet12_4QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_4QNone_Int_1_onehotd = 4'd0;
  assign _17_d = {lizzieLet12_4QNone_Int_1_d[66:1],
                  lizzieLet12_4QNone_Int_1_onehotd[0]};
  assign lizzieLet12_4QNone_Int_1QVal_Int_d = {lizzieLet12_4QNone_Int_1_d[66:1],
                                               lizzieLet12_4QNone_Int_1_onehotd[1]};
  assign lizzieLet12_4QNone_Int_1QNode_Int_d = {lizzieLet12_4QNone_Int_1_d[66:1],
                                                lizzieLet12_4QNone_Int_1_onehotd[2]};
  assign _16_d = {lizzieLet12_4QNone_Int_1_d[66:1],
                  lizzieLet12_4QNone_Int_1_onehotd[3]};
  assign lizzieLet12_4QNone_Int_1_r = (| (lizzieLet12_4QNone_Int_1_onehotd & {_16_r,
                                                                              lizzieLet12_4QNone_Int_1QNode_Int_r,
                                                                              lizzieLet12_4QNone_Int_1QVal_Int_r,
                                                                              _17_r}));
  assign lizzieLet12_4QNone_Int_2_r = lizzieLet12_4QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_4QNone_Int_3,QTree_Int) (lizzieLet12_3QNone_Int,Go) > [(lizzieLet12_4QNone_Int_3QNone_Int,Go),
                                                                                    (lizzieLet12_4QNone_Int_3QVal_Int,Go),
                                                                                    (lizzieLet12_4QNone_Int_3QNode_Int,Go),
                                                                                    (lizzieLet12_4QNone_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QNone_Int_3_d[0] && lizzieLet12_3QNone_Int_d[0]))
      unique case (lizzieLet12_4QNone_Int_3_d[2:1])
        2'd0: lizzieLet12_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QNone_Int_onehotd = 4'd0;
  assign lizzieLet12_4QNone_Int_3QNone_Int_d = lizzieLet12_3QNone_Int_onehotd[0];
  assign lizzieLet12_4QNone_Int_3QVal_Int_d = lizzieLet12_3QNone_Int_onehotd[1];
  assign lizzieLet12_4QNone_Int_3QNode_Int_d = lizzieLet12_3QNone_Int_onehotd[2];
  assign lizzieLet12_4QNone_Int_3QError_Int_d = lizzieLet12_3QNone_Int_onehotd[3];
  assign lizzieLet12_3QNone_Int_r = (| (lizzieLet12_3QNone_Int_onehotd & {lizzieLet12_4QNone_Int_3QError_Int_r,
                                                                          lizzieLet12_4QNone_Int_3QNode_Int_r,
                                                                          lizzieLet12_4QNone_Int_3QVal_Int_r,
                                                                          lizzieLet12_4QNone_Int_3QNone_Int_r}));
  assign lizzieLet12_4QNone_Int_3_r = lizzieLet12_3QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_4QNone_Int_3QError_Int,Go) > [(lizzieLet12_4QNone_Int_3QError_Int_1,Go),
                                                          (lizzieLet12_4QNone_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QNone_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_4QNone_Int_3QError_Int_done;
  assign lizzieLet12_4QNone_Int_3QError_Int_1_d = (lizzieLet12_4QNone_Int_3QError_Int_d[0] && (! lizzieLet12_4QNone_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_4QNone_Int_3QError_Int_2_d = (lizzieLet12_4QNone_Int_3QError_Int_d[0] && (! lizzieLet12_4QNone_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_4QNone_Int_3QError_Int_done = (lizzieLet12_4QNone_Int_3QError_Int_emitted | ({lizzieLet12_4QNone_Int_3QError_Int_2_d[0],
                                                                                                   lizzieLet12_4QNone_Int_3QError_Int_1_d[0]} & {lizzieLet12_4QNone_Int_3QError_Int_2_r,
                                                                                                                                                 lizzieLet12_4QNone_Int_3QError_Int_1_r}));
  assign lizzieLet12_4QNone_Int_3QError_Int_r = (& lizzieLet12_4QNone_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QNone_Int_3QError_Int_emitted <= (lizzieLet12_4QNone_Int_3QError_Int_r ? 2'd0 :
                                                     lizzieLet12_4QNone_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_4QNone_Int_3QError_Int_1,Go)] > (lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_4QNone_Int_3QError_Int_1_d[0]}), lizzieLet12_4QNone_Int_3QError_Int_1_d);
  assign {lizzieLet12_4QNone_Int_3QError_Int_1_r} = {1 {(lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_r && lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet21_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_r = ((! lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_r)
        lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d <= lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_r = (! lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_buf <= lizzieLet12_4QNone_Int_3QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QError_Int_2,Go) > (lizzieLet12_4QNone_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QError_Int_2_r = ((! lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QError_Int_2_r)
        lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d <= lizzieLet12_4QNone_Int_3QError_Int_2_d;
  Go_t lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_d = (lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf :
                                                          lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_r && lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_4QNone_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int,Go) > [(lizzieLet12_4QNone_Int_3QNode_Int_1,Go),
                                                         (lizzieLet12_4QNone_Int_3QNode_Int_2,Go),
                                                         (lizzieLet12_4QNone_Int_3QNode_Int_3,Go),
                                                         (lizzieLet12_4QNone_Int_3QNode_Int_4,Go),
                                                         (lizzieLet12_4QNone_Int_3QNode_Int_5,Go)] */
  logic [4:0] lizzieLet12_4QNone_Int_3QNode_Int_emitted;
  logic [4:0] lizzieLet12_4QNone_Int_3QNode_Int_done;
  assign lizzieLet12_4QNone_Int_3QNode_Int_1_d = (lizzieLet12_4QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNode_Int_emitted[0]));
  assign lizzieLet12_4QNone_Int_3QNode_Int_2_d = (lizzieLet12_4QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNode_Int_emitted[1]));
  assign lizzieLet12_4QNone_Int_3QNode_Int_3_d = (lizzieLet12_4QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNode_Int_emitted[2]));
  assign lizzieLet12_4QNone_Int_3QNode_Int_4_d = (lizzieLet12_4QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNode_Int_emitted[3]));
  assign lizzieLet12_4QNone_Int_3QNode_Int_5_d = (lizzieLet12_4QNone_Int_3QNode_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNode_Int_emitted[4]));
  assign lizzieLet12_4QNone_Int_3QNode_Int_done = (lizzieLet12_4QNone_Int_3QNode_Int_emitted | ({lizzieLet12_4QNone_Int_3QNode_Int_5_d[0],
                                                                                                 lizzieLet12_4QNone_Int_3QNode_Int_4_d[0],
                                                                                                 lizzieLet12_4QNone_Int_3QNode_Int_3_d[0],
                                                                                                 lizzieLet12_4QNone_Int_3QNode_Int_2_d[0],
                                                                                                 lizzieLet12_4QNone_Int_3QNode_Int_1_d[0]} & {lizzieLet12_4QNone_Int_3QNode_Int_5_r,
                                                                                                                                              lizzieLet12_4QNone_Int_3QNode_Int_4_r,
                                                                                                                                              lizzieLet12_4QNone_Int_3QNode_Int_3_r,
                                                                                                                                              lizzieLet12_4QNone_Int_3QNode_Int_2_r,
                                                                                                                                              lizzieLet12_4QNone_Int_3QNode_Int_1_r}));
  assign lizzieLet12_4QNone_Int_3QNode_Int_r = (& lizzieLet12_4QNone_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_emitted <= 5'd0;
    else
      lizzieLet12_4QNone_Int_3QNode_Int_emitted <= (lizzieLet12_4QNone_Int_3QNode_Int_r ? 5'd0 :
                                                    lizzieLet12_4QNone_Int_3QNode_Int_done);
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int_1,Go) > (lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNode_Int_1_r = ((! lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNode_Int_1_r)
        lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d <= lizzieLet12_4QNone_Int_3QNode_Int_1_d;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_r = (! lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_d = (lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_r && lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_buf <= lizzieLet12_4QNone_Int_3QNode_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf,Go),
                                         (braed_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_d[0],
                                                                                               braed_1_argbuf_d[0]}), lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_d, braed_1_argbuf_d);
  assign {lizzieLet12_4QNone_Int_3QNode_Int_1_argbuf_r,
          braed_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int_2,Go) > (lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNode_Int_2_r = ((! lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNode_Int_2_r)
        lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d <= lizzieLet12_4QNone_Int_3QNode_Int_2_d;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_r = (! lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_d = (lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_r && lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_buf <= lizzieLet12_4QNone_Int_3QNode_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf,Go),
                                         (blaec_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int2,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_d[0],
                                                                                              blaec_1_argbuf_d[0]}), lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_d, blaec_1_argbuf_d);
  assign {lizzieLet12_4QNone_Int_3QNode_Int_2_argbuf_r,
          blaec_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int2_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int_3,Go) > (lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNode_Int_3_r = ((! lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNode_Int_3_r)
        lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d <= lizzieLet12_4QNone_Int_3QNode_Int_3_d;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_r = (! lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_d = (lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_r && lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_buf <= lizzieLet12_4QNone_Int_3QNode_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf,Go),
                                         (traeb_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int3,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_d[0],
                                                                                              traeb_1_argbuf_d[0]}), lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_d, traeb_1_argbuf_d);
  assign {lizzieLet12_4QNone_Int_3QNode_Int_3_argbuf_r,
          traeb_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int3_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int_4,Go) > (lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNode_Int_4_r = ((! lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNode_Int_4_r)
        lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d <= lizzieLet12_4QNone_Int_3QNode_Int_4_d;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_r = (! lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_d = (lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_r && lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_buf <= lizzieLet12_4QNone_Int_3QNode_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf,Go),
                                         (tlaea_1_argbuf,Pointer_QTree_Int)] > (f''''''''_f''''''''TupGo___Pointer_QTree_Int4,TupGo___Pointer_QTree_Int) */
  assign \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_d  = TupGo___Pointer_QTree_Int_dc((& {lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_d[0],
                                                                                              tlaea_1_argbuf_d[0]}), lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_d, tlaea_1_argbuf_d);
  assign {lizzieLet12_4QNone_Int_3QNode_Int_4_argbuf_r,
          tlaea_1_argbuf_r} = {2 {(\f''''''''_f''''''''TupGo___Pointer_QTree_Int4_r  && \f''''''''_f''''''''TupGo___Pointer_QTree_Int4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNode_Int_5,Go) > (lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNode_Int_5_r = ((! lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNode_Int_5_r)
        lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d <= lizzieLet12_4QNone_Int_3QNode_Int_5_d;
  Go_t lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_r = (! lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_d = (lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_r && lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_buf <= lizzieLet12_4QNone_Int_3QNode_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_4QNone_Int_3QNone_Int,Go) > [(lizzieLet12_4QNone_Int_3QNone_Int_1,Go),
                                                         (lizzieLet12_4QNone_Int_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QNone_Int_3QNone_Int_emitted;
  logic [1:0] lizzieLet12_4QNone_Int_3QNone_Int_done;
  assign lizzieLet12_4QNone_Int_3QNone_Int_1_d = (lizzieLet12_4QNone_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNone_Int_emitted[0]));
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_d = (lizzieLet12_4QNone_Int_3QNone_Int_d[0] && (! lizzieLet12_4QNone_Int_3QNone_Int_emitted[1]));
  assign lizzieLet12_4QNone_Int_3QNone_Int_done = (lizzieLet12_4QNone_Int_3QNone_Int_emitted | ({lizzieLet12_4QNone_Int_3QNone_Int_2_d[0],
                                                                                                 lizzieLet12_4QNone_Int_3QNone_Int_1_d[0]} & {lizzieLet12_4QNone_Int_3QNone_Int_2_r,
                                                                                                                                              lizzieLet12_4QNone_Int_3QNone_Int_1_r}));
  assign lizzieLet12_4QNone_Int_3QNone_Int_r = (& lizzieLet12_4QNone_Int_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QNone_Int_3QNone_Int_emitted <= (lizzieLet12_4QNone_Int_3QNone_Int_r ? 2'd0 :
                                                    lizzieLet12_4QNone_Int_3QNone_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet12_4QNone_Int_3QNone_Int_1,Go)] > (lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool,QTree_Bool) */
  assign lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet12_4QNone_Int_3QNone_Int_1_d[0]}), lizzieLet12_4QNone_Int_3QNone_Int_1_d);
  assign {lizzieLet12_4QNone_Int_3QNone_Int_1_r} = {1 {(lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_r && lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool,QTree_Bool) > (lizzieLet14_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_r = ((! lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_r)
        lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d <= lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_d;
  QTree_Bool_t lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_r = (! lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf :
                                   lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_buf <= lizzieLet12_4QNone_Int_3QNone_Int_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QNone_Int_3QNone_Int_2,Go) > (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d;
  logic lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_r;
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_r = ((! lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d[0]) || lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QNone_Int_3QNone_Int_2_r)
        lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d <= lizzieLet12_4QNone_Int_3QNone_Int_2_d;
  Go_t lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf;
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_r = (! lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_d = (lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf[0] ? lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_r && lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_r) && (! lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_buf <= lizzieLet12_4QNone_Int_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C16,
           Ty Go) : [(lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf,Go),
                     (lizzieLet53_3Lcall_f_f0_1_argbuf,Go),
                     (lizzieLet17_1MyFalse_2_argbuf,Go),
                     (lizzieLet17_1MyTrue_2_argbuf,Go),
                     (lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf,Go),
                     (lizzieLet12_4QNone_Int_3QError_Int_2_argbuf,Go),
                     (lizzieLet25_1MyFalse_2_argbuf,Go),
                     (lizzieLet25_1MyTrue_2_argbuf,Go),
                     (lizzieLet30_1MyFalse_2_argbuf,Go),
                     (lizzieLet30_1MyTrue_2_argbuf,Go),
                     (lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf,Go),
                     (lizzieLet12_4QVal_Int_3QError_Int_2_argbuf,Go),
                     (lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf,Go),
                     (lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf,Go),
                     (lizzieLet12_4QNode_Int_3QError_Int_2_argbuf,Go),
                     (lizzieLet12_3QError_Int_2_argbuf,Go)] > (go_21_goMux_choice,C16) (go_21_goMux_data,Go) */
  logic [15:0] lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d = ((| lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_q) ? lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_q :
                                                                (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_d[0] ? 16'd1 :
                                                                 (lizzieLet53_3Lcall_f_f0_1_argbuf_d[0] ? 16'd2 :
                                                                  (lizzieLet17_1MyFalse_2_argbuf_d[0] ? 16'd4 :
                                                                   (lizzieLet17_1MyTrue_2_argbuf_d[0] ? 16'd8 :
                                                                    (lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_d[0] ? 16'd16 :
                                                                     (lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_d[0] ? 16'd32 :
                                                                      (lizzieLet25_1MyFalse_2_argbuf_d[0] ? 16'd64 :
                                                                       (lizzieLet25_1MyTrue_2_argbuf_d[0] ? 16'd128 :
                                                                        (lizzieLet30_1MyFalse_2_argbuf_d[0] ? 16'd256 :
                                                                         (lizzieLet30_1MyTrue_2_argbuf_d[0] ? 16'd512 :
                                                                          (lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_d[0] ? 16'd1024 :
                                                                           (lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_d[0] ? 16'd2048 :
                                                                            (lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_d[0] ? 16'd4096 :
                                                                             (lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_d[0] ? 16'd8192 :
                                                                              (lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_d[0] ? 16'd16384 :
                                                                               (lizzieLet12_3QError_Int_2_argbuf_d[0] ? 16'd32768 :
                                                                                16'd0)))))))))))))))));
  logic [15:0] lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_q <= 16'd0;
    else
      lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_q <= (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_done ? 16'd0 :
                                                              lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q <= (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                            lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_d = (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q | ({go_21_goMux_choice_d[0],
                                                                                                                    go_21_goMux_data_d[0]} & {go_21_goMux_choice_r,
                                                                                                                                              go_21_goMux_data_r}));
  logic lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_done;
  assign lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_done = (& lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet12_3QError_Int_2_argbuf_r,
          lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_r,
          lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_r,
          lizzieLet30_1MyTrue_2_argbuf_r,
          lizzieLet30_1MyFalse_2_argbuf_r,
          lizzieLet25_1MyTrue_2_argbuf_r,
          lizzieLet25_1MyFalse_2_argbuf_r,
          lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_r,
          lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_r,
          lizzieLet17_1MyTrue_2_argbuf_r,
          lizzieLet17_1MyFalse_2_argbuf_r,
          lizzieLet53_3Lcall_f_f0_1_argbuf_r,
          lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_r} = (lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_done ? lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d :
                                                           16'd0);
  assign go_21_goMux_data_d = ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_d :
                               ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet53_3Lcall_f_f0_1_argbuf_d :
                                ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_1MyFalse_2_argbuf_d :
                                 ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_1MyTrue_2_argbuf_d :
                                  ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNone_Int_3QNode_Int_5_argbuf_d :
                                   ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[5] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNone_Int_3QError_Int_2_argbuf_d :
                                    ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[6] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet25_1MyFalse_2_argbuf_d :
                                     ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[7] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet25_1MyTrue_2_argbuf_d :
                                      ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[8] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet30_1MyFalse_2_argbuf_d :
                                       ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[9] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet30_1MyTrue_2_argbuf_d :
                                        ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[10] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_d :
                                         ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[11] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_d :
                                          ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[12] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNode_Int_3QNone_Int_5_argbuf_d :
                                           ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[13] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNode_Int_3QVal_Int_2_argbuf_d :
                                            ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[14] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_4QNode_Int_3QError_Int_2_argbuf_d :
                                             ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[15] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet12_3QError_Int_2_argbuf_d :
                                              1'd0))))))))))))))));
  assign go_21_goMux_choice_d = ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C1_16_dc(1'd1) :
                                 ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C2_16_dc(1'd1) :
                                  ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C3_16_dc(1'd1) :
                                   ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C4_16_dc(1'd1) :
                                    ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C5_16_dc(1'd1) :
                                     ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[5] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C6_16_dc(1'd1) :
                                      ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[6] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C7_16_dc(1'd1) :
                                       ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[7] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C8_16_dc(1'd1) :
                                        ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[8] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C9_16_dc(1'd1) :
                                         ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[9] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C10_16_dc(1'd1) :
                                          ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[10] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C11_16_dc(1'd1) :
                                           ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[11] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C12_16_dc(1'd1) :
                                            ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[12] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C13_16_dc(1'd1) :
                                             ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[13] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C14_16_dc(1'd1) :
                                              ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[14] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C15_16_dc(1'd1) :
                                               ((lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_select_d[15] && (! lizzieLet12_4QNone_Int_3QNone_Int_2_argbuf_emit_q[1])) ? C16_16_dc(1'd1) :
                                                {4'd0, 1'd0}))))))))))))))));
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QNone_Int_4,QTree_Int) (lizzieLet12_5QNone_Int,Pointer_CTf_f) > [(lizzieLet12_4QNone_Int_4QNone_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNone_Int_4QVal_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNone_Int_4QNode_Int,Pointer_CTf_f),
                                                                                                          (lizzieLet12_4QNone_Int_4QError_Int,Pointer_CTf_f)] */
  logic [3:0] lizzieLet12_5QNone_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QNone_Int_4_d[0] && lizzieLet12_5QNone_Int_d[0]))
      unique case (lizzieLet12_4QNone_Int_4_d[2:1])
        2'd0: lizzieLet12_5QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QNone_Int_onehotd = 4'd8;
        default: lizzieLet12_5QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QNone_Int_onehotd = 4'd0;
  assign lizzieLet12_4QNone_Int_4QNone_Int_d = {lizzieLet12_5QNone_Int_d[16:1],
                                                lizzieLet12_5QNone_Int_onehotd[0]};
  assign lizzieLet12_4QNone_Int_4QVal_Int_d = {lizzieLet12_5QNone_Int_d[16:1],
                                               lizzieLet12_5QNone_Int_onehotd[1]};
  assign lizzieLet12_4QNone_Int_4QNode_Int_d = {lizzieLet12_5QNone_Int_d[16:1],
                                                lizzieLet12_5QNone_Int_onehotd[2]};
  assign lizzieLet12_4QNone_Int_4QError_Int_d = {lizzieLet12_5QNone_Int_d[16:1],
                                                 lizzieLet12_5QNone_Int_onehotd[3]};
  assign lizzieLet12_5QNone_Int_r = (| (lizzieLet12_5QNone_Int_onehotd & {lizzieLet12_4QNone_Int_4QError_Int_r,
                                                                          lizzieLet12_4QNone_Int_4QNode_Int_r,
                                                                          lizzieLet12_4QNone_Int_4QVal_Int_r,
                                                                          lizzieLet12_4QNone_Int_4QNone_Int_r}));
  assign lizzieLet12_4QNone_Int_4_r = lizzieLet12_5QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNone_Int_4QError_Int,Pointer_CTf_f) > (lizzieLet12_4QNone_Int_4QError_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QError_Int_bufchan_d;
  logic lizzieLet12_4QNone_Int_4QError_Int_bufchan_r;
  assign lizzieLet12_4QNone_Int_4QError_Int_r = ((! lizzieLet12_4QNone_Int_4QError_Int_bufchan_d[0]) || lizzieLet12_4QNone_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNone_Int_4QError_Int_r)
        lizzieLet12_4QNone_Int_4QError_Int_bufchan_d <= lizzieLet12_4QNone_Int_4QError_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf;
  assign lizzieLet12_4QNone_Int_4QError_Int_bufchan_r = (! lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_d = (lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf[0] ? lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf :
                                                          lizzieLet12_4QNone_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_r && lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNone_Int_4QError_Int_1_argbuf_r) && (! lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_4QError_Int_bufchan_buf <= lizzieLet12_4QNone_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNone_Int_4QNode_Int,Pointer_CTf_f) > (lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d;
  logic lizzieLet12_4QNone_Int_4QNode_Int_bufchan_r;
  assign lizzieLet12_4QNone_Int_4QNode_Int_r = ((! lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d[0]) || lizzieLet12_4QNone_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNone_Int_4QNode_Int_r)
        lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d <= lizzieLet12_4QNone_Int_4QNode_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet12_4QNone_Int_4QNode_Int_bufchan_r = (! lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_d = (lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_r && lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNone_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_4QNode_Int_bufchan_buf <= lizzieLet12_4QNone_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QNone_Int_4QNone_Int,Pointer_CTf_f) > (lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d;
  logic lizzieLet12_4QNone_Int_4QNone_Int_bufchan_r;
  assign lizzieLet12_4QNone_Int_4QNone_Int_r = ((! lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d[0]) || lizzieLet12_4QNone_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QNone_Int_4QNone_Int_r)
        lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d <= lizzieLet12_4QNone_Int_4QNone_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet12_4QNone_Int_4QNone_Int_bufchan_r = (! lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_d = (lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf :
                                                         lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_r && lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QNone_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet12_4QNone_Int_4QNone_Int_bufchan_buf <= lizzieLet12_4QNone_Int_4QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet12_4QVal_Int,QTree_Int) > [(lizzieLet12_4QVal_Int_1,QTree_Int),
                                                           (lizzieLet12_4QVal_Int_2,QTree_Int),
                                                           (lizzieLet12_4QVal_Int_3,QTree_Int),
                                                           (lizzieLet12_4QVal_Int_4,QTree_Int),
                                                           (lizzieLet12_4QVal_Int_5,QTree_Int)] */
  logic [4:0] lizzieLet12_4QVal_Int_emitted;
  logic [4:0] lizzieLet12_4QVal_Int_done;
  assign lizzieLet12_4QVal_Int_1_d = {lizzieLet12_4QVal_Int_d[66:1],
                                      (lizzieLet12_4QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_emitted[0]))};
  assign lizzieLet12_4QVal_Int_2_d = {lizzieLet12_4QVal_Int_d[66:1],
                                      (lizzieLet12_4QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_emitted[1]))};
  assign lizzieLet12_4QVal_Int_3_d = {lizzieLet12_4QVal_Int_d[66:1],
                                      (lizzieLet12_4QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_emitted[2]))};
  assign lizzieLet12_4QVal_Int_4_d = {lizzieLet12_4QVal_Int_d[66:1],
                                      (lizzieLet12_4QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_emitted[3]))};
  assign lizzieLet12_4QVal_Int_5_d = {lizzieLet12_4QVal_Int_d[66:1],
                                      (lizzieLet12_4QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_emitted[4]))};
  assign lizzieLet12_4QVal_Int_done = (lizzieLet12_4QVal_Int_emitted | ({lizzieLet12_4QVal_Int_5_d[0],
                                                                         lizzieLet12_4QVal_Int_4_d[0],
                                                                         lizzieLet12_4QVal_Int_3_d[0],
                                                                         lizzieLet12_4QVal_Int_2_d[0],
                                                                         lizzieLet12_4QVal_Int_1_d[0]} & {lizzieLet12_4QVal_Int_5_r,
                                                                                                          lizzieLet12_4QVal_Int_4_r,
                                                                                                          lizzieLet12_4QVal_Int_3_r,
                                                                                                          lizzieLet12_4QVal_Int_2_r,
                                                                                                          lizzieLet12_4QVal_Int_1_r}));
  assign lizzieLet12_4QVal_Int_r = (& lizzieLet12_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_4QVal_Int_emitted <= 5'd0;
    else
      lizzieLet12_4QVal_Int_emitted <= (lizzieLet12_4QVal_Int_r ? 5'd0 :
                                        lizzieLet12_4QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet12_4QVal_Int_1QVal_Int,QTree_Int) > [(vaeg_destruct,Int)] */
  assign vaeg_destruct_d = {lizzieLet12_4QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet12_4QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet12_4QVal_Int_1QVal_Int_r = vaeg_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet12_4QVal_Int_2,QTree_Int) (lizzieLet12_4QVal_Int_1,QTree_Int) > [(_15,QTree_Int),
                                                                                                  (lizzieLet12_4QVal_Int_1QVal_Int,QTree_Int),
                                                                                                  (_14,QTree_Int),
                                                                                                  (_13,QTree_Int)] */
  logic [3:0] lizzieLet12_4QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet12_4QVal_Int_2_d[0] && lizzieLet12_4QVal_Int_1_d[0]))
      unique case (lizzieLet12_4QVal_Int_2_d[2:1])
        2'd0: lizzieLet12_4QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet12_4QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet12_4QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet12_4QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet12_4QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_4QVal_Int_1_onehotd = 4'd0;
  assign _15_d = {lizzieLet12_4QVal_Int_1_d[66:1],
                  lizzieLet12_4QVal_Int_1_onehotd[0]};
  assign lizzieLet12_4QVal_Int_1QVal_Int_d = {lizzieLet12_4QVal_Int_1_d[66:1],
                                              lizzieLet12_4QVal_Int_1_onehotd[1]};
  assign _14_d = {lizzieLet12_4QVal_Int_1_d[66:1],
                  lizzieLet12_4QVal_Int_1_onehotd[2]};
  assign _13_d = {lizzieLet12_4QVal_Int_1_d[66:1],
                  lizzieLet12_4QVal_Int_1_onehotd[3]};
  assign lizzieLet12_4QVal_Int_1_r = (| (lizzieLet12_4QVal_Int_1_onehotd & {_13_r,
                                                                            _14_r,
                                                                            lizzieLet12_4QVal_Int_1QVal_Int_r,
                                                                            _15_r}));
  assign lizzieLet12_4QVal_Int_2_r = lizzieLet12_4QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet12_4QVal_Int_3,QTree_Int) (lizzieLet12_3QVal_Int,Go) > [(lizzieLet12_4QVal_Int_3QNone_Int,Go),
                                                                                  (lizzieLet12_4QVal_Int_3QVal_Int,Go),
                                                                                  (lizzieLet12_4QVal_Int_3QNode_Int,Go),
                                                                                  (lizzieLet12_4QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet12_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QVal_Int_3_d[0] && lizzieLet12_3QVal_Int_d[0]))
      unique case (lizzieLet12_4QVal_Int_3_d[2:1])
        2'd0: lizzieLet12_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_4QVal_Int_3QNone_Int_d = lizzieLet12_3QVal_Int_onehotd[0];
  assign lizzieLet12_4QVal_Int_3QVal_Int_d = lizzieLet12_3QVal_Int_onehotd[1];
  assign lizzieLet12_4QVal_Int_3QNode_Int_d = lizzieLet12_3QVal_Int_onehotd[2];
  assign lizzieLet12_4QVal_Int_3QError_Int_d = lizzieLet12_3QVal_Int_onehotd[3];
  assign lizzieLet12_3QVal_Int_r = (| (lizzieLet12_3QVal_Int_onehotd & {lizzieLet12_4QVal_Int_3QError_Int_r,
                                                                        lizzieLet12_4QVal_Int_3QNode_Int_r,
                                                                        lizzieLet12_4QVal_Int_3QVal_Int_r,
                                                                        lizzieLet12_4QVal_Int_3QNone_Int_r}));
  assign lizzieLet12_4QVal_Int_3_r = lizzieLet12_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet12_4QVal_Int_3QError_Int,Go) > [(lizzieLet12_4QVal_Int_3QError_Int_1,Go),
                                                         (lizzieLet12_4QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet12_4QVal_Int_3QError_Int_done;
  assign lizzieLet12_4QVal_Int_3QError_Int_1_d = (lizzieLet12_4QVal_Int_3QError_Int_d[0] && (! lizzieLet12_4QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet12_4QVal_Int_3QError_Int_2_d = (lizzieLet12_4QVal_Int_3QError_Int_d[0] && (! lizzieLet12_4QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet12_4QVal_Int_3QError_Int_done = (lizzieLet12_4QVal_Int_3QError_Int_emitted | ({lizzieLet12_4QVal_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet12_4QVal_Int_3QError_Int_1_d[0]} & {lizzieLet12_4QVal_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet12_4QVal_Int_3QError_Int_1_r}));
  assign lizzieLet12_4QVal_Int_3QError_Int_r = (& lizzieLet12_4QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QVal_Int_3QError_Int_emitted <= (lizzieLet12_4QVal_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet12_4QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_4QVal_Int_3QError_Int_1,Go)] > (lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_4QVal_Int_3QError_Int_1_d[0]}), lizzieLet12_4QVal_Int_3QError_Int_1_d);
  assign {lizzieLet12_4QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_r && lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet34_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_r = ((! lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_r)
        lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d <= lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_r = (! lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_buf <= lizzieLet12_4QVal_Int_3QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_3QError_Int_2,Go) > (lizzieLet12_4QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet12_4QVal_Int_3QError_Int_2_r = ((! lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QVal_Int_3QError_Int_2_r)
        lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet12_4QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_r && lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet12_4QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_4QVal_Int_3QNode_Int,Go) > [(lizzieLet12_4QVal_Int_3QNode_Int_1,Go),
                                                        (lizzieLet12_4QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet12_4QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet12_4QVal_Int_3QNode_Int_done;
  assign lizzieLet12_4QVal_Int_3QNode_Int_1_d = (lizzieLet12_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet12_4QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet12_4QVal_Int_3QNode_Int_2_d = (lizzieLet12_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet12_4QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet12_4QVal_Int_3QNode_Int_done = (lizzieLet12_4QVal_Int_3QNode_Int_emitted | ({lizzieLet12_4QVal_Int_3QNode_Int_2_d[0],
                                                                                               lizzieLet12_4QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet12_4QVal_Int_3QNode_Int_2_r,
                                                                                                                                           lizzieLet12_4QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet12_4QVal_Int_3QNode_Int_r = (& lizzieLet12_4QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet12_4QVal_Int_3QNode_Int_emitted <= (lizzieLet12_4QVal_Int_3QNode_Int_r ? 2'd0 :
                                                   lizzieLet12_4QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_4QVal_Int_3QNode_Int_1,Go)] > (lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_4QVal_Int_3QNode_Int_1_d[0]}), lizzieLet12_4QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet12_4QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_r && lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool,QTree_Bool) > (lizzieLet33_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_r;
  assign lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_r = ((! lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d[0]) || lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_r)
        lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d <= lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_r = (! lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_buf <= lizzieLet12_4QVal_Int_3QNode_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_3QNode_Int_2,Go) > (lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet12_4QVal_Int_3QNode_Int_2_r = ((! lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_4QVal_Int_3QNode_Int_2_r)
        lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet12_4QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf :
                                                        lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_4QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet12_4QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_4,QTree_Int) (lizzieLet12_5QVal_Int,Pointer_CTf_f) > [(lizzieLet12_4QVal_Int_4QNone_Int,Pointer_CTf_f),
                                                                                                        (lizzieLet12_4QVal_Int_4QVal_Int,Pointer_CTf_f),
                                                                                                        (lizzieLet12_4QVal_Int_4QNode_Int,Pointer_CTf_f),
                                                                                                        (lizzieLet12_4QVal_Int_4QError_Int,Pointer_CTf_f)] */
  logic [3:0] lizzieLet12_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet12_4QVal_Int_4_d[0] && lizzieLet12_5QVal_Int_d[0]))
      unique case (lizzieLet12_4QVal_Int_4_d[2:1])
        2'd0: lizzieLet12_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet12_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet12_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet12_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet12_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet12_5QVal_Int_onehotd = 4'd0;
  assign lizzieLet12_4QVal_Int_4QNone_Int_d = {lizzieLet12_5QVal_Int_d[16:1],
                                               lizzieLet12_5QVal_Int_onehotd[0]};
  assign lizzieLet12_4QVal_Int_4QVal_Int_d = {lizzieLet12_5QVal_Int_d[16:1],
                                              lizzieLet12_5QVal_Int_onehotd[1]};
  assign lizzieLet12_4QVal_Int_4QNode_Int_d = {lizzieLet12_5QVal_Int_d[16:1],
                                               lizzieLet12_5QVal_Int_onehotd[2]};
  assign lizzieLet12_4QVal_Int_4QError_Int_d = {lizzieLet12_5QVal_Int_d[16:1],
                                                lizzieLet12_5QVal_Int_onehotd[3]};
  assign lizzieLet12_5QVal_Int_r = (| (lizzieLet12_5QVal_Int_onehotd & {lizzieLet12_4QVal_Int_4QError_Int_r,
                                                                        lizzieLet12_4QVal_Int_4QNode_Int_r,
                                                                        lizzieLet12_4QVal_Int_4QVal_Int_r,
                                                                        lizzieLet12_4QVal_Int_4QNone_Int_r}));
  assign lizzieLet12_4QVal_Int_4_r = lizzieLet12_5QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_4QError_Int,Pointer_CTf_f) > (lizzieLet12_4QVal_Int_4QError_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QError_Int_bufchan_d;
  logic lizzieLet12_4QVal_Int_4QError_Int_bufchan_r;
  assign lizzieLet12_4QVal_Int_4QError_Int_r = ((! lizzieLet12_4QVal_Int_4QError_Int_bufchan_d[0]) || lizzieLet12_4QVal_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QVal_Int_4QError_Int_r)
        lizzieLet12_4QVal_Int_4QError_Int_bufchan_d <= lizzieLet12_4QVal_Int_4QError_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf;
  assign lizzieLet12_4QVal_Int_4QError_Int_bufchan_r = (! lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_d = (lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf[0] ? lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf :
                                                         lizzieLet12_4QVal_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_r && lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QVal_Int_4QError_Int_1_argbuf_r) && (! lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_4QError_Int_bufchan_buf <= lizzieLet12_4QVal_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_4QNode_Int,Pointer_CTf_f) > (lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d;
  logic lizzieLet12_4QVal_Int_4QNode_Int_bufchan_r;
  assign lizzieLet12_4QVal_Int_4QNode_Int_r = ((! lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d[0]) || lizzieLet12_4QVal_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_4QVal_Int_4QNode_Int_r)
        lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d <= lizzieLet12_4QVal_Int_4QNode_Int_d;
  Pointer_CTf_f_t lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet12_4QVal_Int_4QNode_Int_bufchan_r = (! lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_d = (lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf :
                                                        lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_r && lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_4QVal_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet12_4QVal_Int_4QNode_Int_bufchan_buf <= lizzieLet12_4QVal_Int_4QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet12_4QVal_Int_5,QTree_Int) (v1aee_destruct,Int) > [(lizzieLet12_4QVal_Int_5QNone_Int,Int),
                                                                             (lizzieLet12_4QVal_Int_5QVal_Int,Int),
                                                                             (_12,Int),
                                                                             (_11,Int)] */
  logic [3:0] v1aee_destruct_onehotd;
  always_comb
    if ((lizzieLet12_4QVal_Int_5_d[0] && v1aee_destruct_d[0]))
      unique case (lizzieLet12_4QVal_Int_5_d[2:1])
        2'd0: v1aee_destruct_onehotd = 4'd1;
        2'd1: v1aee_destruct_onehotd = 4'd2;
        2'd2: v1aee_destruct_onehotd = 4'd4;
        2'd3: v1aee_destruct_onehotd = 4'd8;
        default: v1aee_destruct_onehotd = 4'd0;
      endcase
    else v1aee_destruct_onehotd = 4'd0;
  assign lizzieLet12_4QVal_Int_5QNone_Int_d = {v1aee_destruct_d[32:1],
                                               v1aee_destruct_onehotd[0]};
  assign lizzieLet12_4QVal_Int_5QVal_Int_d = {v1aee_destruct_d[32:1],
                                              v1aee_destruct_onehotd[1]};
  assign _12_d = {v1aee_destruct_d[32:1], v1aee_destruct_onehotd[2]};
  assign _11_d = {v1aee_destruct_d[32:1], v1aee_destruct_onehotd[3]};
  assign v1aee_destruct_r = (| (v1aee_destruct_onehotd & {_11_r,
                                                          _12_r,
                                                          lizzieLet12_4QVal_Int_5QVal_Int_r,
                                                          lizzieLet12_4QVal_Int_5QNone_Int_r}));
  assign lizzieLet12_4QVal_Int_5_r = v1aee_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet12_4QVal_Int_5QNone_Int,Int) > [(lizzieLet12_4QVal_Int_5QNone_Int_1,Int),
                                                          (lizzieLet12_4QVal_Int_5QNone_Int_2,Int),
                                                          (lizzieLet12_4QVal_Int_5QNone_Int_3,Int),
                                                          (lizzieLet12_4QVal_Int_5QNone_Int_4,Int)] */
  logic [3:0] lizzieLet12_4QVal_Int_5QNone_Int_emitted;
  logic [3:0] lizzieLet12_4QVal_Int_5QNone_Int_done;
  assign lizzieLet12_4QVal_Int_5QNone_Int_1_d = {lizzieLet12_4QVal_Int_5QNone_Int_d[32:1],
                                                 (lizzieLet12_4QVal_Int_5QNone_Int_d[0] && (! lizzieLet12_4QVal_Int_5QNone_Int_emitted[0]))};
  assign lizzieLet12_4QVal_Int_5QNone_Int_2_d = {lizzieLet12_4QVal_Int_5QNone_Int_d[32:1],
                                                 (lizzieLet12_4QVal_Int_5QNone_Int_d[0] && (! lizzieLet12_4QVal_Int_5QNone_Int_emitted[1]))};
  assign lizzieLet12_4QVal_Int_5QNone_Int_3_d = {lizzieLet12_4QVal_Int_5QNone_Int_d[32:1],
                                                 (lizzieLet12_4QVal_Int_5QNone_Int_d[0] && (! lizzieLet12_4QVal_Int_5QNone_Int_emitted[2]))};
  assign lizzieLet12_4QVal_Int_5QNone_Int_4_d = {lizzieLet12_4QVal_Int_5QNone_Int_d[32:1],
                                                 (lizzieLet12_4QVal_Int_5QNone_Int_d[0] && (! lizzieLet12_4QVal_Int_5QNone_Int_emitted[3]))};
  assign lizzieLet12_4QVal_Int_5QNone_Int_done = (lizzieLet12_4QVal_Int_5QNone_Int_emitted | ({lizzieLet12_4QVal_Int_5QNone_Int_4_d[0],
                                                                                               lizzieLet12_4QVal_Int_5QNone_Int_3_d[0],
                                                                                               lizzieLet12_4QVal_Int_5QNone_Int_2_d[0],
                                                                                               lizzieLet12_4QVal_Int_5QNone_Int_1_d[0]} & {lizzieLet12_4QVal_Int_5QNone_Int_4_r,
                                                                                                                                           lizzieLet12_4QVal_Int_5QNone_Int_3_r,
                                                                                                                                           lizzieLet12_4QVal_Int_5QNone_Int_2_r,
                                                                                                                                           lizzieLet12_4QVal_Int_5QNone_Int_1_r}));
  assign lizzieLet12_4QVal_Int_5QNone_Int_r = (& lizzieLet12_4QVal_Int_5QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_5QNone_Int_emitted <= 4'd0;
    else
      lizzieLet12_4QVal_Int_5QNone_Int_emitted <= (lizzieLet12_4QVal_Int_5QNone_Int_r ? 4'd0 :
                                                   lizzieLet12_4QVal_Int_5QNone_Int_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (lizzieLet12_4QVal_Int_5QNone_Int_1I#,Int) > [(xakK_2_destruct,Int#)] */
  assign xakK_2_destruct_d = {\lizzieLet12_4QVal_Int_5QNone_Int_1I#_d [32:1],
                              \lizzieLet12_4QVal_Int_5QNone_Int_1I#_d [0]};
  assign \lizzieLet12_4QVal_Int_5QNone_Int_1I#_r  = xakK_2_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (lizzieLet12_4QVal_Int_5QNone_Int_2,Int) (lizzieLet12_4QVal_Int_5QNone_Int_1,Int) > [(lizzieLet12_4QVal_Int_5QNone_Int_1I#,Int)] */
  assign \lizzieLet12_4QVal_Int_5QNone_Int_1I#_d  = {lizzieLet12_4QVal_Int_5QNone_Int_1_d[32:1],
                                                     (lizzieLet12_4QVal_Int_5QNone_Int_2_d[0] && lizzieLet12_4QVal_Int_5QNone_Int_1_d[0])};
  assign lizzieLet12_4QVal_Int_5QNone_Int_1_r = (\lizzieLet12_4QVal_Int_5QNone_Int_1I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_2_d[0] && lizzieLet12_4QVal_Int_5QNone_Int_1_d[0]));
  assign lizzieLet12_4QVal_Int_5QNone_Int_2_r = (\lizzieLet12_4QVal_Int_5QNone_Int_1I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_2_d[0] && lizzieLet12_4QVal_Int_5QNone_Int_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (lizzieLet12_4QVal_Int_5QNone_Int_3,Int) (lizzieLet12_4QVal_Int_3QNone_Int,Go) > [(lizzieLet12_4QVal_Int_5QNone_Int_3I#,Go)] */
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_d  = (lizzieLet12_4QVal_Int_5QNone_Int_3_d[0] && lizzieLet12_4QVal_Int_3QNone_Int_d[0]);
  assign lizzieLet12_4QVal_Int_3QNone_Int_r = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_3_d[0] && lizzieLet12_4QVal_Int_3QNone_Int_d[0]));
  assign lizzieLet12_4QVal_Int_5QNone_Int_3_r = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_3_d[0] && lizzieLet12_4QVal_Int_3QNone_Int_d[0]));
  
  /* fork (Ty Go) : (lizzieLet12_4QVal_Int_5QNone_Int_3I#,Go) > [(lizzieLet12_4QVal_Int_5QNone_Int_3I#_1,Go),
                                                            (lizzieLet12_4QVal_Int_5QNone_Int_3I#_2,Go),
                                                            (lizzieLet12_4QVal_Int_5QNone_Int_3I#_3,Go)] */
  logic [2:0] \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted ;
  logic [2:0] \lizzieLet12_4QVal_Int_5QNone_Int_3I#_done ;
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_d  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted [0]));
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_d  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted [1]));
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_d  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted [2]));
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_done  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted  | ({\lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_d [0],
                                                                                                           \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_d [0],
                                                                                                           \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_d [0]} & {\lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_r ,
                                                                                                                                                             \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_r ,
                                                                                                                                                             \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_r }));
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_r  = (& \lizzieLet12_4QVal_Int_5QNone_Int_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted  <= 3'd0;
    else
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_emitted  <= (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_r  ? 3'd0 :
                                                         \lizzieLet12_4QVal_Int_5QNone_Int_3I#_done );
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_5QNone_Int_3I#_1,Go) > (lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf,Go) */
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_r ;
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_r  = ((! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d [0]) || \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_r )
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d  <= \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_d ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf ;
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_r  = (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf [0]);
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_d  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf [0] ? \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf  :
                                                              \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_r  && \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf [0]))
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_r ) && (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf [0])))
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_buf  <= \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf,Go) > (lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0,Int#) */
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_d  = {32'd0,
                                                                \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_d [0]};
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_r  = \lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0,Int#) (xakK_2_destruct,Int#) > (lizzieLet23_1wild3XR_1_1_Eq,Bool) */
  assign lizzieLet23_1wild3XR_1_1_Eq_d = {(\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_d [32:1] == xakK_2_destruct_d[32:1]),
                                          (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_d [0] && xakK_2_destruct_d[0])};
  assign {\lizzieLet12_4QVal_Int_5QNone_Int_3I#_1_argbuf_0_r ,
          xakK_2_destruct_r} = {2 {(lizzieLet23_1wild3XR_1_1_Eq_r && lizzieLet23_1wild3XR_1_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_5QNone_Int_3I#_2,Go) > (lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf,Go) */
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d ;
  logic \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_r ;
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_r  = ((! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d [0]) || \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_r )
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d  <= \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_d ;
  Go_t \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf ;
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_r  = (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf [0]);
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_d  = (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf [0] ? \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf  :
                                                              \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_r  && \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf [0]))
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_r ) && (! \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf [0])))
        \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_buf  <= \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf,Go),
                            (lizzieLet24_1_argbuf,Bool)] > (boolConvert_3TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_3TupGo___Bool_1_d = TupGo___Bool_dc((& {\lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_d [0],
                                                             lizzieLet24_1_argbuf_d[0]}), \lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_d , lizzieLet24_1_argbuf_d);
  assign {\lizzieLet12_4QVal_Int_5QNone_Int_3I#_2_argbuf_r ,
          lizzieLet24_1_argbuf_r} = {2 {(boolConvert_3TupGo___Bool_1_r && boolConvert_3TupGo___Bool_1_d[0])}};
  
  /* demux (Ty Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_5QNone_Int_4,Int) (lizzieLet12_4QVal_Int_4QNone_Int,Pointer_CTf_f) > [(lizzieLet12_4QVal_Int_5QNone_Int_4I#,Pointer_CTf_f)] */
  assign \lizzieLet12_4QVal_Int_5QNone_Int_4I#_d  = {lizzieLet12_4QVal_Int_4QNone_Int_d[16:1],
                                                     (lizzieLet12_4QVal_Int_5QNone_Int_4_d[0] && lizzieLet12_4QVal_Int_4QNone_Int_d[0])};
  assign lizzieLet12_4QVal_Int_4QNone_Int_r = (\lizzieLet12_4QVal_Int_5QNone_Int_4I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_4_d[0] && lizzieLet12_4QVal_Int_4QNone_Int_d[0]));
  assign lizzieLet12_4QVal_Int_5QNone_Int_4_r = (\lizzieLet12_4QVal_Int_5QNone_Int_4I#_r  && (lizzieLet12_4QVal_Int_5QNone_Int_4_d[0] && lizzieLet12_4QVal_Int_4QNone_Int_d[0]));
  
  /* fork (Ty Int) : (lizzieLet12_4QVal_Int_5QVal_Int,Int) > [(lizzieLet12_4QVal_Int_5QVal_Int_1,Int),
                                                         (lizzieLet12_4QVal_Int_5QVal_Int_2,Int),
                                                         (lizzieLet12_4QVal_Int_5QVal_Int_3,Int),
                                                         (lizzieLet12_4QVal_Int_5QVal_Int_4,Int),
                                                         (lizzieLet12_4QVal_Int_5QVal_Int_5,Int)] */
  logic [4:0] lizzieLet12_4QVal_Int_5QVal_Int_emitted;
  logic [4:0] lizzieLet12_4QVal_Int_5QVal_Int_done;
  assign lizzieLet12_4QVal_Int_5QVal_Int_1_d = {lizzieLet12_4QVal_Int_5QVal_Int_d[32:1],
                                                (lizzieLet12_4QVal_Int_5QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_5QVal_Int_emitted[0]))};
  assign lizzieLet12_4QVal_Int_5QVal_Int_2_d = {lizzieLet12_4QVal_Int_5QVal_Int_d[32:1],
                                                (lizzieLet12_4QVal_Int_5QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_5QVal_Int_emitted[1]))};
  assign lizzieLet12_4QVal_Int_5QVal_Int_3_d = {lizzieLet12_4QVal_Int_5QVal_Int_d[32:1],
                                                (lizzieLet12_4QVal_Int_5QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_5QVal_Int_emitted[2]))};
  assign lizzieLet12_4QVal_Int_5QVal_Int_4_d = {lizzieLet12_4QVal_Int_5QVal_Int_d[32:1],
                                                (lizzieLet12_4QVal_Int_5QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_5QVal_Int_emitted[3]))};
  assign lizzieLet12_4QVal_Int_5QVal_Int_5_d = {lizzieLet12_4QVal_Int_5QVal_Int_d[32:1],
                                                (lizzieLet12_4QVal_Int_5QVal_Int_d[0] && (! lizzieLet12_4QVal_Int_5QVal_Int_emitted[4]))};
  assign lizzieLet12_4QVal_Int_5QVal_Int_done = (lizzieLet12_4QVal_Int_5QVal_Int_emitted | ({lizzieLet12_4QVal_Int_5QVal_Int_5_d[0],
                                                                                             lizzieLet12_4QVal_Int_5QVal_Int_4_d[0],
                                                                                             lizzieLet12_4QVal_Int_5QVal_Int_3_d[0],
                                                                                             lizzieLet12_4QVal_Int_5QVal_Int_2_d[0],
                                                                                             lizzieLet12_4QVal_Int_5QVal_Int_1_d[0]} & {lizzieLet12_4QVal_Int_5QVal_Int_5_r,
                                                                                                                                        lizzieLet12_4QVal_Int_5QVal_Int_4_r,
                                                                                                                                        lizzieLet12_4QVal_Int_5QVal_Int_3_r,
                                                                                                                                        lizzieLet12_4QVal_Int_5QVal_Int_2_r,
                                                                                                                                        lizzieLet12_4QVal_Int_5QVal_Int_1_r}));
  assign lizzieLet12_4QVal_Int_5QVal_Int_r = (& lizzieLet12_4QVal_Int_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_4QVal_Int_5QVal_Int_emitted <= 5'd0;
    else
      lizzieLet12_4QVal_Int_5QVal_Int_emitted <= (lizzieLet12_4QVal_Int_5QVal_Int_r ? 5'd0 :
                                                  lizzieLet12_4QVal_Int_5QVal_Int_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (lizzieLet12_4QVal_Int_5QVal_Int_1I#,Int) > [(xakw_destruct,Int#)] */
  assign xakw_destruct_d = {\lizzieLet12_4QVal_Int_5QVal_Int_1I#_d [32:1],
                            \lizzieLet12_4QVal_Int_5QVal_Int_1I#_d [0]};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_1I#_r  = xakw_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (lizzieLet12_4QVal_Int_5QVal_Int_2,Int) (lizzieLet12_4QVal_Int_5QVal_Int_1,Int) > [(lizzieLet12_4QVal_Int_5QVal_Int_1I#,Int)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_1I#_d  = {lizzieLet12_4QVal_Int_5QVal_Int_1_d[32:1],
                                                    (lizzieLet12_4QVal_Int_5QVal_Int_2_d[0] && lizzieLet12_4QVal_Int_5QVal_Int_1_d[0])};
  assign lizzieLet12_4QVal_Int_5QVal_Int_1_r = (\lizzieLet12_4QVal_Int_5QVal_Int_1I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_2_d[0] && lizzieLet12_4QVal_Int_5QVal_Int_1_d[0]));
  assign lizzieLet12_4QVal_Int_5QVal_Int_2_r = (\lizzieLet12_4QVal_Int_5QVal_Int_1I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_2_d[0] && lizzieLet12_4QVal_Int_5QVal_Int_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (lizzieLet12_4QVal_Int_5QVal_Int_3,Int) (lizzieLet12_4QVal_Int_3QVal_Int,Go) > [(lizzieLet12_4QVal_Int_5QVal_Int_3I#,Go)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_3I#_d  = (lizzieLet12_4QVal_Int_5QVal_Int_3_d[0] && lizzieLet12_4QVal_Int_3QVal_Int_d[0]);
  assign lizzieLet12_4QVal_Int_3QVal_Int_r = (\lizzieLet12_4QVal_Int_5QVal_Int_3I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_3_d[0] && lizzieLet12_4QVal_Int_3QVal_Int_d[0]));
  assign lizzieLet12_4QVal_Int_5QVal_Int_3_r = (\lizzieLet12_4QVal_Int_5QVal_Int_3I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_3_d[0] && lizzieLet12_4QVal_Int_3QVal_Int_d[0]));
  
  /* demux (Ty Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_5QVal_Int_4,Int) (lizzieLet12_4QVal_Int_4QVal_Int,Pointer_CTf_f) > [(lizzieLet12_4QVal_Int_5QVal_Int_4I#,Pointer_CTf_f)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_4I#_d  = {lizzieLet12_4QVal_Int_4QVal_Int_d[16:1],
                                                    (lizzieLet12_4QVal_Int_5QVal_Int_4_d[0] && lizzieLet12_4QVal_Int_4QVal_Int_d[0])};
  assign lizzieLet12_4QVal_Int_4QVal_Int_r = (\lizzieLet12_4QVal_Int_5QVal_Int_4I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_4_d[0] && lizzieLet12_4QVal_Int_4QVal_Int_d[0]));
  assign lizzieLet12_4QVal_Int_5QVal_Int_4_r = (\lizzieLet12_4QVal_Int_5QVal_Int_4I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_4_d[0] && lizzieLet12_4QVal_Int_4QVal_Int_d[0]));
  
  /* demux (Ty Int,
       Ty Int) : (lizzieLet12_4QVal_Int_5QVal_Int_5,Int) (vaeg_destruct,Int) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#,Int)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_d  = {vaeg_destruct_d[32:1],
                                                    (lizzieLet12_4QVal_Int_5QVal_Int_5_d[0] && vaeg_destruct_d[0])};
  assign vaeg_destruct_r = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_5_d[0] && vaeg_destruct_d[0]));
  assign lizzieLet12_4QVal_Int_5QVal_Int_5_r = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_r  && (lizzieLet12_4QVal_Int_5QVal_Int_5_d[0] && vaeg_destruct_d[0]));
  
  /* fork (Ty Int) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#,Int) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_1,Int),
                                                             (lizzieLet12_4QVal_Int_5QVal_Int_5I#_2,Int),
                                                             (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3,Int),
                                                             (lizzieLet12_4QVal_Int_5QVal_Int_5I#_4,Int),
                                                             (lizzieLet12_4QVal_Int_5QVal_Int_5I#_5,Int)] */
  logic [4:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted ;
  logic [4:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_done ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [32:1],
                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted [0]))};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [32:1],
                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted [1]))};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [32:1],
                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted [2]))};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [32:1],
                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted [3]))};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [32:1],
                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted [4]))};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_done  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted  | ({\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d [0],
                                                                                                         \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d [0],
                                                                                                         \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d [0],
                                                                                                         \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d [0],
                                                                                                         \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d [0]} & {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_r ,
                                                                                                                                                          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_r ,
                                                                                                                                                          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_r ,
                                                                                                                                                          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_r ,
                                                                                                                                                          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_r }));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_r  = (& \lizzieLet12_4QVal_Int_5QVal_Int_5I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted  <= 5'd0;
    else
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_emitted  <= (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_r  ? 5'd0 :
                                                        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#,Int) > [(yakA_destruct,Int#)] */
  assign yakA_destruct_d = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_d [32:1],
                            \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_d [0]};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_r  = yakA_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_2,Int) (lizzieLet12_4QVal_Int_5QVal_Int_5I#_1,Int) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#,Int)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d [32:1],
                                                        (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d [0])};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d [0]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_1I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_2_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Go) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3,Int) (lizzieLet12_4QVal_Int_5QVal_Int_3I#,Go) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#,Go)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_3I#_d [0]);
  assign \lizzieLet12_4QVal_Int_5QVal_Int_3I#_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_3I#_d [0]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_3I#_d [0]));
  
  /* fork (Ty Go) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#,Go) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1,Go),
                                                               (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2,Go),
                                                               (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3,Go)] */
  logic [2:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted ;
  logic [2:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_done ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted [0]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted [1]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_d [0] && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted [2]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_done  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted  | ({\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_d [0],
                                                                                                                 \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_d [0],
                                                                                                                 \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_d [0]} & {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_r ,
                                                                                                                                                                      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_r ,
                                                                                                                                                                      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_r }));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_r  = (& \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted  <= 3'd0;
    else
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_emitted  <= (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_r  ? 3'd0 :
                                                            \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_done );
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1,Go) > (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf,Go) */
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_r ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_r  = ((! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d [0]) || \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_r )
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d  <= \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_d ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_r  = (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf [0]);
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf [0] ? \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf  :
                                                                 \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_r  && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf [0]))
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_r ) && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf [0])))
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_buf  <= \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf,Go) > (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0,Int#) */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_d  = {32'd0,
                                                                   \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_d [0]};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_r  = \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0,Int#) (lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32,Int#) > (lizzieLet28_1wild4XU_1_Eq,Bool) */
  assign lizzieLet28_1wild4XU_1_Eq_d = {(\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_d [32:1] == \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_d [32:1]),
                                        (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_d [0])};
  assign {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_1_argbuf_0_r ,
          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_r } = {2 {(lizzieLet28_1wild4XU_1_Eq_r && lizzieLet28_1wild4XU_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2,Go) > (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf,Go) */
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d ;
  logic \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_r ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_r  = ((! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d [0]) || \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_r )
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d  <= \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_d ;
  Go_t \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf ;
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_r  = (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf [0]);
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_d  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf [0] ? \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf  :
                                                                 \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_r  && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf [0]))
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_r ) && (! \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf [0])))
        \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_buf  <= \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf,Go),
                            (lizzieLet29_1_argbuf,Bool)] > (boolConvert_4TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_4TupGo___Bool_1_d = TupGo___Bool_dc((& {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_d [0],
                                                             lizzieLet29_1_argbuf_d[0]}), \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_d , lizzieLet29_1_argbuf_d);
  assign {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_2_argbuf_r ,
          lizzieLet29_1_argbuf_r} = {2 {(boolConvert_4TupGo___Bool_1_r && boolConvert_4TupGo___Bool_1_d[0])}};
  
  /* demux (Ty Int,
       Ty Pointer_CTf_f) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_4,Int) (lizzieLet12_4QVal_Int_5QVal_Int_4I#,Pointer_CTf_f) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#,Pointer_CTf_f)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_d  = {\lizzieLet12_4QVal_Int_5QVal_Int_4I#_d [16:1],
                                                        (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_4I#_d [0])};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_4I#_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_4I#_d [0]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4_d [0] && \lizzieLet12_4QVal_Int_5QVal_Int_4I#_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_5,Int) (xakw_destruct,Int#) > [(lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#,Int#)] */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_d  = {xakw_destruct_d[32:1],
                                                        (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d [0] && xakw_destruct_d[0])};
  assign xakw_destruct_r = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d [0] && xakw_destruct_d[0]));
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_r  = (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_r  && (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5_d [0] && xakw_destruct_d[0]));
  
  /* op_add (Ty Int#) : (lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#,Int#) (yakA_destruct,Int#) > (lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32,Int#) */
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_d  = {(\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_d [32:1] + yakA_destruct_d[32:1]),
                                                                      (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_d [0] && yakA_destruct_d[0])};
  assign {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_r ,
          yakA_destruct_r} = {2 {(\lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_r  && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_5I#_1yakA_1_Add32_d [0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f) : (lizzieLet12_5,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTf_f) > [(lizzieLet12_5QNone_Int,Pointer_CTf_f),
                                                                                         (lizzieLet12_5QVal_Int,Pointer_CTf_f),
                                                                                         (lizzieLet12_5QNode_Int,Pointer_CTf_f),
                                                                                         (lizzieLet12_5QError_Int,Pointer_CTf_f)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_5_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet12_5_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_5QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet12_5QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet12_5QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet12_5QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet12_5QError_Int_r,
                                                              lizzieLet12_5QNode_Int_r,
                                                              lizzieLet12_5QVal_Int_r,
                                                              lizzieLet12_5QNone_Int_r}));
  assign lizzieLet12_5_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet12_5QError_Int,Pointer_CTf_f) > (lizzieLet12_5QError_Int_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet12_5QError_Int_bufchan_d;
  logic lizzieLet12_5QError_Int_bufchan_r;
  assign lizzieLet12_5QError_Int_r = ((! lizzieLet12_5QError_Int_bufchan_d[0]) || lizzieLet12_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_5QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_5QError_Int_r)
        lizzieLet12_5QError_Int_bufchan_d <= lizzieLet12_5QError_Int_d;
  Pointer_CTf_f_t lizzieLet12_5QError_Int_bufchan_buf;
  assign lizzieLet12_5QError_Int_bufchan_r = (! lizzieLet12_5QError_Int_bufchan_buf[0]);
  assign lizzieLet12_5QError_Int_1_argbuf_d = (lizzieLet12_5QError_Int_bufchan_buf[0] ? lizzieLet12_5QError_Int_bufchan_buf :
                                               lizzieLet12_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_5QError_Int_1_argbuf_r && lizzieLet12_5QError_Int_bufchan_buf[0]))
        lizzieLet12_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_5QError_Int_1_argbuf_r) && (! lizzieLet12_5QError_Int_bufchan_buf[0])))
        lizzieLet12_5QError_Int_bufchan_buf <= lizzieLet12_5QError_Int_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet15_1wild3XR_1_Eq,Bool) > (lizzieLet16_1_argbuf,Bool) */
  Bool_t lizzieLet15_1wild3XR_1_Eq_bufchan_d;
  logic lizzieLet15_1wild3XR_1_Eq_bufchan_r;
  assign lizzieLet15_1wild3XR_1_Eq_r = ((! lizzieLet15_1wild3XR_1_Eq_bufchan_d[0]) || lizzieLet15_1wild3XR_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_1wild3XR_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet15_1wild3XR_1_Eq_r)
        lizzieLet15_1wild3XR_1_Eq_bufchan_d <= lizzieLet15_1wild3XR_1_Eq_d;
  Bool_t lizzieLet15_1wild3XR_1_Eq_bufchan_buf;
  assign lizzieLet15_1wild3XR_1_Eq_bufchan_r = (! lizzieLet15_1wild3XR_1_Eq_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet15_1wild3XR_1_Eq_bufchan_buf[0] ? lizzieLet15_1wild3XR_1_Eq_bufchan_buf :
                                   lizzieLet15_1wild3XR_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_1wild3XR_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet15_1wild3XR_1_Eq_bufchan_buf[0]))
        lizzieLet15_1wild3XR_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet15_1wild3XR_1_Eq_bufchan_buf[0])))
        lizzieLet15_1wild3XR_1_Eq_bufchan_buf <= lizzieLet15_1wild3XR_1_Eq_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet17_1,MyBool) (vae8_3I#_3,Go) > [(lizzieLet17_1MyFalse,Go),
                                                          (lizzieLet17_1MyTrue,Go)] */
  logic [1:0] \vae8_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet17_1_d[0] && \vae8_3I#_3_d [0]))
      unique case (lizzieLet17_1_d[1:1])
        1'd0: \vae8_3I#_3_onehotd  = 2'd1;
        1'd1: \vae8_3I#_3_onehotd  = 2'd2;
        default: \vae8_3I#_3_onehotd  = 2'd0;
      endcase
    else \vae8_3I#_3_onehotd  = 2'd0;
  assign lizzieLet17_1MyFalse_d = \vae8_3I#_3_onehotd [0];
  assign lizzieLet17_1MyTrue_d = \vae8_3I#_3_onehotd [1];
  assign \vae8_3I#_3_r  = (| (\vae8_3I#_3_onehotd  & {lizzieLet17_1MyTrue_r,
                                                      lizzieLet17_1MyFalse_r}));
  assign lizzieLet17_1_r = \vae8_3I#_3_r ;
  
  /* fork (Ty Go) : (lizzieLet17_1MyFalse,Go) > [(lizzieLet17_1MyFalse_1,Go),
                                            (lizzieLet17_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet17_1MyFalse_emitted;
  logic [1:0] lizzieLet17_1MyFalse_done;
  assign lizzieLet17_1MyFalse_1_d = (lizzieLet17_1MyFalse_d[0] && (! lizzieLet17_1MyFalse_emitted[0]));
  assign lizzieLet17_1MyFalse_2_d = (lizzieLet17_1MyFalse_d[0] && (! lizzieLet17_1MyFalse_emitted[1]));
  assign lizzieLet17_1MyFalse_done = (lizzieLet17_1MyFalse_emitted | ({lizzieLet17_1MyFalse_2_d[0],
                                                                       lizzieLet17_1MyFalse_1_d[0]} & {lizzieLet17_1MyFalse_2_r,
                                                                                                       lizzieLet17_1MyFalse_1_r}));
  assign lizzieLet17_1MyFalse_r = (& lizzieLet17_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet17_1MyFalse_emitted <= (lizzieLet17_1MyFalse_r ? 2'd0 :
                                       lizzieLet17_1MyFalse_done);
  
  /* buf (Ty Go) : (lizzieLet17_1MyFalse_1,Go) > (lizzieLet17_1MyFalse_1_argbuf,Go) */
  Go_t lizzieLet17_1MyFalse_1_bufchan_d;
  logic lizzieLet17_1MyFalse_1_bufchan_r;
  assign lizzieLet17_1MyFalse_1_r = ((! lizzieLet17_1MyFalse_1_bufchan_d[0]) || lizzieLet17_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_1MyFalse_1_r)
        lizzieLet17_1MyFalse_1_bufchan_d <= lizzieLet17_1MyFalse_1_d;
  Go_t lizzieLet17_1MyFalse_1_bufchan_buf;
  assign lizzieLet17_1MyFalse_1_bufchan_r = (! lizzieLet17_1MyFalse_1_bufchan_buf[0]);
  assign lizzieLet17_1MyFalse_1_argbuf_d = (lizzieLet17_1MyFalse_1_bufchan_buf[0] ? lizzieLet17_1MyFalse_1_bufchan_buf :
                                            lizzieLet17_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_1MyFalse_1_argbuf_r && lizzieLet17_1MyFalse_1_bufchan_buf[0]))
        lizzieLet17_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_1MyFalse_1_argbuf_r) && (! lizzieLet17_1MyFalse_1_bufchan_buf[0])))
        lizzieLet17_1MyFalse_1_bufchan_buf <= lizzieLet17_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet17_1MyFalse_1_argbuf,Go)] > (f''''''''1TupGo_1,TupGo) */
  assign \f''''''''1TupGo_1_d  = TupGo_dc((& {lizzieLet17_1MyFalse_1_argbuf_d[0]}), lizzieLet17_1MyFalse_1_argbuf_d);
  assign {lizzieLet17_1MyFalse_1_argbuf_r} = {1 {(\f''''''''1TupGo_1_r  && \f''''''''1TupGo_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet17_1MyFalse_2,Go) > (lizzieLet17_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet17_1MyFalse_2_bufchan_d;
  logic lizzieLet17_1MyFalse_2_bufchan_r;
  assign lizzieLet17_1MyFalse_2_r = ((! lizzieLet17_1MyFalse_2_bufchan_d[0]) || lizzieLet17_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_1MyFalse_2_r)
        lizzieLet17_1MyFalse_2_bufchan_d <= lizzieLet17_1MyFalse_2_d;
  Go_t lizzieLet17_1MyFalse_2_bufchan_buf;
  assign lizzieLet17_1MyFalse_2_bufchan_r = (! lizzieLet17_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet17_1MyFalse_2_argbuf_d = (lizzieLet17_1MyFalse_2_bufchan_buf[0] ? lizzieLet17_1MyFalse_2_bufchan_buf :
                                            lizzieLet17_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_1MyFalse_2_argbuf_r && lizzieLet17_1MyFalse_2_bufchan_buf[0]))
        lizzieLet17_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_1MyFalse_2_argbuf_r) && (! lizzieLet17_1MyFalse_2_bufchan_buf[0])))
        lizzieLet17_1MyFalse_2_bufchan_buf <= lizzieLet17_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_1MyTrue,Go) > [(lizzieLet17_1MyTrue_1,Go),
                                           (lizzieLet17_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet17_1MyTrue_emitted;
  logic [1:0] lizzieLet17_1MyTrue_done;
  assign lizzieLet17_1MyTrue_1_d = (lizzieLet17_1MyTrue_d[0] && (! lizzieLet17_1MyTrue_emitted[0]));
  assign lizzieLet17_1MyTrue_2_d = (lizzieLet17_1MyTrue_d[0] && (! lizzieLet17_1MyTrue_emitted[1]));
  assign lizzieLet17_1MyTrue_done = (lizzieLet17_1MyTrue_emitted | ({lizzieLet17_1MyTrue_2_d[0],
                                                                     lizzieLet17_1MyTrue_1_d[0]} & {lizzieLet17_1MyTrue_2_r,
                                                                                                    lizzieLet17_1MyTrue_1_r}));
  assign lizzieLet17_1MyTrue_r = (& lizzieLet17_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet17_1MyTrue_emitted <= (lizzieLet17_1MyTrue_r ? 2'd0 :
                                      lizzieLet17_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet17_1MyTrue_1,Go)] > (lizzieLet17_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign lizzieLet17_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet17_1MyTrue_1_d[0]}), lizzieLet17_1MyTrue_1_d);
  assign {lizzieLet17_1MyTrue_1_r} = {1 {(lizzieLet17_1MyTrue_1QNone_Bool_r && lizzieLet17_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet17_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet19_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d;
  logic lizzieLet17_1MyTrue_1QNone_Bool_bufchan_r;
  assign lizzieLet17_1MyTrue_1QNone_Bool_r = ((! lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d[0]) || lizzieLet17_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_1MyTrue_1QNone_Bool_r)
        lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d <= lizzieLet17_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf;
  assign lizzieLet17_1MyTrue_1QNone_Bool_bufchan_r = (! lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet19_1_1_argbuf_d = (lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf[0] ? lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf :
                                     lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet19_1_1_argbuf_r && lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet19_1_1_argbuf_r) && (! lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        lizzieLet17_1MyTrue_1QNone_Bool_bufchan_buf <= lizzieLet17_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_1MyTrue_2,Go) > (lizzieLet17_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet17_1MyTrue_2_bufchan_d;
  logic lizzieLet17_1MyTrue_2_bufchan_r;
  assign lizzieLet17_1MyTrue_2_r = ((! lizzieLet17_1MyTrue_2_bufchan_d[0]) || lizzieLet17_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_1MyTrue_2_r)
        lizzieLet17_1MyTrue_2_bufchan_d <= lizzieLet17_1MyTrue_2_d;
  Go_t lizzieLet17_1MyTrue_2_bufchan_buf;
  assign lizzieLet17_1MyTrue_2_bufchan_r = (! lizzieLet17_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet17_1MyTrue_2_argbuf_d = (lizzieLet17_1MyTrue_2_bufchan_buf[0] ? lizzieLet17_1MyTrue_2_bufchan_buf :
                                           lizzieLet17_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_1MyTrue_2_argbuf_r && lizzieLet17_1MyTrue_2_bufchan_buf[0]))
        lizzieLet17_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_1MyTrue_2_argbuf_r) && (! lizzieLet17_1MyTrue_2_bufchan_buf[0])))
        lizzieLet17_1MyTrue_2_bufchan_buf <= lizzieLet17_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f) : (lizzieLet17_2,MyBool) (vae8_4I#,Pointer_CTf_f) > [(lizzieLet17_2MyFalse,Pointer_CTf_f),
                                                                              (lizzieLet17_2MyTrue,Pointer_CTf_f)] */
  logic [1:0] \vae8_4I#_onehotd ;
  always_comb
    if ((lizzieLet17_2_d[0] && \vae8_4I#_d [0]))
      unique case (lizzieLet17_2_d[1:1])
        1'd0: \vae8_4I#_onehotd  = 2'd1;
        1'd1: \vae8_4I#_onehotd  = 2'd2;
        default: \vae8_4I#_onehotd  = 2'd0;
      endcase
    else \vae8_4I#_onehotd  = 2'd0;
  assign lizzieLet17_2MyFalse_d = {\vae8_4I#_d [16:1],
                                   \vae8_4I#_onehotd [0]};
  assign lizzieLet17_2MyTrue_d = {\vae8_4I#_d [16:1],
                                  \vae8_4I#_onehotd [1]};
  assign \vae8_4I#_r  = (| (\vae8_4I#_onehotd  & {lizzieLet17_2MyTrue_r,
                                                  lizzieLet17_2MyFalse_r}));
  assign lizzieLet17_2_r = \vae8_4I#_r ;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet17_2MyFalse,Pointer_CTf_f) > (lizzieLet17_2MyFalse_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet17_2MyFalse_bufchan_d;
  logic lizzieLet17_2MyFalse_bufchan_r;
  assign lizzieLet17_2MyFalse_r = ((! lizzieLet17_2MyFalse_bufchan_d[0]) || lizzieLet17_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_2MyFalse_r)
        lizzieLet17_2MyFalse_bufchan_d <= lizzieLet17_2MyFalse_d;
  Pointer_CTf_f_t lizzieLet17_2MyFalse_bufchan_buf;
  assign lizzieLet17_2MyFalse_bufchan_r = (! lizzieLet17_2MyFalse_bufchan_buf[0]);
  assign lizzieLet17_2MyFalse_1_argbuf_d = (lizzieLet17_2MyFalse_bufchan_buf[0] ? lizzieLet17_2MyFalse_bufchan_buf :
                                            lizzieLet17_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_2MyFalse_1_argbuf_r && lizzieLet17_2MyFalse_bufchan_buf[0]))
        lizzieLet17_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_2MyFalse_1_argbuf_r) && (! lizzieLet17_2MyFalse_bufchan_buf[0])))
        lizzieLet17_2MyFalse_bufchan_buf <= lizzieLet17_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet17_2MyTrue,Pointer_CTf_f) > (lizzieLet17_2MyTrue_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet17_2MyTrue_bufchan_d;
  logic lizzieLet17_2MyTrue_bufchan_r;
  assign lizzieLet17_2MyTrue_r = ((! lizzieLet17_2MyTrue_bufchan_d[0]) || lizzieLet17_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_2MyTrue_r)
        lizzieLet17_2MyTrue_bufchan_d <= lizzieLet17_2MyTrue_d;
  Pointer_CTf_f_t lizzieLet17_2MyTrue_bufchan_buf;
  assign lizzieLet17_2MyTrue_bufchan_r = (! lizzieLet17_2MyTrue_bufchan_buf[0]);
  assign lizzieLet17_2MyTrue_1_argbuf_d = (lizzieLet17_2MyTrue_bufchan_buf[0] ? lizzieLet17_2MyTrue_bufchan_buf :
                                           lizzieLet17_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_2MyTrue_1_argbuf_r && lizzieLet17_2MyTrue_bufchan_buf[0]))
        lizzieLet17_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_2MyTrue_1_argbuf_r) && (! lizzieLet17_2MyTrue_bufchan_buf[0])))
        lizzieLet17_2MyTrue_bufchan_buf <= lizzieLet17_2MyTrue_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet1_1QNode_Bool,QTree_Bool) > [(q1a84_destruct,Pointer_QTree_Bool),
                                                                    (q2a85_destruct,Pointer_QTree_Bool),
                                                                    (q3a86_destruct,Pointer_QTree_Bool),
                                                                    (q4a87_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet1_1QNode_Bool_emitted;
  logic [3:0] lizzieLet1_1QNode_Bool_done;
  assign q1a84_destruct_d = {lizzieLet1_1QNode_Bool_d[18:3],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[0]))};
  assign q2a85_destruct_d = {lizzieLet1_1QNode_Bool_d[34:19],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[1]))};
  assign q3a86_destruct_d = {lizzieLet1_1QNode_Bool_d[50:35],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[2]))};
  assign q4a87_destruct_d = {lizzieLet1_1QNode_Bool_d[66:51],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[3]))};
  assign lizzieLet1_1QNode_Bool_done = (lizzieLet1_1QNode_Bool_emitted | ({q4a87_destruct_d[0],
                                                                           q3a86_destruct_d[0],
                                                                           q2a85_destruct_d[0],
                                                                           q1a84_destruct_d[0]} & {q4a87_destruct_r,
                                                                                                   q3a86_destruct_r,
                                                                                                   q2a85_destruct_r,
                                                                                                   q1a84_destruct_r}));
  assign lizzieLet1_1QNode_Bool_r = (& lizzieLet1_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet1_1QNode_Bool_emitted <= (lizzieLet1_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet1_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet1_2,QTree_Bool) (lizzieLet1_1,QTree_Bool) > [(_10,QTree_Bool),
                                                                               (_9,QTree_Bool),
                                                                               (lizzieLet1_1QNode_Bool,QTree_Bool),
                                                                               (_8,QTree_Bool)] */
  logic [3:0] lizzieLet1_1_onehotd;
  always_comb
    if ((lizzieLet1_2_d[0] && lizzieLet1_1_d[0]))
      unique case (lizzieLet1_2_d[2:1])
        2'd0: lizzieLet1_1_onehotd = 4'd1;
        2'd1: lizzieLet1_1_onehotd = 4'd2;
        2'd2: lizzieLet1_1_onehotd = 4'd4;
        2'd3: lizzieLet1_1_onehotd = 4'd8;
        default: lizzieLet1_1_onehotd = 4'd0;
      endcase
    else lizzieLet1_1_onehotd = 4'd0;
  assign _10_d = {lizzieLet1_1_d[66:1], lizzieLet1_1_onehotd[0]};
  assign _9_d = {lizzieLet1_1_d[66:1], lizzieLet1_1_onehotd[1]};
  assign lizzieLet1_1QNode_Bool_d = {lizzieLet1_1_d[66:1],
                                     lizzieLet1_1_onehotd[2]};
  assign _8_d = {lizzieLet1_1_d[66:1], lizzieLet1_1_onehotd[3]};
  assign lizzieLet1_1_r = (| (lizzieLet1_1_onehotd & {_8_r,
                                                      lizzieLet1_1QNode_Bool_r,
                                                      _9_r,
                                                      _10_r}));
  assign lizzieLet1_2_r = lizzieLet1_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet1_3,QTree_Bool) (go_13_goMux_data,Go) > [(lizzieLet1_3QNone_Bool,Go),
                                                                   (lizzieLet1_3QVal_Bool,Go),
                                                                   (lizzieLet1_3QNode_Bool,Go),
                                                                   (lizzieLet1_3QError_Bool,Go)] */
  logic [3:0] go_13_goMux_data_onehotd;
  always_comb
    if ((lizzieLet1_3_d[0] && go_13_goMux_data_d[0]))
      unique case (lizzieLet1_3_d[2:1])
        2'd0: go_13_goMux_data_onehotd = 4'd1;
        2'd1: go_13_goMux_data_onehotd = 4'd2;
        2'd2: go_13_goMux_data_onehotd = 4'd4;
        2'd3: go_13_goMux_data_onehotd = 4'd8;
        default: go_13_goMux_data_onehotd = 4'd0;
      endcase
    else go_13_goMux_data_onehotd = 4'd0;
  assign lizzieLet1_3QNone_Bool_d = go_13_goMux_data_onehotd[0];
  assign lizzieLet1_3QVal_Bool_d = go_13_goMux_data_onehotd[1];
  assign lizzieLet1_3QNode_Bool_d = go_13_goMux_data_onehotd[2];
  assign lizzieLet1_3QError_Bool_d = go_13_goMux_data_onehotd[3];
  assign go_13_goMux_data_r = (| (go_13_goMux_data_onehotd & {lizzieLet1_3QError_Bool_r,
                                                              lizzieLet1_3QNode_Bool_r,
                                                              lizzieLet1_3QVal_Bool_r,
                                                              lizzieLet1_3QNone_Bool_r}));
  assign lizzieLet1_3_r = go_13_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet1_3QError_Bool,Go) > [(lizzieLet1_3QError_Bool_1,Go),
                                               (lizzieLet1_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet1_3QError_Bool_emitted;
  logic [1:0] lizzieLet1_3QError_Bool_done;
  assign lizzieLet1_3QError_Bool_1_d = (lizzieLet1_3QError_Bool_d[0] && (! lizzieLet1_3QError_Bool_emitted[0]));
  assign lizzieLet1_3QError_Bool_2_d = (lizzieLet1_3QError_Bool_d[0] && (! lizzieLet1_3QError_Bool_emitted[1]));
  assign lizzieLet1_3QError_Bool_done = (lizzieLet1_3QError_Bool_emitted | ({lizzieLet1_3QError_Bool_2_d[0],
                                                                             lizzieLet1_3QError_Bool_1_d[0]} & {lizzieLet1_3QError_Bool_2_r,
                                                                                                                lizzieLet1_3QError_Bool_1_r}));
  assign lizzieLet1_3QError_Bool_r = (& lizzieLet1_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet1_3QError_Bool_emitted <= (lizzieLet1_3QError_Bool_r ? 2'd0 :
                                          lizzieLet1_3QError_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet1_3QError_Bool_1,Go) > (lizzieLet1_3QError_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_3QError_Bool_1_bufchan_d;
  logic lizzieLet1_3QError_Bool_1_bufchan_r;
  assign lizzieLet1_3QError_Bool_1_r = ((! lizzieLet1_3QError_Bool_1_bufchan_d[0]) || lizzieLet1_3QError_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QError_Bool_1_r)
        lizzieLet1_3QError_Bool_1_bufchan_d <= lizzieLet1_3QError_Bool_1_d;
  Go_t lizzieLet1_3QError_Bool_1_bufchan_buf;
  assign lizzieLet1_3QError_Bool_1_bufchan_r = (! lizzieLet1_3QError_Bool_1_bufchan_buf[0]);
  assign lizzieLet1_3QError_Bool_1_argbuf_d = (lizzieLet1_3QError_Bool_1_bufchan_buf[0] ? lizzieLet1_3QError_Bool_1_bufchan_buf :
                                               lizzieLet1_3QError_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QError_Bool_1_argbuf_r && lizzieLet1_3QError_Bool_1_bufchan_buf[0]))
        lizzieLet1_3QError_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QError_Bool_1_argbuf_r) && (! lizzieLet1_3QError_Bool_1_bufchan_buf[0])))
        lizzieLet1_3QError_Bool_1_bufchan_buf <= lizzieLet1_3QError_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet1_3QError_Bool_1_argbuf,Go) > (lizzieLet1_3QError_Bool_1_argbuf_0,Int#) */
  assign lizzieLet1_3QError_Bool_1_argbuf_0_d = {32'd0,
                                                 lizzieLet1_3QError_Bool_1_argbuf_d[0]};
  assign lizzieLet1_3QError_Bool_1_argbuf_r = lizzieLet1_3QError_Bool_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet1_3QError_Bool_1_argbuf_0,Int#) > (lizzieLet18_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d;
  logic lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_r;
  assign lizzieLet1_3QError_Bool_1_argbuf_0_r = ((! lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d[0]) || lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet1_3QError_Bool_1_argbuf_0_r)
        lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d <= lizzieLet1_3QError_Bool_1_argbuf_0_d;
  \Int#_t  lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf;
  assign lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_r = (! lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf[0] ? lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf :
                                     lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf[0]))
        lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf[0])))
        lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_buf <= lizzieLet1_3QError_Bool_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QError_Bool_2,Go) > (lizzieLet1_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_3QError_Bool_2_bufchan_d;
  logic lizzieLet1_3QError_Bool_2_bufchan_r;
  assign lizzieLet1_3QError_Bool_2_r = ((! lizzieLet1_3QError_Bool_2_bufchan_d[0]) || lizzieLet1_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QError_Bool_2_r)
        lizzieLet1_3QError_Bool_2_bufchan_d <= lizzieLet1_3QError_Bool_2_d;
  Go_t lizzieLet1_3QError_Bool_2_bufchan_buf;
  assign lizzieLet1_3QError_Bool_2_bufchan_r = (! lizzieLet1_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_3QError_Bool_2_argbuf_d = (lizzieLet1_3QError_Bool_2_bufchan_buf[0] ? lizzieLet1_3QError_Bool_2_bufchan_buf :
                                               lizzieLet1_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QError_Bool_2_argbuf_r && lizzieLet1_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet1_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QError_Bool_2_argbuf_r) && (! lizzieLet1_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet1_3QError_Bool_2_bufchan_buf <= lizzieLet1_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QNode_Bool,Go) > (lizzieLet1_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_3QNode_Bool_bufchan_d;
  logic lizzieLet1_3QNode_Bool_bufchan_r;
  assign lizzieLet1_3QNode_Bool_r = ((! lizzieLet1_3QNode_Bool_bufchan_d[0]) || lizzieLet1_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QNode_Bool_r)
        lizzieLet1_3QNode_Bool_bufchan_d <= lizzieLet1_3QNode_Bool_d;
  Go_t lizzieLet1_3QNode_Bool_bufchan_buf;
  assign lizzieLet1_3QNode_Bool_bufchan_r = (! lizzieLet1_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet1_3QNode_Bool_1_argbuf_d = (lizzieLet1_3QNode_Bool_bufchan_buf[0] ? lizzieLet1_3QNode_Bool_bufchan_buf :
                                              lizzieLet1_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QNode_Bool_1_argbuf_r && lizzieLet1_3QNode_Bool_bufchan_buf[0]))
        lizzieLet1_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QNode_Bool_1_argbuf_r) && (! lizzieLet1_3QNode_Bool_bufchan_buf[0])))
        lizzieLet1_3QNode_Bool_bufchan_buf <= lizzieLet1_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet1_3QNone_Bool,Go) > [(lizzieLet1_3QNone_Bool_1,Go),
                                              (lizzieLet1_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet1_3QNone_Bool_emitted;
  logic [1:0] lizzieLet1_3QNone_Bool_done;
  assign lizzieLet1_3QNone_Bool_1_d = (lizzieLet1_3QNone_Bool_d[0] && (! lizzieLet1_3QNone_Bool_emitted[0]));
  assign lizzieLet1_3QNone_Bool_2_d = (lizzieLet1_3QNone_Bool_d[0] && (! lizzieLet1_3QNone_Bool_emitted[1]));
  assign lizzieLet1_3QNone_Bool_done = (lizzieLet1_3QNone_Bool_emitted | ({lizzieLet1_3QNone_Bool_2_d[0],
                                                                           lizzieLet1_3QNone_Bool_1_d[0]} & {lizzieLet1_3QNone_Bool_2_r,
                                                                                                             lizzieLet1_3QNone_Bool_1_r}));
  assign lizzieLet1_3QNone_Bool_r = (& lizzieLet1_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet1_3QNone_Bool_emitted <= (lizzieLet1_3QNone_Bool_r ? 2'd0 :
                                         lizzieLet1_3QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet1_3QNone_Bool_1,Go) > (lizzieLet1_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_3QNone_Bool_1_bufchan_d;
  logic lizzieLet1_3QNone_Bool_1_bufchan_r;
  assign lizzieLet1_3QNone_Bool_1_r = ((! lizzieLet1_3QNone_Bool_1_bufchan_d[0]) || lizzieLet1_3QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QNone_Bool_1_r)
        lizzieLet1_3QNone_Bool_1_bufchan_d <= lizzieLet1_3QNone_Bool_1_d;
  Go_t lizzieLet1_3QNone_Bool_1_bufchan_buf;
  assign lizzieLet1_3QNone_Bool_1_bufchan_r = (! lizzieLet1_3QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet1_3QNone_Bool_1_argbuf_d = (lizzieLet1_3QNone_Bool_1_bufchan_buf[0] ? lizzieLet1_3QNone_Bool_1_bufchan_buf :
                                              lizzieLet1_3QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QNone_Bool_1_argbuf_r && lizzieLet1_3QNone_Bool_1_bufchan_buf[0]))
        lizzieLet1_3QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QNone_Bool_1_argbuf_r) && (! lizzieLet1_3QNone_Bool_1_bufchan_buf[0])))
        lizzieLet1_3QNone_Bool_1_bufchan_buf <= lizzieLet1_3QNone_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet1_3QNone_Bool_1_argbuf,Go) > (lizzieLet1_3QNone_Bool_1_argbuf_0,Int#) */
  assign lizzieLet1_3QNone_Bool_1_argbuf_0_d = {32'd0,
                                                lizzieLet1_3QNone_Bool_1_argbuf_d[0]};
  assign lizzieLet1_3QNone_Bool_1_argbuf_r = lizzieLet1_3QNone_Bool_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet1_3QNone_Bool_1_argbuf_0,Int#) > (lizzieLet18_1_argbuf,Int#) */
  \Int#_t  lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d;
  logic lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_r;
  assign lizzieLet1_3QNone_Bool_1_argbuf_0_r = ((! lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d[0]) || lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet1_3QNone_Bool_1_argbuf_0_r)
        lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d <= lizzieLet1_3QNone_Bool_1_argbuf_0_d;
  \Int#_t  lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf;
  assign lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_r = (! lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf[0] ? lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf :
                                   lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf[0]))
        lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf[0])))
        lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_buf <= lizzieLet1_3QNone_Bool_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QNone_Bool_2,Go) > (lizzieLet1_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_3QNone_Bool_2_bufchan_d;
  logic lizzieLet1_3QNone_Bool_2_bufchan_r;
  assign lizzieLet1_3QNone_Bool_2_r = ((! lizzieLet1_3QNone_Bool_2_bufchan_d[0]) || lizzieLet1_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QNone_Bool_2_r)
        lizzieLet1_3QNone_Bool_2_bufchan_d <= lizzieLet1_3QNone_Bool_2_d;
  Go_t lizzieLet1_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet1_3QNone_Bool_2_bufchan_r = (! lizzieLet1_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_3QNone_Bool_2_argbuf_d = (lizzieLet1_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet1_3QNone_Bool_2_bufchan_buf :
                                              lizzieLet1_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QNone_Bool_2_argbuf_r && lizzieLet1_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet1_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QNone_Bool_2_argbuf_r) && (! lizzieLet1_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet1_3QNone_Bool_2_bufchan_buf <= lizzieLet1_3QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet1_3QNone_Bool_2_argbuf,Go),
                           (lizzieLet44_3Lcall_$wnnz0_1_argbuf,Go),
                           (lizzieLet1_3QVal_Bool_2_argbuf,Go),
                           (lizzieLet1_3QError_Bool_2_argbuf,Go)] > (go_19_goMux_choice,C4) (go_19_goMux_data,Go) */
  logic [3:0] lizzieLet1_3QNone_Bool_2_argbuf_select_d;
  assign lizzieLet1_3QNone_Bool_2_argbuf_select_d = ((| lizzieLet1_3QNone_Bool_2_argbuf_select_q) ? lizzieLet1_3QNone_Bool_2_argbuf_select_q :
                                                     (lizzieLet1_3QNone_Bool_2_argbuf_d[0] ? 4'd1 :
                                                      (lizzieLet44_3Lcall_$wnnz0_1_argbuf_d[0] ? 4'd2 :
                                                       (lizzieLet1_3QVal_Bool_2_argbuf_d[0] ? 4'd4 :
                                                        (lizzieLet1_3QError_Bool_2_argbuf_d[0] ? 4'd8 :
                                                         4'd0)))));
  logic [3:0] lizzieLet1_3QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet1_3QNone_Bool_2_argbuf_select_q <= (lizzieLet1_3QNone_Bool_2_argbuf_done ? 4'd0 :
                                                   lizzieLet1_3QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet1_3QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet1_3QNone_Bool_2_argbuf_emit_q <= (lizzieLet1_3QNone_Bool_2_argbuf_done ? 2'd0 :
                                                 lizzieLet1_3QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet1_3QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet1_3QNone_Bool_2_argbuf_emit_d = (lizzieLet1_3QNone_Bool_2_argbuf_emit_q | ({go_19_goMux_choice_d[0],
                                                                                              go_19_goMux_data_d[0]} & {go_19_goMux_choice_r,
                                                                                                                        go_19_goMux_data_r}));
  logic lizzieLet1_3QNone_Bool_2_argbuf_done;
  assign lizzieLet1_3QNone_Bool_2_argbuf_done = (& lizzieLet1_3QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet1_3QError_Bool_2_argbuf_r,
          lizzieLet1_3QVal_Bool_2_argbuf_r,
          lizzieLet44_3Lcall_$wnnz0_1_argbuf_r,
          lizzieLet1_3QNone_Bool_2_argbuf_r} = (lizzieLet1_3QNone_Bool_2_argbuf_done ? lizzieLet1_3QNone_Bool_2_argbuf_select_d :
                                                4'd0);
  assign go_19_goMux_data_d = ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet1_3QNone_Bool_2_argbuf_d :
                               ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet44_3Lcall_$wnnz0_1_argbuf_d :
                                ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet1_3QVal_Bool_2_argbuf_d :
                                 ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet1_3QError_Bool_2_argbuf_d :
                                  1'd0))));
  assign go_19_goMux_choice_d = ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet1_3QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet1_3QNone_Bool_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet1_3QVal_Bool,Go) > [(lizzieLet1_3QVal_Bool_1,Go),
                                             (lizzieLet1_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet1_3QVal_Bool_emitted;
  logic [1:0] lizzieLet1_3QVal_Bool_done;
  assign lizzieLet1_3QVal_Bool_1_d = (lizzieLet1_3QVal_Bool_d[0] && (! lizzieLet1_3QVal_Bool_emitted[0]));
  assign lizzieLet1_3QVal_Bool_2_d = (lizzieLet1_3QVal_Bool_d[0] && (! lizzieLet1_3QVal_Bool_emitted[1]));
  assign lizzieLet1_3QVal_Bool_done = (lizzieLet1_3QVal_Bool_emitted | ({lizzieLet1_3QVal_Bool_2_d[0],
                                                                         lizzieLet1_3QVal_Bool_1_d[0]} & {lizzieLet1_3QVal_Bool_2_r,
                                                                                                          lizzieLet1_3QVal_Bool_1_r}));
  assign lizzieLet1_3QVal_Bool_r = (& lizzieLet1_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet1_3QVal_Bool_emitted <= (lizzieLet1_3QVal_Bool_r ? 2'd0 :
                                        lizzieLet1_3QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet1_3QVal_Bool_1,Go) > (lizzieLet1_3QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_3QVal_Bool_1_bufchan_d;
  logic lizzieLet1_3QVal_Bool_1_bufchan_r;
  assign lizzieLet1_3QVal_Bool_1_r = ((! lizzieLet1_3QVal_Bool_1_bufchan_d[0]) || lizzieLet1_3QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QVal_Bool_1_r)
        lizzieLet1_3QVal_Bool_1_bufchan_d <= lizzieLet1_3QVal_Bool_1_d;
  Go_t lizzieLet1_3QVal_Bool_1_bufchan_buf;
  assign lizzieLet1_3QVal_Bool_1_bufchan_r = (! lizzieLet1_3QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet1_3QVal_Bool_1_argbuf_d = (lizzieLet1_3QVal_Bool_1_bufchan_buf[0] ? lizzieLet1_3QVal_Bool_1_bufchan_buf :
                                             lizzieLet1_3QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QVal_Bool_1_argbuf_r && lizzieLet1_3QVal_Bool_1_bufchan_buf[0]))
        lizzieLet1_3QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QVal_Bool_1_argbuf_r) && (! lizzieLet1_3QVal_Bool_1_bufchan_buf[0])))
        lizzieLet1_3QVal_Bool_1_bufchan_buf <= lizzieLet1_3QVal_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet1_3QVal_Bool_1_argbuf,Go) > (lizzieLet1_3QVal_Bool_1_argbuf_1,Int#) */
  assign lizzieLet1_3QVal_Bool_1_argbuf_1_d = {32'd1,
                                               lizzieLet1_3QVal_Bool_1_argbuf_d[0]};
  assign lizzieLet1_3QVal_Bool_1_argbuf_r = lizzieLet1_3QVal_Bool_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet1_3QVal_Bool_1_argbuf_1,Int#) > (lizzieLet19_1_argbuf,Int#) */
  \Int#_t  lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d;
  logic lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_r;
  assign lizzieLet1_3QVal_Bool_1_argbuf_1_r = ((! lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d[0]) || lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet1_3QVal_Bool_1_argbuf_1_r)
        lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d <= lizzieLet1_3QVal_Bool_1_argbuf_1_d;
  \Int#_t  lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf;
  assign lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_r = (! lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf[0] ? lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf :
                                   lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf[0]))
        lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf[0])))
        lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_buf <= lizzieLet1_3QVal_Bool_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QVal_Bool_2,Go) > (lizzieLet1_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_3QVal_Bool_2_bufchan_d;
  logic lizzieLet1_3QVal_Bool_2_bufchan_r;
  assign lizzieLet1_3QVal_Bool_2_r = ((! lizzieLet1_3QVal_Bool_2_bufchan_d[0]) || lizzieLet1_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QVal_Bool_2_r)
        lizzieLet1_3QVal_Bool_2_bufchan_d <= lizzieLet1_3QVal_Bool_2_d;
  Go_t lizzieLet1_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet1_3QVal_Bool_2_bufchan_r = (! lizzieLet1_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_3QVal_Bool_2_argbuf_d = (lizzieLet1_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet1_3QVal_Bool_2_bufchan_buf :
                                             lizzieLet1_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QVal_Bool_2_argbuf_r && lizzieLet1_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet1_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QVal_Bool_2_argbuf_r) && (! lizzieLet1_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet1_3QVal_Bool_2_bufchan_buf <= lizzieLet1_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CT$wnnz) : (lizzieLet1_4,QTree_Bool) (sc_0_goMux_mux,Pointer_CT$wnnz) > [(lizzieLet1_4QNone_Bool,Pointer_CT$wnnz),
                                                                                           (lizzieLet1_4QVal_Bool,Pointer_CT$wnnz),
                                                                                           (lizzieLet1_4QNode_Bool,Pointer_CT$wnnz),
                                                                                           (lizzieLet1_4QError_Bool,Pointer_CT$wnnz)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet1_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet1_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet1_4QNone_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet1_4QVal_Bool_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet1_4QError_Bool_d = {sc_0_goMux_mux_d[16:1],
                                      sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet1_4QError_Bool_r,
                                                          lizzieLet1_4QNode_Bool_r,
                                                          lizzieLet1_4QVal_Bool_r,
                                                          lizzieLet1_4QNone_Bool_r}));
  assign lizzieLet1_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet1_4QError_Bool,Pointer_CT$wnnz) > (lizzieLet1_4QError_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet1_4QError_Bool_bufchan_d;
  logic lizzieLet1_4QError_Bool_bufchan_r;
  assign lizzieLet1_4QError_Bool_r = ((! lizzieLet1_4QError_Bool_bufchan_d[0]) || lizzieLet1_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QError_Bool_r)
        lizzieLet1_4QError_Bool_bufchan_d <= lizzieLet1_4QError_Bool_d;
  Pointer_CT$wnnz_t lizzieLet1_4QError_Bool_bufchan_buf;
  assign lizzieLet1_4QError_Bool_bufchan_r = (! lizzieLet1_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QError_Bool_1_argbuf_d = (lizzieLet1_4QError_Bool_bufchan_buf[0] ? lizzieLet1_4QError_Bool_bufchan_buf :
                                               lizzieLet1_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QError_Bool_1_argbuf_r && lizzieLet1_4QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QError_Bool_1_argbuf_r) && (! lizzieLet1_4QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QError_Bool_bufchan_buf <= lizzieLet1_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz3) : [(lizzieLet1_4QNode_Bool,Pointer_CT$wnnz),
                            (q4a87_destruct,Pointer_QTree_Bool),
                            (q3a86_destruct,Pointer_QTree_Bool),
                            (q2a85_destruct,Pointer_QTree_Bool)] > (lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3,CT$wnnz) */
  assign lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d = Lcall_$wnnz3_dc((& {lizzieLet1_4QNode_Bool_d[0],
                                                                                           q4a87_destruct_d[0],
                                                                                           q3a86_destruct_d[0],
                                                                                           q2a85_destruct_d[0]}), lizzieLet1_4QNode_Bool_d, q4a87_destruct_d, q3a86_destruct_d, q2a85_destruct_d);
  assign {lizzieLet1_4QNode_Bool_r,
          q4a87_destruct_r,
          q3a86_destruct_r,
          q2a85_destruct_r} = {4 {(lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r && lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3,CT$wnnz) > (lizzieLet2_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d;
  logic lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r;
  assign lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r = ((! lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d[0]) || lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d <= {115'd0,
                                                                              1'd0};
    else
      if (lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_r)
        lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d <= lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_d;
  CT$wnnz_t lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_r = (! lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf :
                                  lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                  1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_buf <= lizzieLet1_4QNode_Bool_1q4a87_1q3a86_1q2a85_1Lcall_$wnnz3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet1_4QNone_Bool,Pointer_CT$wnnz) > (lizzieLet1_4QNone_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet1_4QNone_Bool_bufchan_d;
  logic lizzieLet1_4QNone_Bool_bufchan_r;
  assign lizzieLet1_4QNone_Bool_r = ((! lizzieLet1_4QNone_Bool_bufchan_d[0]) || lizzieLet1_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNone_Bool_r)
        lizzieLet1_4QNone_Bool_bufchan_d <= lizzieLet1_4QNone_Bool_d;
  Pointer_CT$wnnz_t lizzieLet1_4QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QNone_Bool_bufchan_r = (! lizzieLet1_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNone_Bool_1_argbuf_d = (lizzieLet1_4QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QNone_Bool_bufchan_buf :
                                              lizzieLet1_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNone_Bool_1_argbuf_r && lizzieLet1_4QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QNone_Bool_bufchan_buf <= lizzieLet1_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet1_4QVal_Bool,Pointer_CT$wnnz) > (lizzieLet1_4QVal_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet1_4QVal_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_r = ((! lizzieLet1_4QVal_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_r)
        lizzieLet1_4QVal_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_d;
  Pointer_CT$wnnz_t lizzieLet1_4QVal_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_bufchan_buf :
                                             lizzieLet1_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet23_1wild3XR_1_1_Eq,Bool) > (lizzieLet24_1_argbuf,Bool) */
  Bool_t lizzieLet23_1wild3XR_1_1_Eq_bufchan_d;
  logic lizzieLet23_1wild3XR_1_1_Eq_bufchan_r;
  assign lizzieLet23_1wild3XR_1_1_Eq_r = ((! lizzieLet23_1wild3XR_1_1_Eq_bufchan_d[0]) || lizzieLet23_1wild3XR_1_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet23_1wild3XR_1_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet23_1wild3XR_1_1_Eq_r)
        lizzieLet23_1wild3XR_1_1_Eq_bufchan_d <= lizzieLet23_1wild3XR_1_1_Eq_d;
  Bool_t lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf;
  assign lizzieLet23_1wild3XR_1_1_Eq_bufchan_r = (! lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf[0]);
  assign lizzieLet24_1_argbuf_d = (lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf[0] ? lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf :
                                   lizzieLet23_1wild3XR_1_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf[0]))
        lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf[0])))
        lizzieLet23_1wild3XR_1_1_Eq_bufchan_buf <= lizzieLet23_1wild3XR_1_1_Eq_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet25_1,MyBool) (lizzieLet12_4QVal_Int_5QNone_Int_3I#_3,Go) > [(lizzieLet25_1MyFalse,Go),
                                                                                      (lizzieLet25_1MyTrue,Go)] */
  logic [1:0] \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet25_1_d[0] && \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_d [0]))
      unique case (lizzieLet25_1_d[1:1])
        1'd0: \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd  = 2'd1;
        1'd1: \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd  = 2'd2;
        default: \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd  = 2'd0;
      endcase
    else \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd  = 2'd0;
  assign lizzieLet25_1MyFalse_d = \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd [0];
  assign lizzieLet25_1MyTrue_d = \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd [1];
  assign \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_r  = (| (\lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_onehotd  & {lizzieLet25_1MyTrue_r,
                                                                                                              lizzieLet25_1MyFalse_r}));
  assign lizzieLet25_1_r = \lizzieLet12_4QVal_Int_5QNone_Int_3I#_3_r ;
  
  /* fork (Ty Go) : (lizzieLet25_1MyFalse,Go) > [(lizzieLet25_1MyFalse_1,Go),
                                            (lizzieLet25_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet25_1MyFalse_emitted;
  logic [1:0] lizzieLet25_1MyFalse_done;
  assign lizzieLet25_1MyFalse_1_d = (lizzieLet25_1MyFalse_d[0] && (! lizzieLet25_1MyFalse_emitted[0]));
  assign lizzieLet25_1MyFalse_2_d = (lizzieLet25_1MyFalse_d[0] && (! lizzieLet25_1MyFalse_emitted[1]));
  assign lizzieLet25_1MyFalse_done = (lizzieLet25_1MyFalse_emitted | ({lizzieLet25_1MyFalse_2_d[0],
                                                                       lizzieLet25_1MyFalse_1_d[0]} & {lizzieLet25_1MyFalse_2_r,
                                                                                                       lizzieLet25_1MyFalse_1_r}));
  assign lizzieLet25_1MyFalse_r = (& lizzieLet25_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet25_1MyFalse_emitted <= (lizzieLet25_1MyFalse_r ? 2'd0 :
                                       lizzieLet25_1MyFalse_done);
  
  /* buf (Ty Go) : (lizzieLet25_1MyFalse_1,Go) > (lizzieLet25_1MyFalse_1_argbuf,Go) */
  Go_t lizzieLet25_1MyFalse_1_bufchan_d;
  logic lizzieLet25_1MyFalse_1_bufchan_r;
  assign lizzieLet25_1MyFalse_1_r = ((! lizzieLet25_1MyFalse_1_bufchan_d[0]) || lizzieLet25_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_1MyFalse_1_r)
        lizzieLet25_1MyFalse_1_bufchan_d <= lizzieLet25_1MyFalse_1_d;
  Go_t lizzieLet25_1MyFalse_1_bufchan_buf;
  assign lizzieLet25_1MyFalse_1_bufchan_r = (! lizzieLet25_1MyFalse_1_bufchan_buf[0]);
  assign lizzieLet25_1MyFalse_1_argbuf_d = (lizzieLet25_1MyFalse_1_bufchan_buf[0] ? lizzieLet25_1MyFalse_1_bufchan_buf :
                                            lizzieLet25_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_1MyFalse_1_argbuf_r && lizzieLet25_1MyFalse_1_bufchan_buf[0]))
        lizzieLet25_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_1MyFalse_1_argbuf_r) && (! lizzieLet25_1MyFalse_1_bufchan_buf[0])))
        lizzieLet25_1MyFalse_1_bufchan_buf <= lizzieLet25_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet25_1MyFalse_1_argbuf,Go)] > (f''''''''1TupGo3,TupGo) */
  assign \f''''''''1TupGo3_d  = TupGo_dc((& {lizzieLet25_1MyFalse_1_argbuf_d[0]}), lizzieLet25_1MyFalse_1_argbuf_d);
  assign {lizzieLet25_1MyFalse_1_argbuf_r} = {1 {(\f''''''''1TupGo3_r  && \f''''''''1TupGo3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet25_1MyFalse_2,Go) > (lizzieLet25_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet25_1MyFalse_2_bufchan_d;
  logic lizzieLet25_1MyFalse_2_bufchan_r;
  assign lizzieLet25_1MyFalse_2_r = ((! lizzieLet25_1MyFalse_2_bufchan_d[0]) || lizzieLet25_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_1MyFalse_2_r)
        lizzieLet25_1MyFalse_2_bufchan_d <= lizzieLet25_1MyFalse_2_d;
  Go_t lizzieLet25_1MyFalse_2_bufchan_buf;
  assign lizzieLet25_1MyFalse_2_bufchan_r = (! lizzieLet25_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet25_1MyFalse_2_argbuf_d = (lizzieLet25_1MyFalse_2_bufchan_buf[0] ? lizzieLet25_1MyFalse_2_bufchan_buf :
                                            lizzieLet25_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_1MyFalse_2_argbuf_r && lizzieLet25_1MyFalse_2_bufchan_buf[0]))
        lizzieLet25_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_1MyFalse_2_argbuf_r) && (! lizzieLet25_1MyFalse_2_bufchan_buf[0])))
        lizzieLet25_1MyFalse_2_bufchan_buf <= lizzieLet25_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet25_1MyTrue,Go) > [(lizzieLet25_1MyTrue_1,Go),
                                           (lizzieLet25_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet25_1MyTrue_emitted;
  logic [1:0] lizzieLet25_1MyTrue_done;
  assign lizzieLet25_1MyTrue_1_d = (lizzieLet25_1MyTrue_d[0] && (! lizzieLet25_1MyTrue_emitted[0]));
  assign lizzieLet25_1MyTrue_2_d = (lizzieLet25_1MyTrue_d[0] && (! lizzieLet25_1MyTrue_emitted[1]));
  assign lizzieLet25_1MyTrue_done = (lizzieLet25_1MyTrue_emitted | ({lizzieLet25_1MyTrue_2_d[0],
                                                                     lizzieLet25_1MyTrue_1_d[0]} & {lizzieLet25_1MyTrue_2_r,
                                                                                                    lizzieLet25_1MyTrue_1_r}));
  assign lizzieLet25_1MyTrue_r = (& lizzieLet25_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet25_1MyTrue_emitted <= (lizzieLet25_1MyTrue_r ? 2'd0 :
                                      lizzieLet25_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet25_1MyTrue_1,Go)] > (lizzieLet25_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign lizzieLet25_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet25_1MyTrue_1_d[0]}), lizzieLet25_1MyTrue_1_d);
  assign {lizzieLet25_1MyTrue_1_r} = {1 {(lizzieLet25_1MyTrue_1QNone_Bool_r && lizzieLet25_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet25_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet27_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d;
  logic lizzieLet25_1MyTrue_1QNone_Bool_bufchan_r;
  assign lizzieLet25_1MyTrue_1QNone_Bool_r = ((! lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d[0]) || lizzieLet25_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet25_1MyTrue_1QNone_Bool_r)
        lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d <= lizzieLet25_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf;
  assign lizzieLet25_1MyTrue_1QNone_Bool_bufchan_r = (! lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf[0] ? lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf :
                                   lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        lizzieLet25_1MyTrue_1QNone_Bool_bufchan_buf <= lizzieLet25_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet25_1MyTrue_2,Go) > (lizzieLet25_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet25_1MyTrue_2_bufchan_d;
  logic lizzieLet25_1MyTrue_2_bufchan_r;
  assign lizzieLet25_1MyTrue_2_r = ((! lizzieLet25_1MyTrue_2_bufchan_d[0]) || lizzieLet25_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet25_1MyTrue_2_r)
        lizzieLet25_1MyTrue_2_bufchan_d <= lizzieLet25_1MyTrue_2_d;
  Go_t lizzieLet25_1MyTrue_2_bufchan_buf;
  assign lizzieLet25_1MyTrue_2_bufchan_r = (! lizzieLet25_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet25_1MyTrue_2_argbuf_d = (lizzieLet25_1MyTrue_2_bufchan_buf[0] ? lizzieLet25_1MyTrue_2_bufchan_buf :
                                           lizzieLet25_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet25_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet25_1MyTrue_2_argbuf_r && lizzieLet25_1MyTrue_2_bufchan_buf[0]))
        lizzieLet25_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet25_1MyTrue_2_argbuf_r) && (! lizzieLet25_1MyTrue_2_bufchan_buf[0])))
        lizzieLet25_1MyTrue_2_bufchan_buf <= lizzieLet25_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f) : (lizzieLet25_2,MyBool) (lizzieLet12_4QVal_Int_5QNone_Int_4I#,Pointer_CTf_f) > [(lizzieLet25_2MyFalse,Pointer_CTf_f),
                                                                                                          (lizzieLet25_2MyTrue,Pointer_CTf_f)] */
  logic [1:0] \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd ;
  always_comb
    if ((lizzieLet25_2_d[0] && \lizzieLet12_4QVal_Int_5QNone_Int_4I#_d [0]))
      unique case (lizzieLet25_2_d[1:1])
        1'd0: \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd  = 2'd1;
        1'd1: \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd  = 2'd2;
        default: \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd  = 2'd0;
      endcase
    else \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd  = 2'd0;
  assign lizzieLet25_2MyFalse_d = {\lizzieLet12_4QVal_Int_5QNone_Int_4I#_d [16:1],
                                   \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd [0]};
  assign lizzieLet25_2MyTrue_d = {\lizzieLet12_4QVal_Int_5QNone_Int_4I#_d [16:1],
                                  \lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd [1]};
  assign \lizzieLet12_4QVal_Int_5QNone_Int_4I#_r  = (| (\lizzieLet12_4QVal_Int_5QNone_Int_4I#_onehotd  & {lizzieLet25_2MyTrue_r,
                                                                                                          lizzieLet25_2MyFalse_r}));
  assign lizzieLet25_2_r = \lizzieLet12_4QVal_Int_5QNone_Int_4I#_r ;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet25_2MyFalse,Pointer_CTf_f) > (lizzieLet25_2MyFalse_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet25_2MyFalse_bufchan_d;
  logic lizzieLet25_2MyFalse_bufchan_r;
  assign lizzieLet25_2MyFalse_r = ((! lizzieLet25_2MyFalse_bufchan_d[0]) || lizzieLet25_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet25_2MyFalse_r)
        lizzieLet25_2MyFalse_bufchan_d <= lizzieLet25_2MyFalse_d;
  Pointer_CTf_f_t lizzieLet25_2MyFalse_bufchan_buf;
  assign lizzieLet25_2MyFalse_bufchan_r = (! lizzieLet25_2MyFalse_bufchan_buf[0]);
  assign lizzieLet25_2MyFalse_1_argbuf_d = (lizzieLet25_2MyFalse_bufchan_buf[0] ? lizzieLet25_2MyFalse_bufchan_buf :
                                            lizzieLet25_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet25_2MyFalse_1_argbuf_r && lizzieLet25_2MyFalse_bufchan_buf[0]))
        lizzieLet25_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet25_2MyFalse_1_argbuf_r) && (! lizzieLet25_2MyFalse_bufchan_buf[0])))
        lizzieLet25_2MyFalse_bufchan_buf <= lizzieLet25_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet25_2MyTrue,Pointer_CTf_f) > (lizzieLet25_2MyTrue_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet25_2MyTrue_bufchan_d;
  logic lizzieLet25_2MyTrue_bufchan_r;
  assign lizzieLet25_2MyTrue_r = ((! lizzieLet25_2MyTrue_bufchan_d[0]) || lizzieLet25_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet25_2MyTrue_r)
        lizzieLet25_2MyTrue_bufchan_d <= lizzieLet25_2MyTrue_d;
  Pointer_CTf_f_t lizzieLet25_2MyTrue_bufchan_buf;
  assign lizzieLet25_2MyTrue_bufchan_r = (! lizzieLet25_2MyTrue_bufchan_buf[0]);
  assign lizzieLet25_2MyTrue_1_argbuf_d = (lizzieLet25_2MyTrue_bufchan_buf[0] ? lizzieLet25_2MyTrue_bufchan_buf :
                                           lizzieLet25_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet25_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet25_2MyTrue_1_argbuf_r && lizzieLet25_2MyTrue_bufchan_buf[0]))
        lizzieLet25_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet25_2MyTrue_1_argbuf_r) && (! lizzieLet25_2MyTrue_bufchan_buf[0])))
        lizzieLet25_2MyTrue_bufchan_buf <= lizzieLet25_2MyTrue_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet28_1wild4XU_1_Eq,Bool) > (lizzieLet29_1_argbuf,Bool) */
  Bool_t lizzieLet28_1wild4XU_1_Eq_bufchan_d;
  logic lizzieLet28_1wild4XU_1_Eq_bufchan_r;
  assign lizzieLet28_1wild4XU_1_Eq_r = ((! lizzieLet28_1wild4XU_1_Eq_bufchan_d[0]) || lizzieLet28_1wild4XU_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1wild4XU_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet28_1wild4XU_1_Eq_r)
        lizzieLet28_1wild4XU_1_Eq_bufchan_d <= lizzieLet28_1wild4XU_1_Eq_d;
  Bool_t lizzieLet28_1wild4XU_1_Eq_bufchan_buf;
  assign lizzieLet28_1wild4XU_1_Eq_bufchan_r = (! lizzieLet28_1wild4XU_1_Eq_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet28_1wild4XU_1_Eq_bufchan_buf[0] ? lizzieLet28_1wild4XU_1_Eq_bufchan_buf :
                                   lizzieLet28_1wild4XU_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1wild4XU_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet28_1wild4XU_1_Eq_bufchan_buf[0]))
        lizzieLet28_1wild4XU_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet28_1wild4XU_1_Eq_bufchan_buf[0])))
        lizzieLet28_1wild4XU_1_Eq_bufchan_buf <= lizzieLet28_1wild4XU_1_Eq_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet30_1,MyBool) (lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3,Go) > [(lizzieLet30_1MyFalse,Go),
                                                                                         (lizzieLet30_1MyTrue,Go)] */
  logic [1:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet30_1_d[0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_d [0]))
      unique case (lizzieLet30_1_d[1:1])
        1'd0: \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd  = 2'd1;
        1'd1: \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd  = 2'd2;
        default:
          \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd  = 2'd0;
      endcase
    else \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd  = 2'd0;
  assign lizzieLet30_1MyFalse_d = \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd [0];
  assign lizzieLet30_1MyTrue_d = \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd [1];
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_r  = (| (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_onehotd  & {lizzieLet30_1MyTrue_r,
                                                                                                                    lizzieLet30_1MyFalse_r}));
  assign lizzieLet30_1_r = \lizzieLet12_4QVal_Int_5QVal_Int_5I#_3I#_3_r ;
  
  /* fork (Ty Go) : (lizzieLet30_1MyFalse,Go) > [(lizzieLet30_1MyFalse_1,Go),
                                            (lizzieLet30_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet30_1MyFalse_emitted;
  logic [1:0] lizzieLet30_1MyFalse_done;
  assign lizzieLet30_1MyFalse_1_d = (lizzieLet30_1MyFalse_d[0] && (! lizzieLet30_1MyFalse_emitted[0]));
  assign lizzieLet30_1MyFalse_2_d = (lizzieLet30_1MyFalse_d[0] && (! lizzieLet30_1MyFalse_emitted[1]));
  assign lizzieLet30_1MyFalse_done = (lizzieLet30_1MyFalse_emitted | ({lizzieLet30_1MyFalse_2_d[0],
                                                                       lizzieLet30_1MyFalse_1_d[0]} & {lizzieLet30_1MyFalse_2_r,
                                                                                                       lizzieLet30_1MyFalse_1_r}));
  assign lizzieLet30_1MyFalse_r = (& lizzieLet30_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet30_1MyFalse_emitted <= (lizzieLet30_1MyFalse_r ? 2'd0 :
                                       lizzieLet30_1MyFalse_done);
  
  /* buf (Ty Go) : (lizzieLet30_1MyFalse_1,Go) > (lizzieLet30_1MyFalse_1_argbuf,Go) */
  Go_t lizzieLet30_1MyFalse_1_bufchan_d;
  logic lizzieLet30_1MyFalse_1_bufchan_r;
  assign lizzieLet30_1MyFalse_1_r = ((! lizzieLet30_1MyFalse_1_bufchan_d[0]) || lizzieLet30_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_1MyFalse_1_r)
        lizzieLet30_1MyFalse_1_bufchan_d <= lizzieLet30_1MyFalse_1_d;
  Go_t lizzieLet30_1MyFalse_1_bufchan_buf;
  assign lizzieLet30_1MyFalse_1_bufchan_r = (! lizzieLet30_1MyFalse_1_bufchan_buf[0]);
  assign lizzieLet30_1MyFalse_1_argbuf_d = (lizzieLet30_1MyFalse_1_bufchan_buf[0] ? lizzieLet30_1MyFalse_1_bufchan_buf :
                                            lizzieLet30_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_1MyFalse_1_argbuf_r && lizzieLet30_1MyFalse_1_bufchan_buf[0]))
        lizzieLet30_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_1MyFalse_1_argbuf_r) && (! lizzieLet30_1MyFalse_1_bufchan_buf[0])))
        lizzieLet30_1MyFalse_1_bufchan_buf <= lizzieLet30_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet30_1MyFalse_1_argbuf,Go)] > (f''''''''1TupGo4,TupGo) */
  assign \f''''''''1TupGo4_d  = TupGo_dc((& {lizzieLet30_1MyFalse_1_argbuf_d[0]}), lizzieLet30_1MyFalse_1_argbuf_d);
  assign {lizzieLet30_1MyFalse_1_argbuf_r} = {1 {(\f''''''''1TupGo4_r  && \f''''''''1TupGo4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet30_1MyFalse_2,Go) > (lizzieLet30_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet30_1MyFalse_2_bufchan_d;
  logic lizzieLet30_1MyFalse_2_bufchan_r;
  assign lizzieLet30_1MyFalse_2_r = ((! lizzieLet30_1MyFalse_2_bufchan_d[0]) || lizzieLet30_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_1MyFalse_2_r)
        lizzieLet30_1MyFalse_2_bufchan_d <= lizzieLet30_1MyFalse_2_d;
  Go_t lizzieLet30_1MyFalse_2_bufchan_buf;
  assign lizzieLet30_1MyFalse_2_bufchan_r = (! lizzieLet30_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet30_1MyFalse_2_argbuf_d = (lizzieLet30_1MyFalse_2_bufchan_buf[0] ? lizzieLet30_1MyFalse_2_bufchan_buf :
                                            lizzieLet30_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_1MyFalse_2_argbuf_r && lizzieLet30_1MyFalse_2_bufchan_buf[0]))
        lizzieLet30_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_1MyFalse_2_argbuf_r) && (! lizzieLet30_1MyFalse_2_bufchan_buf[0])))
        lizzieLet30_1MyFalse_2_bufchan_buf <= lizzieLet30_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet30_1MyTrue,Go) > [(lizzieLet30_1MyTrue_1,Go),
                                           (lizzieLet30_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet30_1MyTrue_emitted;
  logic [1:0] lizzieLet30_1MyTrue_done;
  assign lizzieLet30_1MyTrue_1_d = (lizzieLet30_1MyTrue_d[0] && (! lizzieLet30_1MyTrue_emitted[0]));
  assign lizzieLet30_1MyTrue_2_d = (lizzieLet30_1MyTrue_d[0] && (! lizzieLet30_1MyTrue_emitted[1]));
  assign lizzieLet30_1MyTrue_done = (lizzieLet30_1MyTrue_emitted | ({lizzieLet30_1MyTrue_2_d[0],
                                                                     lizzieLet30_1MyTrue_1_d[0]} & {lizzieLet30_1MyTrue_2_r,
                                                                                                    lizzieLet30_1MyTrue_1_r}));
  assign lizzieLet30_1MyTrue_r = (& lizzieLet30_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet30_1MyTrue_emitted <= (lizzieLet30_1MyTrue_r ? 2'd0 :
                                      lizzieLet30_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet30_1MyTrue_1,Go)] > (lizzieLet30_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign lizzieLet30_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet30_1MyTrue_1_d[0]}), lizzieLet30_1MyTrue_1_d);
  assign {lizzieLet30_1MyTrue_1_r} = {1 {(lizzieLet30_1MyTrue_1QNone_Bool_r && lizzieLet30_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet30_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet32_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d;
  logic lizzieLet30_1MyTrue_1QNone_Bool_bufchan_r;
  assign lizzieLet30_1MyTrue_1QNone_Bool_r = ((! lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d[0]) || lizzieLet30_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet30_1MyTrue_1QNone_Bool_r)
        lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d <= lizzieLet30_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf;
  assign lizzieLet30_1MyTrue_1QNone_Bool_bufchan_r = (! lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf[0] ? lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf :
                                   lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        lizzieLet30_1MyTrue_1QNone_Bool_bufchan_buf <= lizzieLet30_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet30_1MyTrue_2,Go) > (lizzieLet30_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet30_1MyTrue_2_bufchan_d;
  logic lizzieLet30_1MyTrue_2_bufchan_r;
  assign lizzieLet30_1MyTrue_2_r = ((! lizzieLet30_1MyTrue_2_bufchan_d[0]) || lizzieLet30_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet30_1MyTrue_2_r)
        lizzieLet30_1MyTrue_2_bufchan_d <= lizzieLet30_1MyTrue_2_d;
  Go_t lizzieLet30_1MyTrue_2_bufchan_buf;
  assign lizzieLet30_1MyTrue_2_bufchan_r = (! lizzieLet30_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet30_1MyTrue_2_argbuf_d = (lizzieLet30_1MyTrue_2_bufchan_buf[0] ? lizzieLet30_1MyTrue_2_bufchan_buf :
                                           lizzieLet30_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet30_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet30_1MyTrue_2_argbuf_r && lizzieLet30_1MyTrue_2_bufchan_buf[0]))
        lizzieLet30_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet30_1MyTrue_2_argbuf_r) && (! lizzieLet30_1MyTrue_2_bufchan_buf[0])))
        lizzieLet30_1MyTrue_2_bufchan_buf <= lizzieLet30_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f) : (lizzieLet30_2,MyBool) (lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#,Pointer_CTf_f) > [(lizzieLet30_2MyFalse,Pointer_CTf_f),
                                                                                                             (lizzieLet30_2MyTrue,Pointer_CTf_f)] */
  logic [1:0] \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd ;
  always_comb
    if ((lizzieLet30_2_d[0] && \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_d [0]))
      unique case (lizzieLet30_2_d[1:1])
        1'd0: \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd  = 2'd1;
        1'd1: \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd  = 2'd2;
        default: \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd  = 2'd0;
      endcase
    else \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd  = 2'd0;
  assign lizzieLet30_2MyFalse_d = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_d [16:1],
                                   \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd [0]};
  assign lizzieLet30_2MyTrue_d = {\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_d [16:1],
                                  \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd [1]};
  assign \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_r  = (| (\lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_onehotd  & {lizzieLet30_2MyTrue_r,
                                                                                                                lizzieLet30_2MyFalse_r}));
  assign lizzieLet30_2_r = \lizzieLet12_4QVal_Int_5QVal_Int_5I#_4I#_r ;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet30_2MyFalse,Pointer_CTf_f) > (lizzieLet30_2MyFalse_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet30_2MyFalse_bufchan_d;
  logic lizzieLet30_2MyFalse_bufchan_r;
  assign lizzieLet30_2MyFalse_r = ((! lizzieLet30_2MyFalse_bufchan_d[0]) || lizzieLet30_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet30_2MyFalse_r)
        lizzieLet30_2MyFalse_bufchan_d <= lizzieLet30_2MyFalse_d;
  Pointer_CTf_f_t lizzieLet30_2MyFalse_bufchan_buf;
  assign lizzieLet30_2MyFalse_bufchan_r = (! lizzieLet30_2MyFalse_bufchan_buf[0]);
  assign lizzieLet30_2MyFalse_1_argbuf_d = (lizzieLet30_2MyFalse_bufchan_buf[0] ? lizzieLet30_2MyFalse_bufchan_buf :
                                            lizzieLet30_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet30_2MyFalse_1_argbuf_r && lizzieLet30_2MyFalse_bufchan_buf[0]))
        lizzieLet30_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet30_2MyFalse_1_argbuf_r) && (! lizzieLet30_2MyFalse_bufchan_buf[0])))
        lizzieLet30_2MyFalse_bufchan_buf <= lizzieLet30_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (lizzieLet30_2MyTrue,Pointer_CTf_f) > (lizzieLet30_2MyTrue_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t lizzieLet30_2MyTrue_bufchan_d;
  logic lizzieLet30_2MyTrue_bufchan_r;
  assign lizzieLet30_2MyTrue_r = ((! lizzieLet30_2MyTrue_bufchan_d[0]) || lizzieLet30_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet30_2MyTrue_r)
        lizzieLet30_2MyTrue_bufchan_d <= lizzieLet30_2MyTrue_d;
  Pointer_CTf_f_t lizzieLet30_2MyTrue_bufchan_buf;
  assign lizzieLet30_2MyTrue_bufchan_r = (! lizzieLet30_2MyTrue_bufchan_buf[0]);
  assign lizzieLet30_2MyTrue_1_argbuf_d = (lizzieLet30_2MyTrue_bufchan_buf[0] ? lizzieLet30_2MyTrue_bufchan_buf :
                                           lizzieLet30_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet30_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet30_2MyTrue_1_argbuf_r && lizzieLet30_2MyTrue_bufchan_buf[0]))
        lizzieLet30_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet30_2MyTrue_1_argbuf_r) && (! lizzieLet30_2MyTrue_bufchan_buf[0])))
        lizzieLet30_2MyTrue_bufchan_buf <= lizzieLet30_2MyTrue_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet3_1QNode_Int,QTree_Int) > [(tlae2_destruct,Pointer_QTree_Int),
                                                                 (trae3_destruct,Pointer_QTree_Int),
                                                                 (blae4_destruct,Pointer_QTree_Int),
                                                                 (brae5_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet3_1QNode_Int_emitted;
  logic [3:0] lizzieLet3_1QNode_Int_done;
  assign tlae2_destruct_d = {lizzieLet3_1QNode_Int_d[18:3],
                             (lizzieLet3_1QNode_Int_d[0] && (! lizzieLet3_1QNode_Int_emitted[0]))};
  assign trae3_destruct_d = {lizzieLet3_1QNode_Int_d[34:19],
                             (lizzieLet3_1QNode_Int_d[0] && (! lizzieLet3_1QNode_Int_emitted[1]))};
  assign blae4_destruct_d = {lizzieLet3_1QNode_Int_d[50:35],
                             (lizzieLet3_1QNode_Int_d[0] && (! lizzieLet3_1QNode_Int_emitted[2]))};
  assign brae5_destruct_d = {lizzieLet3_1QNode_Int_d[66:51],
                             (lizzieLet3_1QNode_Int_d[0] && (! lizzieLet3_1QNode_Int_emitted[3]))};
  assign lizzieLet3_1QNode_Int_done = (lizzieLet3_1QNode_Int_emitted | ({brae5_destruct_d[0],
                                                                         blae4_destruct_d[0],
                                                                         trae3_destruct_d[0],
                                                                         tlae2_destruct_d[0]} & {brae5_destruct_r,
                                                                                                 blae4_destruct_r,
                                                                                                 trae3_destruct_r,
                                                                                                 tlae2_destruct_r}));
  assign lizzieLet3_1QNode_Int_r = (& lizzieLet3_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet3_1QNode_Int_emitted <= (lizzieLet3_1QNode_Int_r ? 4'd0 :
                                        lizzieLet3_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet3_1QVal_Int,QTree_Int) > [(va8v_destruct,Int)] */
  assign va8v_destruct_d = {lizzieLet3_1QVal_Int_d[34:3],
                            lizzieLet3_1QVal_Int_d[0]};
  assign lizzieLet3_1QVal_Int_r = va8v_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet3_2,QTree_Int) (lizzieLet3_1,QTree_Int) > [(_7,QTree_Int),
                                                                            (lizzieLet3_1QVal_Int,QTree_Int),
                                                                            (lizzieLet3_1QNode_Int,QTree_Int),
                                                                            (_6,QTree_Int)] */
  logic [3:0] lizzieLet3_1_onehotd;
  always_comb
    if ((lizzieLet3_2_d[0] && lizzieLet3_1_d[0]))
      unique case (lizzieLet3_2_d[2:1])
        2'd0: lizzieLet3_1_onehotd = 4'd1;
        2'd1: lizzieLet3_1_onehotd = 4'd2;
        2'd2: lizzieLet3_1_onehotd = 4'd4;
        2'd3: lizzieLet3_1_onehotd = 4'd8;
        default: lizzieLet3_1_onehotd = 4'd0;
      endcase
    else lizzieLet3_1_onehotd = 4'd0;
  assign _7_d = {lizzieLet3_1_d[66:1], lizzieLet3_1_onehotd[0]};
  assign lizzieLet3_1QVal_Int_d = {lizzieLet3_1_d[66:1],
                                   lizzieLet3_1_onehotd[1]};
  assign lizzieLet3_1QNode_Int_d = {lizzieLet3_1_d[66:1],
                                    lizzieLet3_1_onehotd[2]};
  assign _6_d = {lizzieLet3_1_d[66:1], lizzieLet3_1_onehotd[3]};
  assign lizzieLet3_1_r = (| (lizzieLet3_1_onehotd & {_6_r,
                                                      lizzieLet3_1QNode_Int_r,
                                                      lizzieLet3_1QVal_Int_r,
                                                      _7_r}));
  assign lizzieLet3_2_r = lizzieLet3_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet3_3,QTree_Int) (go_14_goMux_data,Go) > [(lizzieLet3_3QNone_Int,Go),
                                                                  (lizzieLet3_3QVal_Int,Go),
                                                                  (lizzieLet3_3QNode_Int,Go),
                                                                  (lizzieLet3_3QError_Int,Go)] */
  logic [3:0] go_14_goMux_data_onehotd;
  always_comb
    if ((lizzieLet3_3_d[0] && go_14_goMux_data_d[0]))
      unique case (lizzieLet3_3_d[2:1])
        2'd0: go_14_goMux_data_onehotd = 4'd1;
        2'd1: go_14_goMux_data_onehotd = 4'd2;
        2'd2: go_14_goMux_data_onehotd = 4'd4;
        2'd3: go_14_goMux_data_onehotd = 4'd8;
        default: go_14_goMux_data_onehotd = 4'd0;
      endcase
    else go_14_goMux_data_onehotd = 4'd0;
  assign lizzieLet3_3QNone_Int_d = go_14_goMux_data_onehotd[0];
  assign lizzieLet3_3QVal_Int_d = go_14_goMux_data_onehotd[1];
  assign lizzieLet3_3QNode_Int_d = go_14_goMux_data_onehotd[2];
  assign lizzieLet3_3QError_Int_d = go_14_goMux_data_onehotd[3];
  assign go_14_goMux_data_r = (| (go_14_goMux_data_onehotd & {lizzieLet3_3QError_Int_r,
                                                              lizzieLet3_3QNode_Int_r,
                                                              lizzieLet3_3QVal_Int_r,
                                                              lizzieLet3_3QNone_Int_r}));
  assign lizzieLet3_3_r = go_14_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet3_3QError_Int,Go) > [(lizzieLet3_3QError_Int_1,Go),
                                              (lizzieLet3_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet3_3QError_Int_emitted;
  logic [1:0] lizzieLet3_3QError_Int_done;
  assign lizzieLet3_3QError_Int_1_d = (lizzieLet3_3QError_Int_d[0] && (! lizzieLet3_3QError_Int_emitted[0]));
  assign lizzieLet3_3QError_Int_2_d = (lizzieLet3_3QError_Int_d[0] && (! lizzieLet3_3QError_Int_emitted[1]));
  assign lizzieLet3_3QError_Int_done = (lizzieLet3_3QError_Int_emitted | ({lizzieLet3_3QError_Int_2_d[0],
                                                                           lizzieLet3_3QError_Int_1_d[0]} & {lizzieLet3_3QError_Int_2_r,
                                                                                                             lizzieLet3_3QError_Int_1_r}));
  assign lizzieLet3_3QError_Int_r = (& lizzieLet3_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet3_3QError_Int_emitted <= (lizzieLet3_3QError_Int_r ? 2'd0 :
                                         lizzieLet3_3QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet3_3QError_Int_1,Go)] > (lizzieLet3_3QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet3_3QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet3_3QError_Int_1_d[0]}), lizzieLet3_3QError_Int_1_d);
  assign {lizzieLet3_3QError_Int_1_r} = {1 {(lizzieLet3_3QError_Int_1QError_Bool_r && lizzieLet3_3QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet3_3QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet11_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet3_3QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet3_3QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet3_3QError_Int_1QError_Bool_r = ((! lizzieLet3_3QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet3_3QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_3QError_Int_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet3_3QError_Int_1QError_Bool_r)
        lizzieLet3_3QError_Int_1QError_Bool_bufchan_d <= lizzieLet3_3QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet3_3QError_Int_1QError_Bool_bufchan_r = (! lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet3_3QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet3_3QError_Int_1QError_Bool_bufchan_buf <= lizzieLet3_3QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet3_3QError_Int_2,Go) > (lizzieLet3_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet3_3QError_Int_2_bufchan_d;
  logic lizzieLet3_3QError_Int_2_bufchan_r;
  assign lizzieLet3_3QError_Int_2_r = ((! lizzieLet3_3QError_Int_2_bufchan_d[0]) || lizzieLet3_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet3_3QError_Int_2_r)
        lizzieLet3_3QError_Int_2_bufchan_d <= lizzieLet3_3QError_Int_2_d;
  Go_t lizzieLet3_3QError_Int_2_bufchan_buf;
  assign lizzieLet3_3QError_Int_2_bufchan_r = (! lizzieLet3_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet3_3QError_Int_2_argbuf_d = (lizzieLet3_3QError_Int_2_bufchan_buf[0] ? lizzieLet3_3QError_Int_2_bufchan_buf :
                                              lizzieLet3_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet3_3QError_Int_2_argbuf_r && lizzieLet3_3QError_Int_2_bufchan_buf[0]))
        lizzieLet3_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet3_3QError_Int_2_argbuf_r) && (! lizzieLet3_3QError_Int_2_bufchan_buf[0])))
        lizzieLet3_3QError_Int_2_bufchan_buf <= lizzieLet3_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet3_3QNode_Int,Go) > (lizzieLet3_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet3_3QNode_Int_bufchan_d;
  logic lizzieLet3_3QNode_Int_bufchan_r;
  assign lizzieLet3_3QNode_Int_r = ((! lizzieLet3_3QNode_Int_bufchan_d[0]) || lizzieLet3_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet3_3QNode_Int_r)
        lizzieLet3_3QNode_Int_bufchan_d <= lizzieLet3_3QNode_Int_d;
  Go_t lizzieLet3_3QNode_Int_bufchan_buf;
  assign lizzieLet3_3QNode_Int_bufchan_r = (! lizzieLet3_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet3_3QNode_Int_1_argbuf_d = (lizzieLet3_3QNode_Int_bufchan_buf[0] ? lizzieLet3_3QNode_Int_bufchan_buf :
                                             lizzieLet3_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet3_3QNode_Int_1_argbuf_r && lizzieLet3_3QNode_Int_bufchan_buf[0]))
        lizzieLet3_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet3_3QNode_Int_1_argbuf_r) && (! lizzieLet3_3QNode_Int_bufchan_buf[0])))
        lizzieLet3_3QNode_Int_bufchan_buf <= lizzieLet3_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet3_3QNone_Int,Go) > [(lizzieLet3_3QNone_Int_1,Go),
                                             (lizzieLet3_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet3_3QNone_Int_emitted;
  logic [1:0] lizzieLet3_3QNone_Int_done;
  assign lizzieLet3_3QNone_Int_1_d = (lizzieLet3_3QNone_Int_d[0] && (! lizzieLet3_3QNone_Int_emitted[0]));
  assign lizzieLet3_3QNone_Int_2_d = (lizzieLet3_3QNone_Int_d[0] && (! lizzieLet3_3QNone_Int_emitted[1]));
  assign lizzieLet3_3QNone_Int_done = (lizzieLet3_3QNone_Int_emitted | ({lizzieLet3_3QNone_Int_2_d[0],
                                                                         lizzieLet3_3QNone_Int_1_d[0]} & {lizzieLet3_3QNone_Int_2_r,
                                                                                                          lizzieLet3_3QNone_Int_1_r}));
  assign lizzieLet3_3QNone_Int_r = (& lizzieLet3_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet3_3QNone_Int_emitted <= (lizzieLet3_3QNone_Int_r ? 2'd0 :
                                        lizzieLet3_3QNone_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet3_3QNone_Int_1,Go)] > (lizzieLet3_3QNone_Int_1QNone_Bool,QTree_Bool) */
  assign lizzieLet3_3QNone_Int_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet3_3QNone_Int_1_d[0]}), lizzieLet3_3QNone_Int_1_d);
  assign {lizzieLet3_3QNone_Int_1_r} = {1 {(lizzieLet3_3QNone_Int_1QNone_Bool_r && lizzieLet3_3QNone_Int_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet3_3QNone_Int_1QNone_Bool,QTree_Bool) > (lizzieLet4_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d;
  logic lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_r;
  assign lizzieLet3_3QNone_Int_1QNone_Bool_r = ((! lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d[0]) || lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet3_3QNone_Int_1QNone_Bool_r)
        lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d <= lizzieLet3_3QNone_Int_1QNone_Bool_d;
  QTree_Bool_t lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf;
  assign lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_r = (! lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet4_1_argbuf_d = (lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf[0] ? lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf :
                                  lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf[0]))
        lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf[0])))
        lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_buf <= lizzieLet3_3QNone_Int_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet3_3QNone_Int_2,Go) > (lizzieLet3_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet3_3QNone_Int_2_bufchan_d;
  logic lizzieLet3_3QNone_Int_2_bufchan_r;
  assign lizzieLet3_3QNone_Int_2_r = ((! lizzieLet3_3QNone_Int_2_bufchan_d[0]) || lizzieLet3_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet3_3QNone_Int_2_r)
        lizzieLet3_3QNone_Int_2_bufchan_d <= lizzieLet3_3QNone_Int_2_d;
  Go_t lizzieLet3_3QNone_Int_2_bufchan_buf;
  assign lizzieLet3_3QNone_Int_2_bufchan_r = (! lizzieLet3_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet3_3QNone_Int_2_argbuf_d = (lizzieLet3_3QNone_Int_2_bufchan_buf[0] ? lizzieLet3_3QNone_Int_2_bufchan_buf :
                                             lizzieLet3_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet3_3QNone_Int_2_argbuf_r && lizzieLet3_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet3_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet3_3QNone_Int_2_argbuf_r) && (! lizzieLet3_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet3_3QNone_Int_2_bufchan_buf <= lizzieLet3_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet3_3QNone_Int_2_argbuf,Go),
                           (lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf,Go),
                           (lizzieLet7_1MyFalse_2_argbuf,Go),
                           (lizzieLet7_1MyTrue_2_argbuf,Go),
                           (lizzieLet3_3QError_Int_2_argbuf,Go)] > (go_20_goMux_choice,C5) (go_20_goMux_data,Go) */
  logic [4:0] lizzieLet3_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet3_3QNone_Int_2_argbuf_select_d = ((| lizzieLet3_3QNone_Int_2_argbuf_select_q) ? lizzieLet3_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet3_3QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                     (\lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_d [0] ? 5'd2 :
                                                      (lizzieLet7_1MyFalse_2_argbuf_d[0] ? 5'd4 :
                                                       (lizzieLet7_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                        (lizzieLet3_3QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                         5'd0))))));
  logic [4:0] lizzieLet3_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_3QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet3_3QNone_Int_2_argbuf_select_q <= (lizzieLet3_3QNone_Int_2_argbuf_done ? 5'd0 :
                                                  lizzieLet3_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet3_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet3_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet3_3QNone_Int_2_argbuf_emit_q <= (lizzieLet3_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet3_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet3_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet3_3QNone_Int_2_argbuf_emit_d = (lizzieLet3_3QNone_Int_2_argbuf_emit_q | ({go_20_goMux_choice_d[0],
                                                                                            go_20_goMux_data_d[0]} & {go_20_goMux_choice_r,
                                                                                                                      go_20_goMux_data_r}));
  logic lizzieLet3_3QNone_Int_2_argbuf_done;
  assign lizzieLet3_3QNone_Int_2_argbuf_done = (& lizzieLet3_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet3_3QError_Int_2_argbuf_r,
          lizzieLet7_1MyTrue_2_argbuf_r,
          lizzieLet7_1MyFalse_2_argbuf_r,
          \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_r ,
          lizzieLet3_3QNone_Int_2_argbuf_r} = (lizzieLet3_3QNone_Int_2_argbuf_done ? lizzieLet3_3QNone_Int_2_argbuf_select_d :
                                               5'd0);
  assign go_20_goMux_data_d = ((lizzieLet3_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet3_3QNone_Int_2_argbuf_d :
                               ((lizzieLet3_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_d  :
                                ((lizzieLet3_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet7_1MyFalse_2_argbuf_d :
                                 ((lizzieLet3_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet7_1MyTrue_2_argbuf_d :
                                  ((lizzieLet3_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet3_3QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_20_goMux_choice_d = ((lizzieLet3_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet3_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet3_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet3_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet3_3QNone_Int_2_argbuf_select_d[4] && (! lizzieLet3_3QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet3_4,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTf''''''''_f'''''''') > [(lizzieLet3_4QNone_Int,Pointer_CTf''''''''_f''''''''),
                                                                                                                        (lizzieLet3_4QVal_Int,Pointer_CTf''''''''_f''''''''),
                                                                                                                        (lizzieLet3_4QNode_Int,Pointer_CTf''''''''_f''''''''),
                                                                                                                        (lizzieLet3_4QError_Int,Pointer_CTf''''''''_f'''''''')] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet3_4_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet3_4_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet3_4QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet3_4QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet3_4QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet3_4QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet3_4QError_Int_r,
                                                              lizzieLet3_4QNode_Int_r,
                                                              lizzieLet3_4QVal_Int_r,
                                                              lizzieLet3_4QNone_Int_r}));
  assign lizzieLet3_4_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet3_4QError_Int,Pointer_CTf''''''''_f'''''''') > (lizzieLet3_4QError_Int_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QError_Int_bufchan_d;
  logic lizzieLet3_4QError_Int_bufchan_r;
  assign lizzieLet3_4QError_Int_r = ((! lizzieLet3_4QError_Int_bufchan_d[0]) || lizzieLet3_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet3_4QError_Int_r)
        lizzieLet3_4QError_Int_bufchan_d <= lizzieLet3_4QError_Int_d;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QError_Int_bufchan_buf;
  assign lizzieLet3_4QError_Int_bufchan_r = (! lizzieLet3_4QError_Int_bufchan_buf[0]);
  assign lizzieLet3_4QError_Int_1_argbuf_d = (lizzieLet3_4QError_Int_bufchan_buf[0] ? lizzieLet3_4QError_Int_bufchan_buf :
                                              lizzieLet3_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet3_4QError_Int_1_argbuf_r && lizzieLet3_4QError_Int_bufchan_buf[0]))
        lizzieLet3_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet3_4QError_Int_1_argbuf_r) && (! lizzieLet3_4QError_Int_bufchan_buf[0])))
        lizzieLet3_4QError_Int_bufchan_buf <= lizzieLet3_4QError_Int_bufchan_d;
  
  /* dcon (Ty CTf''''''''_f'''''''',
      Dcon Lcall_f''''''''_f''''''''3) : [(lizzieLet3_4QNode_Int,Pointer_CTf''''''''_f''''''''),
                                          (tlae2_destruct,Pointer_QTree_Int),
                                          (trae3_destruct,Pointer_QTree_Int),
                                          (blae4_destruct,Pointer_QTree_Int)] > (lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3,CTf''''''''_f'''''''') */
  assign \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_d  = \Lcall_f''''''''_f''''''''3_dc ((& {lizzieLet3_4QNode_Int_d[0],
                                                                                                                          tlae2_destruct_d[0],
                                                                                                                          trae3_destruct_d[0],
                                                                                                                          blae4_destruct_d[0]}), lizzieLet3_4QNode_Int_d, tlae2_destruct_d, trae3_destruct_d, blae4_destruct_d);
  assign {lizzieLet3_4QNode_Int_r,
          tlae2_destruct_r,
          trae3_destruct_r,
          blae4_destruct_r} = {4 {(\lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_r  && \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_d [0])}};
  
  /* buf (Ty CTf''''''''_f'''''''') : (lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3,CTf''''''''_f'''''''') > (lizzieLet10_1_argbuf,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d ;
  logic \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_r ;
  assign \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_r  = ((! \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d [0]) || \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d  <= {67'd0,
                                                                                             1'd0};
    else
      if (\lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_r )
        \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d  <= \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_d ;
  \CTf''''''''_f''''''''_t  \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf ;
  assign \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_r  = (! \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf [0]);
  assign lizzieLet10_1_argbuf_d = (\lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf [0] ? \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf  :
                                   \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf  <= {67'd0,
                                                                                               1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf [0]))
        \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf  <= {67'd0,
                                                                                                 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf [0])))
        \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_buf  <= \lizzieLet3_4QNode_Int_1tlae2_1trae3_1blae4_1Lcall_f''''''''_f''''''''3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet3_4QNone_Int,Pointer_CTf''''''''_f'''''''') > (lizzieLet3_4QNone_Int_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QNone_Int_bufchan_d;
  logic lizzieLet3_4QNone_Int_bufchan_r;
  assign lizzieLet3_4QNone_Int_r = ((! lizzieLet3_4QNone_Int_bufchan_d[0]) || lizzieLet3_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet3_4QNone_Int_r)
        lizzieLet3_4QNone_Int_bufchan_d <= lizzieLet3_4QNone_Int_d;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet3_4QNone_Int_bufchan_buf;
  assign lizzieLet3_4QNone_Int_bufchan_r = (! lizzieLet3_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet3_4QNone_Int_1_argbuf_d = (lizzieLet3_4QNone_Int_bufchan_buf[0] ? lizzieLet3_4QNone_Int_bufchan_buf :
                                             lizzieLet3_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet3_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet3_4QNone_Int_1_argbuf_r && lizzieLet3_4QNone_Int_bufchan_buf[0]))
        lizzieLet3_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet3_4QNone_Int_1_argbuf_r) && (! lizzieLet3_4QNone_Int_bufchan_buf[0])))
        lizzieLet3_4QNone_Int_bufchan_buf <= lizzieLet3_4QNone_Int_bufchan_d;
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz0) : (lizzieLet44_1Lcall_$wnnz0,CT$wnnz) > [(wwspI_4_destruct,Int#),
                                                                      (ww1Xqr_2_destruct,Int#),
                                                                      (ww2Xqu_1_destruct,Int#),
                                                                      (sc_0_6_destruct,Pointer_CT$wnnz)] */
  logic [3:0] lizzieLet44_1Lcall_$wnnz0_emitted;
  logic [3:0] lizzieLet44_1Lcall_$wnnz0_done;
  assign wwspI_4_destruct_d = {lizzieLet44_1Lcall_$wnnz0_d[35:4],
                               (lizzieLet44_1Lcall_$wnnz0_d[0] && (! lizzieLet44_1Lcall_$wnnz0_emitted[0]))};
  assign ww1Xqr_2_destruct_d = {lizzieLet44_1Lcall_$wnnz0_d[67:36],
                                (lizzieLet44_1Lcall_$wnnz0_d[0] && (! lizzieLet44_1Lcall_$wnnz0_emitted[1]))};
  assign ww2Xqu_1_destruct_d = {lizzieLet44_1Lcall_$wnnz0_d[99:68],
                                (lizzieLet44_1Lcall_$wnnz0_d[0] && (! lizzieLet44_1Lcall_$wnnz0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet44_1Lcall_$wnnz0_d[115:100],
                              (lizzieLet44_1Lcall_$wnnz0_d[0] && (! lizzieLet44_1Lcall_$wnnz0_emitted[3]))};
  assign lizzieLet44_1Lcall_$wnnz0_done = (lizzieLet44_1Lcall_$wnnz0_emitted | ({sc_0_6_destruct_d[0],
                                                                                 ww2Xqu_1_destruct_d[0],
                                                                                 ww1Xqr_2_destruct_d[0],
                                                                                 wwspI_4_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                           ww2Xqu_1_destruct_r,
                                                                                                           ww1Xqr_2_destruct_r,
                                                                                                           wwspI_4_destruct_r}));
  assign lizzieLet44_1Lcall_$wnnz0_r = (& lizzieLet44_1Lcall_$wnnz0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_1Lcall_$wnnz0_emitted <= 4'd0;
    else
      lizzieLet44_1Lcall_$wnnz0_emitted <= (lizzieLet44_1Lcall_$wnnz0_r ? 4'd0 :
                                            lizzieLet44_1Lcall_$wnnz0_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz1) : (lizzieLet44_1Lcall_$wnnz1,CT$wnnz) > [(wwspI_3_destruct,Int#),
                                                                      (ww1Xqr_1_destruct,Int#),
                                                                      (sc_0_5_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_3_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet44_1Lcall_$wnnz1_emitted;
  logic [3:0] lizzieLet44_1Lcall_$wnnz1_done;
  assign wwspI_3_destruct_d = {lizzieLet44_1Lcall_$wnnz1_d[35:4],
                               (lizzieLet44_1Lcall_$wnnz1_d[0] && (! lizzieLet44_1Lcall_$wnnz1_emitted[0]))};
  assign ww1Xqr_1_destruct_d = {lizzieLet44_1Lcall_$wnnz1_d[67:36],
                                (lizzieLet44_1Lcall_$wnnz1_d[0] && (! lizzieLet44_1Lcall_$wnnz1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet44_1Lcall_$wnnz1_d[83:68],
                              (lizzieLet44_1Lcall_$wnnz1_d[0] && (! lizzieLet44_1Lcall_$wnnz1_emitted[2]))};
  assign q4a87_3_destruct_d = {lizzieLet44_1Lcall_$wnnz1_d[99:84],
                               (lizzieLet44_1Lcall_$wnnz1_d[0] && (! lizzieLet44_1Lcall_$wnnz1_emitted[3]))};
  assign lizzieLet44_1Lcall_$wnnz1_done = (lizzieLet44_1Lcall_$wnnz1_emitted | ({q4a87_3_destruct_d[0],
                                                                                 sc_0_5_destruct_d[0],
                                                                                 ww1Xqr_1_destruct_d[0],
                                                                                 wwspI_3_destruct_d[0]} & {q4a87_3_destruct_r,
                                                                                                           sc_0_5_destruct_r,
                                                                                                           ww1Xqr_1_destruct_r,
                                                                                                           wwspI_3_destruct_r}));
  assign lizzieLet44_1Lcall_$wnnz1_r = (& lizzieLet44_1Lcall_$wnnz1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_1Lcall_$wnnz1_emitted <= 4'd0;
    else
      lizzieLet44_1Lcall_$wnnz1_emitted <= (lizzieLet44_1Lcall_$wnnz1_r ? 4'd0 :
                                            lizzieLet44_1Lcall_$wnnz1_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz2) : (lizzieLet44_1Lcall_$wnnz2,CT$wnnz) > [(wwspI_2_destruct,Int#),
                                                                      (sc_0_4_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_2_destruct,Pointer_QTree_Bool),
                                                                      (q3a86_2_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet44_1Lcall_$wnnz2_emitted;
  logic [3:0] lizzieLet44_1Lcall_$wnnz2_done;
  assign wwspI_2_destruct_d = {lizzieLet44_1Lcall_$wnnz2_d[35:4],
                               (lizzieLet44_1Lcall_$wnnz2_d[0] && (! lizzieLet44_1Lcall_$wnnz2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet44_1Lcall_$wnnz2_d[51:36],
                              (lizzieLet44_1Lcall_$wnnz2_d[0] && (! lizzieLet44_1Lcall_$wnnz2_emitted[1]))};
  assign q4a87_2_destruct_d = {lizzieLet44_1Lcall_$wnnz2_d[67:52],
                               (lizzieLet44_1Lcall_$wnnz2_d[0] && (! lizzieLet44_1Lcall_$wnnz2_emitted[2]))};
  assign q3a86_2_destruct_d = {lizzieLet44_1Lcall_$wnnz2_d[83:68],
                               (lizzieLet44_1Lcall_$wnnz2_d[0] && (! lizzieLet44_1Lcall_$wnnz2_emitted[3]))};
  assign lizzieLet44_1Lcall_$wnnz2_done = (lizzieLet44_1Lcall_$wnnz2_emitted | ({q3a86_2_destruct_d[0],
                                                                                 q4a87_2_destruct_d[0],
                                                                                 sc_0_4_destruct_d[0],
                                                                                 wwspI_2_destruct_d[0]} & {q3a86_2_destruct_r,
                                                                                                           q4a87_2_destruct_r,
                                                                                                           sc_0_4_destruct_r,
                                                                                                           wwspI_2_destruct_r}));
  assign lizzieLet44_1Lcall_$wnnz2_r = (& lizzieLet44_1Lcall_$wnnz2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_1Lcall_$wnnz2_emitted <= 4'd0;
    else
      lizzieLet44_1Lcall_$wnnz2_emitted <= (lizzieLet44_1Lcall_$wnnz2_r ? 4'd0 :
                                            lizzieLet44_1Lcall_$wnnz2_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz3) : (lizzieLet44_1Lcall_$wnnz3,CT$wnnz) > [(sc_0_3_destruct,Pointer_CT$wnnz),
                                                                      (q4a87_1_destruct,Pointer_QTree_Bool),
                                                                      (q3a86_1_destruct,Pointer_QTree_Bool),
                                                                      (q2a85_1_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet44_1Lcall_$wnnz3_emitted;
  logic [3:0] lizzieLet44_1Lcall_$wnnz3_done;
  assign sc_0_3_destruct_d = {lizzieLet44_1Lcall_$wnnz3_d[19:4],
                              (lizzieLet44_1Lcall_$wnnz3_d[0] && (! lizzieLet44_1Lcall_$wnnz3_emitted[0]))};
  assign q4a87_1_destruct_d = {lizzieLet44_1Lcall_$wnnz3_d[35:20],
                               (lizzieLet44_1Lcall_$wnnz3_d[0] && (! lizzieLet44_1Lcall_$wnnz3_emitted[1]))};
  assign q3a86_1_destruct_d = {lizzieLet44_1Lcall_$wnnz3_d[51:36],
                               (lizzieLet44_1Lcall_$wnnz3_d[0] && (! lizzieLet44_1Lcall_$wnnz3_emitted[2]))};
  assign q2a85_1_destruct_d = {lizzieLet44_1Lcall_$wnnz3_d[67:52],
                               (lizzieLet44_1Lcall_$wnnz3_d[0] && (! lizzieLet44_1Lcall_$wnnz3_emitted[3]))};
  assign lizzieLet44_1Lcall_$wnnz3_done = (lizzieLet44_1Lcall_$wnnz3_emitted | ({q2a85_1_destruct_d[0],
                                                                                 q3a86_1_destruct_d[0],
                                                                                 q4a87_1_destruct_d[0],
                                                                                 sc_0_3_destruct_d[0]} & {q2a85_1_destruct_r,
                                                                                                          q3a86_1_destruct_r,
                                                                                                          q4a87_1_destruct_r,
                                                                                                          sc_0_3_destruct_r}));
  assign lizzieLet44_1Lcall_$wnnz3_r = (& lizzieLet44_1Lcall_$wnnz3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_1Lcall_$wnnz3_emitted <= 4'd0;
    else
      lizzieLet44_1Lcall_$wnnz3_emitted <= (lizzieLet44_1Lcall_$wnnz3_r ? 4'd0 :
                                            lizzieLet44_1Lcall_$wnnz3_done);
  
  /* demux (Ty CT$wnnz,
       Ty CT$wnnz) : (lizzieLet44_2,CT$wnnz) (lizzieLet44_1,CT$wnnz) > [(_5,CT$wnnz),
                                                                        (lizzieLet44_1Lcall_$wnnz3,CT$wnnz),
                                                                        (lizzieLet44_1Lcall_$wnnz2,CT$wnnz),
                                                                        (lizzieLet44_1Lcall_$wnnz1,CT$wnnz),
                                                                        (lizzieLet44_1Lcall_$wnnz0,CT$wnnz)] */
  logic [4:0] lizzieLet44_1_onehotd;
  always_comb
    if ((lizzieLet44_2_d[0] && lizzieLet44_1_d[0]))
      unique case (lizzieLet44_2_d[3:1])
        3'd0: lizzieLet44_1_onehotd = 5'd1;
        3'd1: lizzieLet44_1_onehotd = 5'd2;
        3'd2: lizzieLet44_1_onehotd = 5'd4;
        3'd3: lizzieLet44_1_onehotd = 5'd8;
        3'd4: lizzieLet44_1_onehotd = 5'd16;
        default: lizzieLet44_1_onehotd = 5'd0;
      endcase
    else lizzieLet44_1_onehotd = 5'd0;
  assign _5_d = {lizzieLet44_1_d[115:1], lizzieLet44_1_onehotd[0]};
  assign lizzieLet44_1Lcall_$wnnz3_d = {lizzieLet44_1_d[115:1],
                                        lizzieLet44_1_onehotd[1]};
  assign lizzieLet44_1Lcall_$wnnz2_d = {lizzieLet44_1_d[115:1],
                                        lizzieLet44_1_onehotd[2]};
  assign lizzieLet44_1Lcall_$wnnz1_d = {lizzieLet44_1_d[115:1],
                                        lizzieLet44_1_onehotd[3]};
  assign lizzieLet44_1Lcall_$wnnz0_d = {lizzieLet44_1_d[115:1],
                                        lizzieLet44_1_onehotd[4]};
  assign lizzieLet44_1_r = (| (lizzieLet44_1_onehotd & {lizzieLet44_1Lcall_$wnnz0_r,
                                                        lizzieLet44_1Lcall_$wnnz1_r,
                                                        lizzieLet44_1Lcall_$wnnz2_r,
                                                        lizzieLet44_1Lcall_$wnnz3_r,
                                                        _5_r}));
  assign lizzieLet44_2_r = lizzieLet44_1_r;
  
  /* demux (Ty CT$wnnz,
       Ty Go) : (lizzieLet44_3,CT$wnnz) (go_19_goMux_data,Go) > [(_4,Go),
                                                                 (lizzieLet44_3Lcall_$wnnz3,Go),
                                                                 (lizzieLet44_3Lcall_$wnnz2,Go),
                                                                 (lizzieLet44_3Lcall_$wnnz1,Go),
                                                                 (lizzieLet44_3Lcall_$wnnz0,Go)] */
  logic [4:0] go_19_goMux_data_onehotd;
  always_comb
    if ((lizzieLet44_3_d[0] && go_19_goMux_data_d[0]))
      unique case (lizzieLet44_3_d[3:1])
        3'd0: go_19_goMux_data_onehotd = 5'd1;
        3'd1: go_19_goMux_data_onehotd = 5'd2;
        3'd2: go_19_goMux_data_onehotd = 5'd4;
        3'd3: go_19_goMux_data_onehotd = 5'd8;
        3'd4: go_19_goMux_data_onehotd = 5'd16;
        default: go_19_goMux_data_onehotd = 5'd0;
      endcase
    else go_19_goMux_data_onehotd = 5'd0;
  assign _4_d = go_19_goMux_data_onehotd[0];
  assign lizzieLet44_3Lcall_$wnnz3_d = go_19_goMux_data_onehotd[1];
  assign lizzieLet44_3Lcall_$wnnz2_d = go_19_goMux_data_onehotd[2];
  assign lizzieLet44_3Lcall_$wnnz1_d = go_19_goMux_data_onehotd[3];
  assign lizzieLet44_3Lcall_$wnnz0_d = go_19_goMux_data_onehotd[4];
  assign go_19_goMux_data_r = (| (go_19_goMux_data_onehotd & {lizzieLet44_3Lcall_$wnnz0_r,
                                                              lizzieLet44_3Lcall_$wnnz1_r,
                                                              lizzieLet44_3Lcall_$wnnz2_r,
                                                              lizzieLet44_3Lcall_$wnnz3_r,
                                                              _4_r}));
  assign lizzieLet44_3_r = go_19_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_$wnnz0,Go) > (lizzieLet44_3Lcall_$wnnz0_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_$wnnz0_bufchan_d;
  logic lizzieLet44_3Lcall_$wnnz0_bufchan_r;
  assign lizzieLet44_3Lcall_$wnnz0_r = ((! lizzieLet44_3Lcall_$wnnz0_bufchan_d[0]) || lizzieLet44_3Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz0_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_$wnnz0_r)
        lizzieLet44_3Lcall_$wnnz0_bufchan_d <= lizzieLet44_3Lcall_$wnnz0_d;
  Go_t lizzieLet44_3Lcall_$wnnz0_bufchan_buf;
  assign lizzieLet44_3Lcall_$wnnz0_bufchan_r = (! lizzieLet44_3Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_$wnnz0_1_argbuf_d = (lizzieLet44_3Lcall_$wnnz0_bufchan_buf[0] ? lizzieLet44_3Lcall_$wnnz0_bufchan_buf :
                                                 lizzieLet44_3Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_$wnnz0_1_argbuf_r && lizzieLet44_3Lcall_$wnnz0_bufchan_buf[0]))
        lizzieLet44_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_$wnnz0_1_argbuf_r) && (! lizzieLet44_3Lcall_$wnnz0_bufchan_buf[0])))
        lizzieLet44_3Lcall_$wnnz0_bufchan_buf <= lizzieLet44_3Lcall_$wnnz0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_$wnnz1,Go) > (lizzieLet44_3Lcall_$wnnz1_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_$wnnz1_bufchan_d;
  logic lizzieLet44_3Lcall_$wnnz1_bufchan_r;
  assign lizzieLet44_3Lcall_$wnnz1_r = ((! lizzieLet44_3Lcall_$wnnz1_bufchan_d[0]) || lizzieLet44_3Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz1_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_$wnnz1_r)
        lizzieLet44_3Lcall_$wnnz1_bufchan_d <= lizzieLet44_3Lcall_$wnnz1_d;
  Go_t lizzieLet44_3Lcall_$wnnz1_bufchan_buf;
  assign lizzieLet44_3Lcall_$wnnz1_bufchan_r = (! lizzieLet44_3Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_$wnnz1_1_argbuf_d = (lizzieLet44_3Lcall_$wnnz1_bufchan_buf[0] ? lizzieLet44_3Lcall_$wnnz1_bufchan_buf :
                                                 lizzieLet44_3Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_$wnnz1_1_argbuf_r && lizzieLet44_3Lcall_$wnnz1_bufchan_buf[0]))
        lizzieLet44_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_$wnnz1_1_argbuf_r) && (! lizzieLet44_3Lcall_$wnnz1_bufchan_buf[0])))
        lizzieLet44_3Lcall_$wnnz1_bufchan_buf <= lizzieLet44_3Lcall_$wnnz1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_$wnnz2,Go) > (lizzieLet44_3Lcall_$wnnz2_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_$wnnz2_bufchan_d;
  logic lizzieLet44_3Lcall_$wnnz2_bufchan_r;
  assign lizzieLet44_3Lcall_$wnnz2_r = ((! lizzieLet44_3Lcall_$wnnz2_bufchan_d[0]) || lizzieLet44_3Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz2_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_$wnnz2_r)
        lizzieLet44_3Lcall_$wnnz2_bufchan_d <= lizzieLet44_3Lcall_$wnnz2_d;
  Go_t lizzieLet44_3Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet44_3Lcall_$wnnz2_bufchan_r = (! lizzieLet44_3Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_$wnnz2_1_argbuf_d = (lizzieLet44_3Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet44_3Lcall_$wnnz2_bufchan_buf :
                                                 lizzieLet44_3Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_$wnnz2_1_argbuf_r && lizzieLet44_3Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet44_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_$wnnz2_1_argbuf_r) && (! lizzieLet44_3Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet44_3Lcall_$wnnz2_bufchan_buf <= lizzieLet44_3Lcall_$wnnz2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet44_3Lcall_$wnnz3,Go) > (lizzieLet44_3Lcall_$wnnz3_1_argbuf,Go) */
  Go_t lizzieLet44_3Lcall_$wnnz3_bufchan_d;
  logic lizzieLet44_3Lcall_$wnnz3_bufchan_r;
  assign lizzieLet44_3Lcall_$wnnz3_r = ((! lizzieLet44_3Lcall_$wnnz3_bufchan_d[0]) || lizzieLet44_3Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz3_bufchan_d <= 1'd0;
    else
      if (lizzieLet44_3Lcall_$wnnz3_r)
        lizzieLet44_3Lcall_$wnnz3_bufchan_d <= lizzieLet44_3Lcall_$wnnz3_d;
  Go_t lizzieLet44_3Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet44_3Lcall_$wnnz3_bufchan_r = (! lizzieLet44_3Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet44_3Lcall_$wnnz3_1_argbuf_d = (lizzieLet44_3Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet44_3Lcall_$wnnz3_bufchan_buf :
                                                 lizzieLet44_3Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet44_3Lcall_$wnnz3_1_argbuf_r && lizzieLet44_3Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet44_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet44_3Lcall_$wnnz3_1_argbuf_r) && (! lizzieLet44_3Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet44_3Lcall_$wnnz3_bufchan_buf <= lizzieLet44_3Lcall_$wnnz3_bufchan_d;
  
  /* demux (Ty CT$wnnz,
       Ty Int#) : (lizzieLet44_4,CT$wnnz) (srtarg_0_goMux_mux,Int#) > [(lizzieLet44_4L$wnnzsbos,Int#),
                                                                       (lizzieLet44_4Lcall_$wnnz3,Int#),
                                                                       (lizzieLet44_4Lcall_$wnnz2,Int#),
                                                                       (lizzieLet44_4Lcall_$wnnz1,Int#),
                                                                       (lizzieLet44_4Lcall_$wnnz0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet44_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet44_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet44_4L$wnnzsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                      srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet44_4Lcall_$wnnz3_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet44_4Lcall_$wnnz2_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet44_4Lcall_$wnnz1_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet44_4Lcall_$wnnz0_d = {srtarg_0_goMux_mux_d[32:1],
                                        srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet44_4Lcall_$wnnz0_r,
                                                                  lizzieLet44_4Lcall_$wnnz1_r,
                                                                  lizzieLet44_4Lcall_$wnnz2_r,
                                                                  lizzieLet44_4Lcall_$wnnz3_r,
                                                                  lizzieLet44_4L$wnnzsbos_r}));
  assign lizzieLet44_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet44_4L$wnnzsbos,Int#) > [(lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1,Int#),
                                                   (lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet44_4L$wnnzsbos_emitted;
  logic [1:0] lizzieLet44_4L$wnnzsbos_done;
  assign lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_d = {lizzieLet44_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet44_4L$wnnzsbos_d[0] && (! lizzieLet44_4L$wnnzsbos_emitted[0]))};
  assign lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_d = {lizzieLet44_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet44_4L$wnnzsbos_d[0] && (! lizzieLet44_4L$wnnzsbos_emitted[1]))};
  assign lizzieLet44_4L$wnnzsbos_done = (lizzieLet44_4L$wnnzsbos_emitted | ({lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_d[0],
                                                                             lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_r,
                                                                                                                                   lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet44_4L$wnnzsbos_r = (& lizzieLet44_4L$wnnzsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet44_4L$wnnzsbos_emitted <= 2'd0;
    else
      lizzieLet44_4L$wnnzsbos_emitted <= (lizzieLet44_4L$wnnzsbos_r ? 2'd0 :
                                          lizzieLet44_4L$wnnzsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_goConst,Go) */
  assign call_$wnnz_goConst_d = lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_1_r = call_$wnnz_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2,Int#) > ($wnnz_resbuf,Int#) */
  \Int#_t  lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_r = ((! lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_r)
        lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_resbuf_d  = (lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf :
                             lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((\$wnnz_resbuf_r  && lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! \$wnnz_resbuf_r ) && (! lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet44_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz2) : [(lizzieLet44_4Lcall_$wnnz3,Int#),
                            (sc_0_3_destruct,Pointer_CT$wnnz),
                            (q4a87_1_destruct,Pointer_QTree_Bool),
                            (q3a86_1_destruct,Pointer_QTree_Bool)] > (lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2,CT$wnnz) */
  assign lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d = Lcall_$wnnz2_dc((& {lizzieLet44_4Lcall_$wnnz3_d[0],
                                                                                                   sc_0_3_destruct_d[0],
                                                                                                   q4a87_1_destruct_d[0],
                                                                                                   q3a86_1_destruct_d[0]}), lizzieLet44_4Lcall_$wnnz3_d, sc_0_3_destruct_d, q4a87_1_destruct_d, q3a86_1_destruct_d);
  assign {lizzieLet44_4Lcall_$wnnz3_r,
          sc_0_3_destruct_r,
          q4a87_1_destruct_r,
          q3a86_1_destruct_r} = {4 {(lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r && lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2,CT$wnnz) > (lizzieLet45_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d;
  logic lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r;
  assign lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r = ((! lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d[0]) || lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_r)
        lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d <= lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_d;
  CT$wnnz_t lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_r = (! lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet45_1_argbuf_d = (lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf :
                                   lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet45_1_argbuf_r && lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet45_1_argbuf_r) && (! lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_buf <= lizzieLet44_4Lcall_$wnnz3_1sc_0_3_1q4a87_1_1q3a86_1_1Lcall_$wnnz2_bufchan_d;
  
  /* destruct (Ty CTf''''''''_f'''''''',
          Dcon Lcall_f''''''''_f''''''''0) : (lizzieLet48_1Lcall_f''''''''_f''''''''0,CTf''''''''_f'''''''') > [(es_1_2_destruct,Pointer_QTree_Bool),
                                                                                                                (es_2_2_destruct,Pointer_QTree_Bool),
                                                                                                                (es_3_3_destruct,Pointer_QTree_Bool),
                                                                                                                (sc_0_10_destruct,Pointer_CTf''''''''_f'''''''')] */
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted ;
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''0_done ;
  assign es_1_2_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [19:4],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted [0]))};
  assign es_2_2_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [35:20],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted [1]))};
  assign es_3_3_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [51:36],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [67:52],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''0_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted [3]))};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''0_done  = (\lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted  | ({sc_0_10_destruct_d[0],
                                                                                                                 es_3_3_destruct_d[0],
                                                                                                                 es_2_2_destruct_d[0],
                                                                                                                 es_1_2_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                                          es_3_3_destruct_r,
                                                                                                                                          es_2_2_destruct_r,
                                                                                                                                          es_1_2_destruct_r}));
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''0_r  = (& \lizzieLet48_1Lcall_f''''''''_f''''''''0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted  <= 4'd0;
    else
      \lizzieLet48_1Lcall_f''''''''_f''''''''0_emitted  <= (\lizzieLet48_1Lcall_f''''''''_f''''''''0_r  ? 4'd0 :
                                                            \lizzieLet48_1Lcall_f''''''''_f''''''''0_done );
  
  /* destruct (Ty CTf''''''''_f'''''''',
          Dcon Lcall_f''''''''_f''''''''1) : (lizzieLet48_1Lcall_f''''''''_f''''''''1,CTf''''''''_f'''''''') > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                                                                                (es_3_2_destruct,Pointer_QTree_Bool),
                                                                                                                (sc_0_9_destruct,Pointer_CTf''''''''_f''''''''),
                                                                                                                (tlae2_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted ;
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''1_done ;
  assign es_2_1_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [19:4],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted [0]))};
  assign es_3_2_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [35:20],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [51:36],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted [2]))};
  assign tlae2_3_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [67:52],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''1_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted [3]))};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''1_done  = (\lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted  | ({tlae2_3_destruct_d[0],
                                                                                                                 sc_0_9_destruct_d[0],
                                                                                                                 es_3_2_destruct_d[0],
                                                                                                                 es_2_1_destruct_d[0]} & {tlae2_3_destruct_r,
                                                                                                                                          sc_0_9_destruct_r,
                                                                                                                                          es_3_2_destruct_r,
                                                                                                                                          es_2_1_destruct_r}));
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''1_r  = (& \lizzieLet48_1Lcall_f''''''''_f''''''''1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted  <= 4'd0;
    else
      \lizzieLet48_1Lcall_f''''''''_f''''''''1_emitted  <= (\lizzieLet48_1Lcall_f''''''''_f''''''''1_r  ? 4'd0 :
                                                            \lizzieLet48_1Lcall_f''''''''_f''''''''1_done );
  
  /* destruct (Ty CTf''''''''_f'''''''',
          Dcon Lcall_f''''''''_f''''''''2) : (lizzieLet48_1Lcall_f''''''''_f''''''''2,CTf''''''''_f'''''''') > [(es_3_1_destruct,Pointer_QTree_Bool),
                                                                                                                (sc_0_8_destruct,Pointer_CTf''''''''_f''''''''),
                                                                                                                (tlae2_2_destruct,Pointer_QTree_Int),
                                                                                                                (trae3_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted ;
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''2_done ;
  assign es_3_1_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [19:4],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [35:20],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted [1]))};
  assign tlae2_2_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [51:36],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted [2]))};
  assign trae3_2_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [67:52],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''2_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted [3]))};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''2_done  = (\lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted  | ({trae3_2_destruct_d[0],
                                                                                                                 tlae2_2_destruct_d[0],
                                                                                                                 sc_0_8_destruct_d[0],
                                                                                                                 es_3_1_destruct_d[0]} & {trae3_2_destruct_r,
                                                                                                                                          tlae2_2_destruct_r,
                                                                                                                                          sc_0_8_destruct_r,
                                                                                                                                          es_3_1_destruct_r}));
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''2_r  = (& \lizzieLet48_1Lcall_f''''''''_f''''''''2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted  <= 4'd0;
    else
      \lizzieLet48_1Lcall_f''''''''_f''''''''2_emitted  <= (\lizzieLet48_1Lcall_f''''''''_f''''''''2_r  ? 4'd0 :
                                                            \lizzieLet48_1Lcall_f''''''''_f''''''''2_done );
  
  /* destruct (Ty CTf''''''''_f'''''''',
          Dcon Lcall_f''''''''_f''''''''3) : (lizzieLet48_1Lcall_f''''''''_f''''''''3,CTf''''''''_f'''''''') > [(sc_0_7_destruct,Pointer_CTf''''''''_f''''''''),
                                                                                                                (tlae2_1_destruct,Pointer_QTree_Int),
                                                                                                                (trae3_1_destruct,Pointer_QTree_Int),
                                                                                                                (blae4_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted ;
  logic [3:0] \lizzieLet48_1Lcall_f''''''''_f''''''''3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [19:4],
                              (\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted [0]))};
  assign tlae2_1_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [35:20],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted [1]))};
  assign trae3_1_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [51:36],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted [2]))};
  assign blae4_1_destruct_d = {\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [67:52],
                               (\lizzieLet48_1Lcall_f''''''''_f''''''''3_d [0] && (! \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted [3]))};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''3_done  = (\lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted  | ({blae4_1_destruct_d[0],
                                                                                                                 trae3_1_destruct_d[0],
                                                                                                                 tlae2_1_destruct_d[0],
                                                                                                                 sc_0_7_destruct_d[0]} & {blae4_1_destruct_r,
                                                                                                                                          trae3_1_destruct_r,
                                                                                                                                          tlae2_1_destruct_r,
                                                                                                                                          sc_0_7_destruct_r}));
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''3_r  = (& \lizzieLet48_1Lcall_f''''''''_f''''''''3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted  <= 4'd0;
    else
      \lizzieLet48_1Lcall_f''''''''_f''''''''3_emitted  <= (\lizzieLet48_1Lcall_f''''''''_f''''''''3_r  ? 4'd0 :
                                                            \lizzieLet48_1Lcall_f''''''''_f''''''''3_done );
  
  /* demux (Ty CTf''''''''_f'''''''',
       Ty CTf''''''''_f'''''''') : (lizzieLet48_2,CTf''''''''_f'''''''') (lizzieLet48_1,CTf''''''''_f'''''''') > [(_3,CTf''''''''_f''''''''),
                                                                                                                  (lizzieLet48_1Lcall_f''''''''_f''''''''3,CTf''''''''_f''''''''),
                                                                                                                  (lizzieLet48_1Lcall_f''''''''_f''''''''2,CTf''''''''_f''''''''),
                                                                                                                  (lizzieLet48_1Lcall_f''''''''_f''''''''1,CTf''''''''_f''''''''),
                                                                                                                  (lizzieLet48_1Lcall_f''''''''_f''''''''0,CTf''''''''_f'''''''')] */
  logic [4:0] lizzieLet48_1_onehotd;
  always_comb
    if ((lizzieLet48_2_d[0] && lizzieLet48_1_d[0]))
      unique case (lizzieLet48_2_d[3:1])
        3'd0: lizzieLet48_1_onehotd = 5'd1;
        3'd1: lizzieLet48_1_onehotd = 5'd2;
        3'd2: lizzieLet48_1_onehotd = 5'd4;
        3'd3: lizzieLet48_1_onehotd = 5'd8;
        3'd4: lizzieLet48_1_onehotd = 5'd16;
        default: lizzieLet48_1_onehotd = 5'd0;
      endcase
    else lizzieLet48_1_onehotd = 5'd0;
  assign _3_d = {lizzieLet48_1_d[67:1], lizzieLet48_1_onehotd[0]};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''3_d  = {lizzieLet48_1_d[67:1],
                                                        lizzieLet48_1_onehotd[1]};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''2_d  = {lizzieLet48_1_d[67:1],
                                                        lizzieLet48_1_onehotd[2]};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''1_d  = {lizzieLet48_1_d[67:1],
                                                        lizzieLet48_1_onehotd[3]};
  assign \lizzieLet48_1Lcall_f''''''''_f''''''''0_d  = {lizzieLet48_1_d[67:1],
                                                        lizzieLet48_1_onehotd[4]};
  assign lizzieLet48_1_r = (| (lizzieLet48_1_onehotd & {\lizzieLet48_1Lcall_f''''''''_f''''''''0_r ,
                                                        \lizzieLet48_1Lcall_f''''''''_f''''''''1_r ,
                                                        \lizzieLet48_1Lcall_f''''''''_f''''''''2_r ,
                                                        \lizzieLet48_1Lcall_f''''''''_f''''''''3_r ,
                                                        _3_r}));
  assign lizzieLet48_2_r = lizzieLet48_1_r;
  
  /* demux (Ty CTf''''''''_f'''''''',
       Ty Go) : (lizzieLet48_3,CTf''''''''_f'''''''') (go_20_goMux_data,Go) > [(_2,Go),
                                                                               (lizzieLet48_3Lcall_f''''''''_f''''''''3,Go),
                                                                               (lizzieLet48_3Lcall_f''''''''_f''''''''2,Go),
                                                                               (lizzieLet48_3Lcall_f''''''''_f''''''''1,Go),
                                                                               (lizzieLet48_3Lcall_f''''''''_f''''''''0,Go)] */
  logic [4:0] go_20_goMux_data_onehotd;
  always_comb
    if ((lizzieLet48_3_d[0] && go_20_goMux_data_d[0]))
      unique case (lizzieLet48_3_d[3:1])
        3'd0: go_20_goMux_data_onehotd = 5'd1;
        3'd1: go_20_goMux_data_onehotd = 5'd2;
        3'd2: go_20_goMux_data_onehotd = 5'd4;
        3'd3: go_20_goMux_data_onehotd = 5'd8;
        3'd4: go_20_goMux_data_onehotd = 5'd16;
        default: go_20_goMux_data_onehotd = 5'd0;
      endcase
    else go_20_goMux_data_onehotd = 5'd0;
  assign _2_d = go_20_goMux_data_onehotd[0];
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''3_d  = go_20_goMux_data_onehotd[1];
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''2_d  = go_20_goMux_data_onehotd[2];
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''1_d  = go_20_goMux_data_onehotd[3];
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''0_d  = go_20_goMux_data_onehotd[4];
  assign go_20_goMux_data_r = (| (go_20_goMux_data_onehotd & {\lizzieLet48_3Lcall_f''''''''_f''''''''0_r ,
                                                              \lizzieLet48_3Lcall_f''''''''_f''''''''1_r ,
                                                              \lizzieLet48_3Lcall_f''''''''_f''''''''2_r ,
                                                              \lizzieLet48_3Lcall_f''''''''_f''''''''3_r ,
                                                              _2_r}));
  assign lizzieLet48_3_r = go_20_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f''''''''_f''''''''0,Go) > (lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_r ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''0_r  = ((! \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d [0]) || \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f''''''''_f''''''''0_r )
        \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d  <= \lizzieLet48_3Lcall_f''''''''_f''''''''0_d ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_r  = (! \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_d  = (\lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf [0] ? \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf  :
                                                                 \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_r  && \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f''''''''_f''''''''0_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_buf  <= \lizzieLet48_3Lcall_f''''''''_f''''''''0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f''''''''_f''''''''1,Go) > (lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_r ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''1_r  = ((! \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d [0]) || \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f''''''''_f''''''''1_r )
        \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d  <= \lizzieLet48_3Lcall_f''''''''_f''''''''1_d ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_r  = (! \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_d  = (\lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf [0] ? \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf  :
                                                                 \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_r  && \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f''''''''_f''''''''1_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_buf  <= \lizzieLet48_3Lcall_f''''''''_f''''''''1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f''''''''_f''''''''2,Go) > (lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_r ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''2_r  = ((! \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d [0]) || \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f''''''''_f''''''''2_r )
        \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d  <= \lizzieLet48_3Lcall_f''''''''_f''''''''2_d ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_r  = (! \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_d  = (\lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf [0] ? \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf  :
                                                                 \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_r  && \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f''''''''_f''''''''2_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_buf  <= \lizzieLet48_3Lcall_f''''''''_f''''''''2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet48_3Lcall_f''''''''_f''''''''3,Go) > (lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf,Go) */
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d ;
  logic \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_r ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''3_r  = ((! \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d [0]) || \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet48_3Lcall_f''''''''_f''''''''3_r )
        \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d  <= \lizzieLet48_3Lcall_f''''''''_f''''''''3_d ;
  Go_t \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf ;
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_r  = (! \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf [0]);
  assign \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_d  = (\lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf [0] ? \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf  :
                                                                 \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_r  && \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf [0]))
        \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet48_3Lcall_f''''''''_f''''''''3_1_argbuf_r ) && (! \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf [0])))
        \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_buf  <= \lizzieLet48_3Lcall_f''''''''_f''''''''3_bufchan_d ;
  
  /* demux (Ty CTf''''''''_f'''''''',
       Ty Pointer_QTree_Bool) : (lizzieLet48_4,CTf''''''''_f'''''''') (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet48_4Lf''''''''_f''''''''sbos,Pointer_QTree_Bool),
                                                                                                                   (lizzieLet48_4Lcall_f''''''''_f''''''''3,Pointer_QTree_Bool),
                                                                                                                   (lizzieLet48_4Lcall_f''''''''_f''''''''2,Pointer_QTree_Bool),
                                                                                                                   (lizzieLet48_4Lcall_f''''''''_f''''''''1,Pointer_QTree_Bool),
                                                                                                                   (lizzieLet48_4Lcall_f''''''''_f''''''''0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet48_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet48_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                      srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet48_4Lcall_f''''''''_f''''''''0_r ,
                                                                      \lizzieLet48_4Lcall_f''''''''_f''''''''1_r ,
                                                                      \lizzieLet48_4Lcall_f''''''''_f''''''''2_r ,
                                                                      \lizzieLet48_4Lcall_f''''''''_f''''''''3_r ,
                                                                      \lizzieLet48_4Lf''''''''_f''''''''sbos_r }));
  assign lizzieLet48_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet48_4Lcall_f''''''''_f''''''''0,Pointer_QTree_Bool),
                          (es_1_2_destruct,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_3_destruct,Pointer_QTree_Bool)] > (lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet48_4Lcall_f''''''''_f''''''''0_d [0],
                                                                                                             es_1_2_destruct_d[0],
                                                                                                             es_2_2_destruct_d[0],
                                                                                                             es_3_3_destruct_d[0]}), \lizzieLet48_4Lcall_f''''''''_f''''''''0_d , es_1_2_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {\lizzieLet48_4Lcall_f''''''''_f''''''''0_r ,
          es_1_2_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(\lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r  && \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) > (lizzieLet52_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r  = ((! \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d [0]) || \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                                  1'd0};
    else
      if (\lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r )
        \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d  <= \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r  = (! \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet52_1_argbuf_d = (\lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0] ? \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                    1'd0};
    else
      if ((lizzieLet52_1_argbuf_r && \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                      1'd0};
      else if (((! lizzieLet52_1_argbuf_r) && (! \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf  <= \lizzieLet48_4Lcall_f''''''''_f''''''''0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f'''''''',
      Dcon Lcall_f''''''''_f''''''''0) : [(lizzieLet48_4Lcall_f''''''''_f''''''''1,Pointer_QTree_Bool),
                                          (es_2_1_destruct,Pointer_QTree_Bool),
                                          (es_3_2_destruct,Pointer_QTree_Bool),
                                          (sc_0_9_destruct,Pointer_CTf''''''''_f'''''''')] > (lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0,CTf''''''''_f'''''''') */
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_d  = \Lcall_f''''''''_f''''''''0_dc ((& {\lizzieLet48_4Lcall_f''''''''_f''''''''1_d [0],
                                                                                                                                               es_2_1_destruct_d[0],
                                                                                                                                               es_3_2_destruct_d[0],
                                                                                                                                               sc_0_9_destruct_d[0]}), \lizzieLet48_4Lcall_f''''''''_f''''''''1_d , es_2_1_destruct_d, es_3_2_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet48_4Lcall_f''''''''_f''''''''1_r ,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_r  && \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_d [0])}};
  
  /* buf (Ty CTf''''''''_f'''''''') : (lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0,CTf''''''''_f'''''''') > (lizzieLet51_1_argbuf,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_r ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_r  = ((! \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d [0]) || \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d  <= {67'd0,
                                                                                                                  1'd0};
    else
      if (\lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_r )
        \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d  <= \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_d ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_r  = (! \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf [0]);
  assign lizzieLet51_1_argbuf_d = (\lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf [0] ? \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf  <= {67'd0,
                                                                                                                    1'd0};
    else
      if ((lizzieLet51_1_argbuf_r && \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf  <= {67'd0,
                                                                                                                      1'd0};
      else if (((! lizzieLet51_1_argbuf_r) && (! \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_buf  <= \lizzieLet48_4Lcall_f''''''''_f''''''''1_1es_2_1_1es_3_2_1sc_0_9_1Lcall_f''''''''_f''''''''0_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f'''''''',
      Dcon Lcall_f''''''''_f''''''''1) : [(lizzieLet48_4Lcall_f''''''''_f''''''''2,Pointer_QTree_Bool),
                                          (es_3_1_destruct,Pointer_QTree_Bool),
                                          (sc_0_8_destruct,Pointer_CTf''''''''_f''''''''),
                                          (tlae2_2_destruct,Pointer_QTree_Int)] > (lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1,CTf''''''''_f'''''''') */
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_d  = \Lcall_f''''''''_f''''''''1_dc ((& {\lizzieLet48_4Lcall_f''''''''_f''''''''2_d [0],
                                                                                                                                                es_3_1_destruct_d[0],
                                                                                                                                                sc_0_8_destruct_d[0],
                                                                                                                                                tlae2_2_destruct_d[0]}), \lizzieLet48_4Lcall_f''''''''_f''''''''2_d , es_3_1_destruct_d, sc_0_8_destruct_d, tlae2_2_destruct_d);
  assign {\lizzieLet48_4Lcall_f''''''''_f''''''''2_r ,
          es_3_1_destruct_r,
          sc_0_8_destruct_r,
          tlae2_2_destruct_r} = {4 {(\lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_r  && \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_d [0])}};
  
  /* buf (Ty CTf''''''''_f'''''''') : (lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1,CTf''''''''_f'''''''') > (lizzieLet50_1_argbuf,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_r ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_r  = ((! \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d [0]) || \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d  <= {67'd0,
                                                                                                                   1'd0};
    else
      if (\lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_r )
        \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d  <= \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_d ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_r  = (! \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf [0]);
  assign lizzieLet50_1_argbuf_d = (\lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf [0] ? \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf  <= {67'd0,
                                                                                                                     1'd0};
    else
      if ((lizzieLet50_1_argbuf_r && \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf  <= {67'd0,
                                                                                                                       1'd0};
      else if (((! lizzieLet50_1_argbuf_r) && (! \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_buf  <= \lizzieLet48_4Lcall_f''''''''_f''''''''2_1es_3_1_1sc_0_8_1tlae2_2_1Lcall_f''''''''_f''''''''1_bufchan_d ;
  
  /* dcon (Ty CTf''''''''_f'''''''',
      Dcon Lcall_f''''''''_f''''''''2) : [(lizzieLet48_4Lcall_f''''''''_f''''''''3,Pointer_QTree_Bool),
                                          (sc_0_7_destruct,Pointer_CTf''''''''_f''''''''),
                                          (tlae2_1_destruct,Pointer_QTree_Int),
                                          (trae3_1_destruct,Pointer_QTree_Int)] > (lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2,CTf''''''''_f'''''''') */
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_d  = \Lcall_f''''''''_f''''''''2_dc ((& {\lizzieLet48_4Lcall_f''''''''_f''''''''3_d [0],
                                                                                                                                                 sc_0_7_destruct_d[0],
                                                                                                                                                 tlae2_1_destruct_d[0],
                                                                                                                                                 trae3_1_destruct_d[0]}), \lizzieLet48_4Lcall_f''''''''_f''''''''3_d , sc_0_7_destruct_d, tlae2_1_destruct_d, trae3_1_destruct_d);
  assign {\lizzieLet48_4Lcall_f''''''''_f''''''''3_r ,
          sc_0_7_destruct_r,
          tlae2_1_destruct_r,
          trae3_1_destruct_r} = {4 {(\lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_r  && \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_d [0])}};
  
  /* buf (Ty CTf''''''''_f'''''''') : (lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2,CTf''''''''_f'''''''') > (lizzieLet49_1_argbuf,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d ;
  logic \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_r ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_r  = ((! \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d [0]) || \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d  <= {67'd0,
                                                                                                                    1'd0};
    else
      if (\lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_r )
        \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d  <= \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_d ;
  \CTf''''''''_f''''''''_t  \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf ;
  assign \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_r  = (! \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf [0]);
  assign lizzieLet49_1_argbuf_d = (\lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf [0] ? \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf  :
                                   \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf  <= {67'd0,
                                                                                                                      1'd0};
    else
      if ((lizzieLet49_1_argbuf_r && \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf [0]))
        \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf  <= {67'd0,
                                                                                                                        1'd0};
      else if (((! lizzieLet49_1_argbuf_r) && (! \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf [0])))
        \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_buf  <= \lizzieLet48_4Lcall_f''''''''_f''''''''3_1sc_0_7_1tlae2_1_1trae3_1_1Lcall_f''''''''_f''''''''2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet48_4Lf''''''''_f''''''''sbos,Pointer_QTree_Bool) > [(lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                             (lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet48_4Lf''''''''_f''''''''sbos_emitted ;
  logic [1:0] \lizzieLet48_4Lf''''''''_f''''''''sbos_done ;
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_d [16:1],
                                                                           (\lizzieLet48_4Lf''''''''_f''''''''sbos_d [0] && (! \lizzieLet48_4Lf''''''''_f''''''''sbos_emitted [0]))};
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d  = {\lizzieLet48_4Lf''''''''_f''''''''sbos_d [16:1],
                                                                           (\lizzieLet48_4Lf''''''''_f''''''''sbos_d [0] && (! \lizzieLet48_4Lf''''''''_f''''''''sbos_emitted [1]))};
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_done  = (\lizzieLet48_4Lf''''''''_f''''''''sbos_emitted  | ({\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_d [0],
                                                                                                             \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                   \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_r  = (& \lizzieLet48_4Lf''''''''_f''''''''sbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet48_4Lf''''''''_f''''''''sbos_emitted  <= 2'd0;
    else
      \lizzieLet48_4Lf''''''''_f''''''''sbos_emitted  <= (\lizzieLet48_4Lf''''''''_f''''''''sbos_r  ? 2'd0 :
                                                          \lizzieLet48_4Lf''''''''_f''''''''sbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f''''''''_f''''''''_goConst,Go) */
  assign \call_f''''''''_f''''''''_goConst_d  = \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet48_4Lf''''''''_f''''''''sbos_1_merge_merge_fork_1_r  = \call_f''''''''_f''''''''_goConst_r ;
  
  /* destruct (Ty CTf_f,
          Dcon Lcall_f_f0) : (lizzieLet53_1Lcall_f_f0,CTf_f) > [(es_10_destruct,Pointer_QTree_Bool),
                                                                (es_11_1_destruct,Pointer_QTree_Bool),
                                                                (es_12_2_destruct,Pointer_QTree_Bool),
                                                                (sc_0_14_destruct,Pointer_CTf_f)] */
  logic [3:0] lizzieLet53_1Lcall_f_f0_emitted;
  logic [3:0] lizzieLet53_1Lcall_f_f0_done;
  assign es_10_destruct_d = {lizzieLet53_1Lcall_f_f0_d[19:4],
                             (lizzieLet53_1Lcall_f_f0_d[0] && (! lizzieLet53_1Lcall_f_f0_emitted[0]))};
  assign es_11_1_destruct_d = {lizzieLet53_1Lcall_f_f0_d[35:20],
                               (lizzieLet53_1Lcall_f_f0_d[0] && (! lizzieLet53_1Lcall_f_f0_emitted[1]))};
  assign es_12_2_destruct_d = {lizzieLet53_1Lcall_f_f0_d[51:36],
                               (lizzieLet53_1Lcall_f_f0_d[0] && (! lizzieLet53_1Lcall_f_f0_emitted[2]))};
  assign sc_0_14_destruct_d = {lizzieLet53_1Lcall_f_f0_d[67:52],
                               (lizzieLet53_1Lcall_f_f0_d[0] && (! lizzieLet53_1Lcall_f_f0_emitted[3]))};
  assign lizzieLet53_1Lcall_f_f0_done = (lizzieLet53_1Lcall_f_f0_emitted | ({sc_0_14_destruct_d[0],
                                                                             es_12_2_destruct_d[0],
                                                                             es_11_1_destruct_d[0],
                                                                             es_10_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                     es_12_2_destruct_r,
                                                                                                     es_11_1_destruct_r,
                                                                                                     es_10_destruct_r}));
  assign lizzieLet53_1Lcall_f_f0_r = (& lizzieLet53_1Lcall_f_f0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_1Lcall_f_f0_emitted <= 4'd0;
    else
      lizzieLet53_1Lcall_f_f0_emitted <= (lizzieLet53_1Lcall_f_f0_r ? 4'd0 :
                                          lizzieLet53_1Lcall_f_f0_done);
  
  /* destruct (Ty CTf_f,
          Dcon Lcall_f_f1) : (lizzieLet53_1Lcall_f_f1,CTf_f) > [(es_11_destruct,Pointer_QTree_Bool),
                                                                (es_12_1_destruct,Pointer_QTree_Bool),
                                                                (sc_0_13_destruct,Pointer_CTf_f),
                                                                (q1aen_3_destruct,Pointer_QTree_Int),
                                                                (t1aes_3_destruct,Pointer_QTree_Int)] */
  logic [4:0] lizzieLet53_1Lcall_f_f1_emitted;
  logic [4:0] lizzieLet53_1Lcall_f_f1_done;
  assign es_11_destruct_d = {lizzieLet53_1Lcall_f_f1_d[19:4],
                             (lizzieLet53_1Lcall_f_f1_d[0] && (! lizzieLet53_1Lcall_f_f1_emitted[0]))};
  assign es_12_1_destruct_d = {lizzieLet53_1Lcall_f_f1_d[35:20],
                               (lizzieLet53_1Lcall_f_f1_d[0] && (! lizzieLet53_1Lcall_f_f1_emitted[1]))};
  assign sc_0_13_destruct_d = {lizzieLet53_1Lcall_f_f1_d[51:36],
                               (lizzieLet53_1Lcall_f_f1_d[0] && (! lizzieLet53_1Lcall_f_f1_emitted[2]))};
  assign q1aen_3_destruct_d = {lizzieLet53_1Lcall_f_f1_d[67:52],
                               (lizzieLet53_1Lcall_f_f1_d[0] && (! lizzieLet53_1Lcall_f_f1_emitted[3]))};
  assign t1aes_3_destruct_d = {lizzieLet53_1Lcall_f_f1_d[83:68],
                               (lizzieLet53_1Lcall_f_f1_d[0] && (! lizzieLet53_1Lcall_f_f1_emitted[4]))};
  assign lizzieLet53_1Lcall_f_f1_done = (lizzieLet53_1Lcall_f_f1_emitted | ({t1aes_3_destruct_d[0],
                                                                             q1aen_3_destruct_d[0],
                                                                             sc_0_13_destruct_d[0],
                                                                             es_12_1_destruct_d[0],
                                                                             es_11_destruct_d[0]} & {t1aes_3_destruct_r,
                                                                                                     q1aen_3_destruct_r,
                                                                                                     sc_0_13_destruct_r,
                                                                                                     es_12_1_destruct_r,
                                                                                                     es_11_destruct_r}));
  assign lizzieLet53_1Lcall_f_f1_r = (& lizzieLet53_1Lcall_f_f1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_1Lcall_f_f1_emitted <= 5'd0;
    else
      lizzieLet53_1Lcall_f_f1_emitted <= (lizzieLet53_1Lcall_f_f1_r ? 5'd0 :
                                          lizzieLet53_1Lcall_f_f1_done);
  
  /* destruct (Ty CTf_f,
          Dcon Lcall_f_f2) : (lizzieLet53_1Lcall_f_f2,CTf_f) > [(es_12_destruct,Pointer_QTree_Bool),
                                                                (sc_0_12_destruct,Pointer_CTf_f),
                                                                (q1aen_2_destruct,Pointer_QTree_Int),
                                                                (t1aes_2_destruct,Pointer_QTree_Int),
                                                                (q2aeo_2_destruct,Pointer_QTree_Int),
                                                                (t2aet_2_destruct,Pointer_QTree_Int)] */
  logic [5:0] lizzieLet53_1Lcall_f_f2_emitted;
  logic [5:0] lizzieLet53_1Lcall_f_f2_done;
  assign es_12_destruct_d = {lizzieLet53_1Lcall_f_f2_d[19:4],
                             (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[0]))};
  assign sc_0_12_destruct_d = {lizzieLet53_1Lcall_f_f2_d[35:20],
                               (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[1]))};
  assign q1aen_2_destruct_d = {lizzieLet53_1Lcall_f_f2_d[51:36],
                               (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[2]))};
  assign t1aes_2_destruct_d = {lizzieLet53_1Lcall_f_f2_d[67:52],
                               (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[3]))};
  assign q2aeo_2_destruct_d = {lizzieLet53_1Lcall_f_f2_d[83:68],
                               (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[4]))};
  assign t2aet_2_destruct_d = {lizzieLet53_1Lcall_f_f2_d[99:84],
                               (lizzieLet53_1Lcall_f_f2_d[0] && (! lizzieLet53_1Lcall_f_f2_emitted[5]))};
  assign lizzieLet53_1Lcall_f_f2_done = (lizzieLet53_1Lcall_f_f2_emitted | ({t2aet_2_destruct_d[0],
                                                                             q2aeo_2_destruct_d[0],
                                                                             t1aes_2_destruct_d[0],
                                                                             q1aen_2_destruct_d[0],
                                                                             sc_0_12_destruct_d[0],
                                                                             es_12_destruct_d[0]} & {t2aet_2_destruct_r,
                                                                                                     q2aeo_2_destruct_r,
                                                                                                     t1aes_2_destruct_r,
                                                                                                     q1aen_2_destruct_r,
                                                                                                     sc_0_12_destruct_r,
                                                                                                     es_12_destruct_r}));
  assign lizzieLet53_1Lcall_f_f2_r = (& lizzieLet53_1Lcall_f_f2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_1Lcall_f_f2_emitted <= 6'd0;
    else
      lizzieLet53_1Lcall_f_f2_emitted <= (lizzieLet53_1Lcall_f_f2_r ? 6'd0 :
                                          lizzieLet53_1Lcall_f_f2_done);
  
  /* destruct (Ty CTf_f,
          Dcon Lcall_f_f3) : (lizzieLet53_1Lcall_f_f3,CTf_f) > [(sc_0_11_destruct,Pointer_CTf_f),
                                                                (q1aen_1_destruct,Pointer_QTree_Int),
                                                                (t1aes_1_destruct,Pointer_QTree_Int),
                                                                (q2aeo_1_destruct,Pointer_QTree_Int),
                                                                (t2aet_1_destruct,Pointer_QTree_Int),
                                                                (q3aep_1_destruct,Pointer_QTree_Int),
                                                                (t3aeu_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet53_1Lcall_f_f3_emitted;
  logic [6:0] lizzieLet53_1Lcall_f_f3_done;
  assign sc_0_11_destruct_d = {lizzieLet53_1Lcall_f_f3_d[19:4],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[0]))};
  assign q1aen_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[35:20],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[1]))};
  assign t1aes_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[51:36],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[2]))};
  assign q2aeo_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[67:52],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[3]))};
  assign t2aet_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[83:68],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[4]))};
  assign q3aep_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[99:84],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[5]))};
  assign t3aeu_1_destruct_d = {lizzieLet53_1Lcall_f_f3_d[115:100],
                               (lizzieLet53_1Lcall_f_f3_d[0] && (! lizzieLet53_1Lcall_f_f3_emitted[6]))};
  assign lizzieLet53_1Lcall_f_f3_done = (lizzieLet53_1Lcall_f_f3_emitted | ({t3aeu_1_destruct_d[0],
                                                                             q3aep_1_destruct_d[0],
                                                                             t2aet_1_destruct_d[0],
                                                                             q2aeo_1_destruct_d[0],
                                                                             t1aes_1_destruct_d[0],
                                                                             q1aen_1_destruct_d[0],
                                                                             sc_0_11_destruct_d[0]} & {t3aeu_1_destruct_r,
                                                                                                       q3aep_1_destruct_r,
                                                                                                       t2aet_1_destruct_r,
                                                                                                       q2aeo_1_destruct_r,
                                                                                                       t1aes_1_destruct_r,
                                                                                                       q1aen_1_destruct_r,
                                                                                                       sc_0_11_destruct_r}));
  assign lizzieLet53_1Lcall_f_f3_r = (& lizzieLet53_1Lcall_f_f3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_1Lcall_f_f3_emitted <= 7'd0;
    else
      lizzieLet53_1Lcall_f_f3_emitted <= (lizzieLet53_1Lcall_f_f3_r ? 7'd0 :
                                          lizzieLet53_1Lcall_f_f3_done);
  
  /* demux (Ty CTf_f,
       Ty CTf_f) : (lizzieLet53_2,CTf_f) (lizzieLet53_1,CTf_f) > [(_1,CTf_f),
                                                                  (lizzieLet53_1Lcall_f_f3,CTf_f),
                                                                  (lizzieLet53_1Lcall_f_f2,CTf_f),
                                                                  (lizzieLet53_1Lcall_f_f1,CTf_f),
                                                                  (lizzieLet53_1Lcall_f_f0,CTf_f)] */
  logic [4:0] lizzieLet53_1_onehotd;
  always_comb
    if ((lizzieLet53_2_d[0] && lizzieLet53_1_d[0]))
      unique case (lizzieLet53_2_d[3:1])
        3'd0: lizzieLet53_1_onehotd = 5'd1;
        3'd1: lizzieLet53_1_onehotd = 5'd2;
        3'd2: lizzieLet53_1_onehotd = 5'd4;
        3'd3: lizzieLet53_1_onehotd = 5'd8;
        3'd4: lizzieLet53_1_onehotd = 5'd16;
        default: lizzieLet53_1_onehotd = 5'd0;
      endcase
    else lizzieLet53_1_onehotd = 5'd0;
  assign _1_d = {lizzieLet53_1_d[115:1], lizzieLet53_1_onehotd[0]};
  assign lizzieLet53_1Lcall_f_f3_d = {lizzieLet53_1_d[115:1],
                                      lizzieLet53_1_onehotd[1]};
  assign lizzieLet53_1Lcall_f_f2_d = {lizzieLet53_1_d[115:1],
                                      lizzieLet53_1_onehotd[2]};
  assign lizzieLet53_1Lcall_f_f1_d = {lizzieLet53_1_d[115:1],
                                      lizzieLet53_1_onehotd[3]};
  assign lizzieLet53_1Lcall_f_f0_d = {lizzieLet53_1_d[115:1],
                                      lizzieLet53_1_onehotd[4]};
  assign lizzieLet53_1_r = (| (lizzieLet53_1_onehotd & {lizzieLet53_1Lcall_f_f0_r,
                                                        lizzieLet53_1Lcall_f_f1_r,
                                                        lizzieLet53_1Lcall_f_f2_r,
                                                        lizzieLet53_1Lcall_f_f3_r,
                                                        _1_r}));
  assign lizzieLet53_2_r = lizzieLet53_1_r;
  
  /* demux (Ty CTf_f,
       Ty Go) : (lizzieLet53_3,CTf_f) (go_21_goMux_data,Go) > [(_0,Go),
                                                               (lizzieLet53_3Lcall_f_f3,Go),
                                                               (lizzieLet53_3Lcall_f_f2,Go),
                                                               (lizzieLet53_3Lcall_f_f1,Go),
                                                               (lizzieLet53_3Lcall_f_f0,Go)] */
  logic [4:0] go_21_goMux_data_onehotd;
  always_comb
    if ((lizzieLet53_3_d[0] && go_21_goMux_data_d[0]))
      unique case (lizzieLet53_3_d[3:1])
        3'd0: go_21_goMux_data_onehotd = 5'd1;
        3'd1: go_21_goMux_data_onehotd = 5'd2;
        3'd2: go_21_goMux_data_onehotd = 5'd4;
        3'd3: go_21_goMux_data_onehotd = 5'd8;
        3'd4: go_21_goMux_data_onehotd = 5'd16;
        default: go_21_goMux_data_onehotd = 5'd0;
      endcase
    else go_21_goMux_data_onehotd = 5'd0;
  assign _0_d = go_21_goMux_data_onehotd[0];
  assign lizzieLet53_3Lcall_f_f3_d = go_21_goMux_data_onehotd[1];
  assign lizzieLet53_3Lcall_f_f2_d = go_21_goMux_data_onehotd[2];
  assign lizzieLet53_3Lcall_f_f1_d = go_21_goMux_data_onehotd[3];
  assign lizzieLet53_3Lcall_f_f0_d = go_21_goMux_data_onehotd[4];
  assign go_21_goMux_data_r = (| (go_21_goMux_data_onehotd & {lizzieLet53_3Lcall_f_f0_r,
                                                              lizzieLet53_3Lcall_f_f1_r,
                                                              lizzieLet53_3Lcall_f_f2_r,
                                                              lizzieLet53_3Lcall_f_f3_r,
                                                              _0_r}));
  assign lizzieLet53_3_r = go_21_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f_f0,Go) > (lizzieLet53_3Lcall_f_f0_1_argbuf,Go) */
  Go_t lizzieLet53_3Lcall_f_f0_bufchan_d;
  logic lizzieLet53_3Lcall_f_f0_bufchan_r;
  assign lizzieLet53_3Lcall_f_f0_r = ((! lizzieLet53_3Lcall_f_f0_bufchan_d[0]) || lizzieLet53_3Lcall_f_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f0_bufchan_d <= 1'd0;
    else
      if (lizzieLet53_3Lcall_f_f0_r)
        lizzieLet53_3Lcall_f_f0_bufchan_d <= lizzieLet53_3Lcall_f_f0_d;
  Go_t lizzieLet53_3Lcall_f_f0_bufchan_buf;
  assign lizzieLet53_3Lcall_f_f0_bufchan_r = (! lizzieLet53_3Lcall_f_f0_bufchan_buf[0]);
  assign lizzieLet53_3Lcall_f_f0_1_argbuf_d = (lizzieLet53_3Lcall_f_f0_bufchan_buf[0] ? lizzieLet53_3Lcall_f_f0_bufchan_buf :
                                               lizzieLet53_3Lcall_f_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet53_3Lcall_f_f0_1_argbuf_r && lizzieLet53_3Lcall_f_f0_bufchan_buf[0]))
        lizzieLet53_3Lcall_f_f0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet53_3Lcall_f_f0_1_argbuf_r) && (! lizzieLet53_3Lcall_f_f0_bufchan_buf[0])))
        lizzieLet53_3Lcall_f_f0_bufchan_buf <= lizzieLet53_3Lcall_f_f0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f_f1,Go) > (lizzieLet53_3Lcall_f_f1_1_argbuf,Go) */
  Go_t lizzieLet53_3Lcall_f_f1_bufchan_d;
  logic lizzieLet53_3Lcall_f_f1_bufchan_r;
  assign lizzieLet53_3Lcall_f_f1_r = ((! lizzieLet53_3Lcall_f_f1_bufchan_d[0]) || lizzieLet53_3Lcall_f_f1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f1_bufchan_d <= 1'd0;
    else
      if (lizzieLet53_3Lcall_f_f1_r)
        lizzieLet53_3Lcall_f_f1_bufchan_d <= lizzieLet53_3Lcall_f_f1_d;
  Go_t lizzieLet53_3Lcall_f_f1_bufchan_buf;
  assign lizzieLet53_3Lcall_f_f1_bufchan_r = (! lizzieLet53_3Lcall_f_f1_bufchan_buf[0]);
  assign lizzieLet53_3Lcall_f_f1_1_argbuf_d = (lizzieLet53_3Lcall_f_f1_bufchan_buf[0] ? lizzieLet53_3Lcall_f_f1_bufchan_buf :
                                               lizzieLet53_3Lcall_f_f1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet53_3Lcall_f_f1_1_argbuf_r && lizzieLet53_3Lcall_f_f1_bufchan_buf[0]))
        lizzieLet53_3Lcall_f_f1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet53_3Lcall_f_f1_1_argbuf_r) && (! lizzieLet53_3Lcall_f_f1_bufchan_buf[0])))
        lizzieLet53_3Lcall_f_f1_bufchan_buf <= lizzieLet53_3Lcall_f_f1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f_f2,Go) > (lizzieLet53_3Lcall_f_f2_1_argbuf,Go) */
  Go_t lizzieLet53_3Lcall_f_f2_bufchan_d;
  logic lizzieLet53_3Lcall_f_f2_bufchan_r;
  assign lizzieLet53_3Lcall_f_f2_r = ((! lizzieLet53_3Lcall_f_f2_bufchan_d[0]) || lizzieLet53_3Lcall_f_f2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f2_bufchan_d <= 1'd0;
    else
      if (lizzieLet53_3Lcall_f_f2_r)
        lizzieLet53_3Lcall_f_f2_bufchan_d <= lizzieLet53_3Lcall_f_f2_d;
  Go_t lizzieLet53_3Lcall_f_f2_bufchan_buf;
  assign lizzieLet53_3Lcall_f_f2_bufchan_r = (! lizzieLet53_3Lcall_f_f2_bufchan_buf[0]);
  assign lizzieLet53_3Lcall_f_f2_1_argbuf_d = (lizzieLet53_3Lcall_f_f2_bufchan_buf[0] ? lizzieLet53_3Lcall_f_f2_bufchan_buf :
                                               lizzieLet53_3Lcall_f_f2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet53_3Lcall_f_f2_1_argbuf_r && lizzieLet53_3Lcall_f_f2_bufchan_buf[0]))
        lizzieLet53_3Lcall_f_f2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet53_3Lcall_f_f2_1_argbuf_r) && (! lizzieLet53_3Lcall_f_f2_bufchan_buf[0])))
        lizzieLet53_3Lcall_f_f2_bufchan_buf <= lizzieLet53_3Lcall_f_f2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet53_3Lcall_f_f3,Go) > (lizzieLet53_3Lcall_f_f3_1_argbuf,Go) */
  Go_t lizzieLet53_3Lcall_f_f3_bufchan_d;
  logic lizzieLet53_3Lcall_f_f3_bufchan_r;
  assign lizzieLet53_3Lcall_f_f3_r = ((! lizzieLet53_3Lcall_f_f3_bufchan_d[0]) || lizzieLet53_3Lcall_f_f3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f3_bufchan_d <= 1'd0;
    else
      if (lizzieLet53_3Lcall_f_f3_r)
        lizzieLet53_3Lcall_f_f3_bufchan_d <= lizzieLet53_3Lcall_f_f3_d;
  Go_t lizzieLet53_3Lcall_f_f3_bufchan_buf;
  assign lizzieLet53_3Lcall_f_f3_bufchan_r = (! lizzieLet53_3Lcall_f_f3_bufchan_buf[0]);
  assign lizzieLet53_3Lcall_f_f3_1_argbuf_d = (lizzieLet53_3Lcall_f_f3_bufchan_buf[0] ? lizzieLet53_3Lcall_f_f3_bufchan_buf :
                                               lizzieLet53_3Lcall_f_f3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_3Lcall_f_f3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet53_3Lcall_f_f3_1_argbuf_r && lizzieLet53_3Lcall_f_f3_bufchan_buf[0]))
        lizzieLet53_3Lcall_f_f3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet53_3Lcall_f_f3_1_argbuf_r) && (! lizzieLet53_3Lcall_f_f3_bufchan_buf[0])))
        lizzieLet53_3Lcall_f_f3_bufchan_buf <= lizzieLet53_3Lcall_f_f3_bufchan_d;
  
  /* demux (Ty CTf_f,
       Ty Pointer_QTree_Bool) : (lizzieLet53_4,CTf_f) (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet53_4Lf_fsbos,Pointer_QTree_Bool),
                                                                                                   (lizzieLet53_4Lcall_f_f3,Pointer_QTree_Bool),
                                                                                                   (lizzieLet53_4Lcall_f_f2,Pointer_QTree_Bool),
                                                                                                   (lizzieLet53_4Lcall_f_f1,Pointer_QTree_Bool),
                                                                                                   (lizzieLet53_4Lcall_f_f0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet53_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet53_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet53_4Lf_fsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                    srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet53_4Lcall_f_f3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                      srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet53_4Lcall_f_f2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                      srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet53_4Lcall_f_f1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                      srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet53_4Lcall_f_f0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                      srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet53_4Lcall_f_f0_r,
                                                                      lizzieLet53_4Lcall_f_f1_r,
                                                                      lizzieLet53_4Lcall_f_f2_r,
                                                                      lizzieLet53_4Lcall_f_f3_r,
                                                                      lizzieLet53_4Lf_fsbos_r}));
  assign lizzieLet53_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet53_4Lcall_f_f0,Pointer_QTree_Bool),
                          (es_10_destruct,Pointer_QTree_Bool),
                          (es_11_1_destruct,Pointer_QTree_Bool),
                          (es_12_2_destruct,Pointer_QTree_Bool)] > (lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool,QTree_Bool) */
  assign lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet53_4Lcall_f_f0_d[0],
                                                                                            es_10_destruct_d[0],
                                                                                            es_11_1_destruct_d[0],
                                                                                            es_12_2_destruct_d[0]}), lizzieLet53_4Lcall_f_f0_d, es_10_destruct_d, es_11_1_destruct_d, es_12_2_destruct_d);
  assign {lizzieLet53_4Lcall_f_f0_r,
          es_10_destruct_r,
          es_11_1_destruct_r,
          es_12_2_destruct_r} = {4 {(lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_r && lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool,QTree_Bool) > (lizzieLet57_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d;
  logic lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_r;
  assign lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_r = ((! lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d[0]) || lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                 1'd0};
    else
      if (lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_r)
        lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d <= lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_d;
  QTree_Bool_t lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf;
  assign lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_r = (! lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet57_1_argbuf_d = (lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf[0] ? lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf :
                                   lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet57_1_argbuf_r && lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf[0]))
        lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                     1'd0};
      else if (((! lizzieLet57_1_argbuf_r) && (! lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf[0])))
        lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_buf <= lizzieLet53_4Lcall_f_f0_1es_10_1es_11_1_1es_12_2_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTf_f,
      Dcon Lcall_f_f0) : [(lizzieLet53_4Lcall_f_f1,Pointer_QTree_Bool),
                          (es_11_destruct,Pointer_QTree_Bool),
                          (es_12_1_destruct,Pointer_QTree_Bool),
                          (sc_0_13_destruct,Pointer_CTf_f)] > (lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0,CTf_f) */
  assign lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_d = Lcall_f_f0_dc((& {lizzieLet53_4Lcall_f_f1_d[0],
                                                                                            es_11_destruct_d[0],
                                                                                            es_12_1_destruct_d[0],
                                                                                            sc_0_13_destruct_d[0]}), lizzieLet53_4Lcall_f_f1_d, es_11_destruct_d, es_12_1_destruct_d, sc_0_13_destruct_d);
  assign {lizzieLet53_4Lcall_f_f1_r,
          es_11_destruct_r,
          es_12_1_destruct_r,
          sc_0_13_destruct_r} = {4 {(lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_r && lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_d[0])}};
  
  /* buf (Ty CTf_f) : (lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0,CTf_f) > (lizzieLet56_1_argbuf,CTf_f) */
  CTf_f_t lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d;
  logic lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_r;
  assign lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_r = ((! lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d[0]) || lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d <= {115'd0,
                                                                                 1'd0};
    else
      if (lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_r)
        lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d <= lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_d;
  CTf_f_t lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf;
  assign lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_r = (! lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf[0]);
  assign lizzieLet56_1_argbuf_d = (lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf[0] ? lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf :
                                   lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf <= {115'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet56_1_argbuf_r && lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf[0]))
        lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf <= {115'd0,
                                                                                     1'd0};
      else if (((! lizzieLet56_1_argbuf_r) && (! lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf[0])))
        lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_buf <= lizzieLet53_4Lcall_f_f1_1es_11_1es_12_1_1sc_0_13_1Lcall_f_f0_bufchan_d;
  
  /* dcon (Ty CTf_f,
      Dcon Lcall_f_f1) : [(lizzieLet53_4Lcall_f_f2,Pointer_QTree_Bool),
                          (es_12_destruct,Pointer_QTree_Bool),
                          (sc_0_12_destruct,Pointer_CTf_f),
                          (q1aen_2_destruct,Pointer_QTree_Int),
                          (t1aes_2_destruct,Pointer_QTree_Int)] > (lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1,CTf_f) */
  assign lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_d = Lcall_f_f1_dc((& {lizzieLet53_4Lcall_f_f2_d[0],
                                                                                                     es_12_destruct_d[0],
                                                                                                     sc_0_12_destruct_d[0],
                                                                                                     q1aen_2_destruct_d[0],
                                                                                                     t1aes_2_destruct_d[0]}), lizzieLet53_4Lcall_f_f2_d, es_12_destruct_d, sc_0_12_destruct_d, q1aen_2_destruct_d, t1aes_2_destruct_d);
  assign {lizzieLet53_4Lcall_f_f2_r,
          es_12_destruct_r,
          sc_0_12_destruct_r,
          q1aen_2_destruct_r,
          t1aes_2_destruct_r} = {5 {(lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_r && lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_d[0])}};
  
  /* buf (Ty CTf_f) : (lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1,CTf_f) > (lizzieLet55_1_argbuf,CTf_f) */
  CTf_f_t lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d;
  logic lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_r;
  assign lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_r = ((! lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d[0]) || lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d <= {115'd0,
                                                                                          1'd0};
    else
      if (lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_r)
        lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d <= lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_d;
  CTf_f_t lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf;
  assign lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_r = (! lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf[0]);
  assign lizzieLet55_1_argbuf_d = (lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf[0] ? lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf :
                                   lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf <= {115'd0,
                                                                                            1'd0};
    else
      if ((lizzieLet55_1_argbuf_r && lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf[0]))
        lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf <= {115'd0,
                                                                                              1'd0};
      else if (((! lizzieLet55_1_argbuf_r) && (! lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf[0])))
        lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_buf <= lizzieLet53_4Lcall_f_f2_1es_12_1sc_0_12_1q1aen_2_1t1aes_2_1Lcall_f_f1_bufchan_d;
  
  /* dcon (Ty CTf_f,
      Dcon Lcall_f_f2) : [(lizzieLet53_4Lcall_f_f3,Pointer_QTree_Bool),
                          (sc_0_11_destruct,Pointer_CTf_f),
                          (q1aen_1_destruct,Pointer_QTree_Int),
                          (t1aes_1_destruct,Pointer_QTree_Int),
                          (q2aeo_1_destruct,Pointer_QTree_Int),
                          (t2aet_1_destruct,Pointer_QTree_Int)] > (lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2,CTf_f) */
  assign lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_d = Lcall_f_f2_dc((& {lizzieLet53_4Lcall_f_f3_d[0],
                                                                                                                sc_0_11_destruct_d[0],
                                                                                                                q1aen_1_destruct_d[0],
                                                                                                                t1aes_1_destruct_d[0],
                                                                                                                q2aeo_1_destruct_d[0],
                                                                                                                t2aet_1_destruct_d[0]}), lizzieLet53_4Lcall_f_f3_d, sc_0_11_destruct_d, q1aen_1_destruct_d, t1aes_1_destruct_d, q2aeo_1_destruct_d, t2aet_1_destruct_d);
  assign {lizzieLet53_4Lcall_f_f3_r,
          sc_0_11_destruct_r,
          q1aen_1_destruct_r,
          t1aes_1_destruct_r,
          q2aeo_1_destruct_r,
          t2aet_1_destruct_r} = {6 {(lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_r && lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_d[0])}};
  
  /* buf (Ty CTf_f) : (lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2,CTf_f) > (lizzieLet54_1_argbuf,CTf_f) */
  CTf_f_t lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d;
  logic lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_r;
  assign lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_r = ((! lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d[0]) || lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d <= {115'd0,
                                                                                                     1'd0};
    else
      if (lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_r)
        lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d <= lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_d;
  CTf_f_t lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf;
  assign lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_r = (! lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf[0]);
  assign lizzieLet54_1_argbuf_d = (lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf[0] ? lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf :
                                   lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf <= {115'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet54_1_argbuf_r && lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf[0]))
        lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf <= {115'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet54_1_argbuf_r) && (! lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf[0])))
        lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_buf <= lizzieLet53_4Lcall_f_f3_1sc_0_11_1q1aen_1_1t1aes_1_1q2aeo_1_1t2aet_1_1Lcall_f_f2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet53_4Lf_fsbos,Pointer_QTree_Bool) > [(lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                             (lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet53_4Lf_fsbos_emitted;
  logic [1:0] lizzieLet53_4Lf_fsbos_done;
  assign lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_d = {lizzieLet53_4Lf_fsbos_d[16:1],
                                                               (lizzieLet53_4Lf_fsbos_d[0] && (! lizzieLet53_4Lf_fsbos_emitted[0]))};
  assign lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_d = {lizzieLet53_4Lf_fsbos_d[16:1],
                                                               (lizzieLet53_4Lf_fsbos_d[0] && (! lizzieLet53_4Lf_fsbos_emitted[1]))};
  assign lizzieLet53_4Lf_fsbos_done = (lizzieLet53_4Lf_fsbos_emitted | ({lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_d[0],
                                                                         lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_d[0]} & {lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_r,
                                                                                                                                   lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_r}));
  assign lizzieLet53_4Lf_fsbos_r = (& lizzieLet53_4Lf_fsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet53_4Lf_fsbos_emitted <= 2'd0;
    else
      lizzieLet53_4Lf_fsbos_emitted <= (lizzieLet53_4Lf_fsbos_r ? 2'd0 :
                                        lizzieLet53_4Lf_fsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1,Pointer_QTree_Bool) > (call_f_f_goConst,Go) */
  assign call_f_f_goConst_d = lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_d[0];
  assign lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_1_r = call_f_f_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2,Pointer_QTree_Bool) > (f_f_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d;
  logic lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_r;
  assign lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_r = ((! lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d[0]) || lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                     1'd0};
    else
      if (lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_r)
        lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d <= lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_r = (! lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]);
  assign f_f_resbuf_d = (lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf :
                         lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                       1'd0};
    else
      if ((f_f_resbuf_r && lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                         1'd0};
      else if (((! f_f_resbuf_r) && (! lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_buf <= lizzieLet53_4Lf_fsbos_1_merge_merge_merge_fork_2_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet5_1wild2XE_1_Eq,Bool) > (lizzieLet6_1_argbuf,Bool) */
  Bool_t lizzieLet5_1wild2XE_1_Eq_bufchan_d;
  logic lizzieLet5_1wild2XE_1_Eq_bufchan_r;
  assign lizzieLet5_1wild2XE_1_Eq_r = ((! lizzieLet5_1wild2XE_1_Eq_bufchan_d[0]) || lizzieLet5_1wild2XE_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_1wild2XE_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet5_1wild2XE_1_Eq_r)
        lizzieLet5_1wild2XE_1_Eq_bufchan_d <= lizzieLet5_1wild2XE_1_Eq_d;
  Bool_t lizzieLet5_1wild2XE_1_Eq_bufchan_buf;
  assign lizzieLet5_1wild2XE_1_Eq_bufchan_r = (! lizzieLet5_1wild2XE_1_Eq_bufchan_buf[0]);
  assign lizzieLet6_1_argbuf_d = (lizzieLet5_1wild2XE_1_Eq_bufchan_buf[0] ? lizzieLet5_1wild2XE_1_Eq_bufchan_buf :
                                  lizzieLet5_1wild2XE_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_1wild2XE_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet6_1_argbuf_r && lizzieLet5_1wild2XE_1_Eq_bufchan_buf[0]))
        lizzieLet5_1wild2XE_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet6_1_argbuf_r) && (! lizzieLet5_1wild2XE_1_Eq_bufchan_buf[0])))
        lizzieLet5_1wild2XE_1_Eq_bufchan_buf <= lizzieLet5_1wild2XE_1_Eq_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet7_1,MyBool) (va8v_3I#_3,Go) > [(lizzieLet7_1MyFalse,Go),
                                                         (lizzieLet7_1MyTrue,Go)] */
  logic [1:0] \va8v_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet7_1_d[0] && \va8v_3I#_3_d [0]))
      unique case (lizzieLet7_1_d[1:1])
        1'd0: \va8v_3I#_3_onehotd  = 2'd1;
        1'd1: \va8v_3I#_3_onehotd  = 2'd2;
        default: \va8v_3I#_3_onehotd  = 2'd0;
      endcase
    else \va8v_3I#_3_onehotd  = 2'd0;
  assign lizzieLet7_1MyFalse_d = \va8v_3I#_3_onehotd [0];
  assign lizzieLet7_1MyTrue_d = \va8v_3I#_3_onehotd [1];
  assign \va8v_3I#_3_r  = (| (\va8v_3I#_3_onehotd  & {lizzieLet7_1MyTrue_r,
                                                      lizzieLet7_1MyFalse_r}));
  assign lizzieLet7_1_r = \va8v_3I#_3_r ;
  
  /* fork (Ty Go) : (lizzieLet7_1MyFalse,Go) > [(lizzieLet7_1MyFalse_1,Go),
                                           (lizzieLet7_1MyFalse_2,Go)] */
  logic [1:0] lizzieLet7_1MyFalse_emitted;
  logic [1:0] lizzieLet7_1MyFalse_done;
  assign lizzieLet7_1MyFalse_1_d = (lizzieLet7_1MyFalse_d[0] && (! lizzieLet7_1MyFalse_emitted[0]));
  assign lizzieLet7_1MyFalse_2_d = (lizzieLet7_1MyFalse_d[0] && (! lizzieLet7_1MyFalse_emitted[1]));
  assign lizzieLet7_1MyFalse_done = (lizzieLet7_1MyFalse_emitted | ({lizzieLet7_1MyFalse_2_d[0],
                                                                     lizzieLet7_1MyFalse_1_d[0]} & {lizzieLet7_1MyFalse_2_r,
                                                                                                    lizzieLet7_1MyFalse_1_r}));
  assign lizzieLet7_1MyFalse_r = (& lizzieLet7_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyFalse_emitted <= 2'd0;
    else
      lizzieLet7_1MyFalse_emitted <= (lizzieLet7_1MyFalse_r ? 2'd0 :
                                      lizzieLet7_1MyFalse_done);
  
  /* buf (Ty Go) : (lizzieLet7_1MyFalse_1,Go) > (lizzieLet7_1MyFalse_1_argbuf,Go) */
  Go_t lizzieLet7_1MyFalse_1_bufchan_d;
  logic lizzieLet7_1MyFalse_1_bufchan_r;
  assign lizzieLet7_1MyFalse_1_r = ((! lizzieLet7_1MyFalse_1_bufchan_d[0]) || lizzieLet7_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet7_1MyFalse_1_r)
        lizzieLet7_1MyFalse_1_bufchan_d <= lizzieLet7_1MyFalse_1_d;
  Go_t lizzieLet7_1MyFalse_1_bufchan_buf;
  assign lizzieLet7_1MyFalse_1_bufchan_r = (! lizzieLet7_1MyFalse_1_bufchan_buf[0]);
  assign lizzieLet7_1MyFalse_1_argbuf_d = (lizzieLet7_1MyFalse_1_bufchan_buf[0] ? lizzieLet7_1MyFalse_1_bufchan_buf :
                                           lizzieLet7_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet7_1MyFalse_1_argbuf_r && lizzieLet7_1MyFalse_1_bufchan_buf[0]))
        lizzieLet7_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet7_1MyFalse_1_argbuf_r) && (! lizzieLet7_1MyFalse_1_bufchan_buf[0])))
        lizzieLet7_1MyFalse_1_bufchan_buf <= lizzieLet7_1MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(lizzieLet7_1MyFalse_1_argbuf,Go)] > (f''''''''1TupGo2,TupGo) */
  assign \f''''''''1TupGo2_d  = TupGo_dc((& {lizzieLet7_1MyFalse_1_argbuf_d[0]}), lizzieLet7_1MyFalse_1_argbuf_d);
  assign {lizzieLet7_1MyFalse_1_argbuf_r} = {1 {(\f''''''''1TupGo2_r  && \f''''''''1TupGo2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet7_1MyFalse_2,Go) > (lizzieLet7_1MyFalse_2_argbuf,Go) */
  Go_t lizzieLet7_1MyFalse_2_bufchan_d;
  logic lizzieLet7_1MyFalse_2_bufchan_r;
  assign lizzieLet7_1MyFalse_2_r = ((! lizzieLet7_1MyFalse_2_bufchan_d[0]) || lizzieLet7_1MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyFalse_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet7_1MyFalse_2_r)
        lizzieLet7_1MyFalse_2_bufchan_d <= lizzieLet7_1MyFalse_2_d;
  Go_t lizzieLet7_1MyFalse_2_bufchan_buf;
  assign lizzieLet7_1MyFalse_2_bufchan_r = (! lizzieLet7_1MyFalse_2_bufchan_buf[0]);
  assign lizzieLet7_1MyFalse_2_argbuf_d = (lizzieLet7_1MyFalse_2_bufchan_buf[0] ? lizzieLet7_1MyFalse_2_bufchan_buf :
                                           lizzieLet7_1MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet7_1MyFalse_2_argbuf_r && lizzieLet7_1MyFalse_2_bufchan_buf[0]))
        lizzieLet7_1MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet7_1MyFalse_2_argbuf_r) && (! lizzieLet7_1MyFalse_2_bufchan_buf[0])))
        lizzieLet7_1MyFalse_2_bufchan_buf <= lizzieLet7_1MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet7_1MyTrue,Go) > [(lizzieLet7_1MyTrue_1,Go),
                                          (lizzieLet7_1MyTrue_2,Go)] */
  logic [1:0] lizzieLet7_1MyTrue_emitted;
  logic [1:0] lizzieLet7_1MyTrue_done;
  assign lizzieLet7_1MyTrue_1_d = (lizzieLet7_1MyTrue_d[0] && (! lizzieLet7_1MyTrue_emitted[0]));
  assign lizzieLet7_1MyTrue_2_d = (lizzieLet7_1MyTrue_d[0] && (! lizzieLet7_1MyTrue_emitted[1]));
  assign lizzieLet7_1MyTrue_done = (lizzieLet7_1MyTrue_emitted | ({lizzieLet7_1MyTrue_2_d[0],
                                                                   lizzieLet7_1MyTrue_1_d[0]} & {lizzieLet7_1MyTrue_2_r,
                                                                                                 lizzieLet7_1MyTrue_1_r}));
  assign lizzieLet7_1MyTrue_r = (& lizzieLet7_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyTrue_emitted <= 2'd0;
    else
      lizzieLet7_1MyTrue_emitted <= (lizzieLet7_1MyTrue_r ? 2'd0 :
                                     lizzieLet7_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet7_1MyTrue_1,Go)] > (lizzieLet7_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign lizzieLet7_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet7_1MyTrue_1_d[0]}), lizzieLet7_1MyTrue_1_d);
  assign {lizzieLet7_1MyTrue_1_r} = {1 {(lizzieLet7_1MyTrue_1QNone_Bool_r && lizzieLet7_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet7_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet9_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d;
  logic lizzieLet7_1MyTrue_1QNone_Bool_bufchan_r;
  assign lizzieLet7_1MyTrue_1QNone_Bool_r = ((! lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d[0]) || lizzieLet7_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet7_1MyTrue_1QNone_Bool_r)
        lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d <= lizzieLet7_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf;
  assign lizzieLet7_1MyTrue_1QNone_Bool_bufchan_r = (! lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf[0] ? lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf :
                                  lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        lizzieLet7_1MyTrue_1QNone_Bool_bufchan_buf <= lizzieLet7_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet7_1MyTrue_2,Go) > (lizzieLet7_1MyTrue_2_argbuf,Go) */
  Go_t lizzieLet7_1MyTrue_2_bufchan_d;
  logic lizzieLet7_1MyTrue_2_bufchan_r;
  assign lizzieLet7_1MyTrue_2_r = ((! lizzieLet7_1MyTrue_2_bufchan_d[0]) || lizzieLet7_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet7_1MyTrue_2_r)
        lizzieLet7_1MyTrue_2_bufchan_d <= lizzieLet7_1MyTrue_2_d;
  Go_t lizzieLet7_1MyTrue_2_bufchan_buf;
  assign lizzieLet7_1MyTrue_2_bufchan_r = (! lizzieLet7_1MyTrue_2_bufchan_buf[0]);
  assign lizzieLet7_1MyTrue_2_argbuf_d = (lizzieLet7_1MyTrue_2_bufchan_buf[0] ? lizzieLet7_1MyTrue_2_bufchan_buf :
                                          lizzieLet7_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet7_1MyTrue_2_argbuf_r && lizzieLet7_1MyTrue_2_bufchan_buf[0]))
        lizzieLet7_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet7_1MyTrue_2_argbuf_r) && (! lizzieLet7_1MyTrue_2_bufchan_buf[0])))
        lizzieLet7_1MyTrue_2_bufchan_buf <= lizzieLet7_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet7_2,MyBool) (va8v_4I#,Pointer_CTf''''''''_f'''''''') > [(lizzieLet7_2MyFalse,Pointer_CTf''''''''_f''''''''),
                                                                                                             (lizzieLet7_2MyTrue,Pointer_CTf''''''''_f'''''''')] */
  logic [1:0] \va8v_4I#_onehotd ;
  always_comb
    if ((lizzieLet7_2_d[0] && \va8v_4I#_d [0]))
      unique case (lizzieLet7_2_d[1:1])
        1'd0: \va8v_4I#_onehotd  = 2'd1;
        1'd1: \va8v_4I#_onehotd  = 2'd2;
        default: \va8v_4I#_onehotd  = 2'd0;
      endcase
    else \va8v_4I#_onehotd  = 2'd0;
  assign lizzieLet7_2MyFalse_d = {\va8v_4I#_d [16:1],
                                  \va8v_4I#_onehotd [0]};
  assign lizzieLet7_2MyTrue_d = {\va8v_4I#_d [16:1],
                                 \va8v_4I#_onehotd [1]};
  assign \va8v_4I#_r  = (| (\va8v_4I#_onehotd  & {lizzieLet7_2MyTrue_r,
                                                  lizzieLet7_2MyFalse_r}));
  assign lizzieLet7_2_r = \va8v_4I#_r ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet7_2MyFalse,Pointer_CTf''''''''_f'''''''') > (lizzieLet7_2MyFalse_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyFalse_bufchan_d;
  logic lizzieLet7_2MyFalse_bufchan_r;
  assign lizzieLet7_2MyFalse_r = ((! lizzieLet7_2MyFalse_bufchan_d[0]) || lizzieLet7_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet7_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet7_2MyFalse_r)
        lizzieLet7_2MyFalse_bufchan_d <= lizzieLet7_2MyFalse_d;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyFalse_bufchan_buf;
  assign lizzieLet7_2MyFalse_bufchan_r = (! lizzieLet7_2MyFalse_bufchan_buf[0]);
  assign lizzieLet7_2MyFalse_1_argbuf_d = (lizzieLet7_2MyFalse_bufchan_buf[0] ? lizzieLet7_2MyFalse_bufchan_buf :
                                           lizzieLet7_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet7_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet7_2MyFalse_1_argbuf_r && lizzieLet7_2MyFalse_bufchan_buf[0]))
        lizzieLet7_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet7_2MyFalse_1_argbuf_r) && (! lizzieLet7_2MyFalse_bufchan_buf[0])))
        lizzieLet7_2MyFalse_bufchan_buf <= lizzieLet7_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (lizzieLet7_2MyTrue,Pointer_CTf''''''''_f'''''''') > (lizzieLet7_2MyTrue_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyTrue_bufchan_d;
  logic lizzieLet7_2MyTrue_bufchan_r;
  assign lizzieLet7_2MyTrue_r = ((! lizzieLet7_2MyTrue_bufchan_d[0]) || lizzieLet7_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet7_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet7_2MyTrue_r)
        lizzieLet7_2MyTrue_bufchan_d <= lizzieLet7_2MyTrue_d;
  \Pointer_CTf''''''''_f''''''''_t  lizzieLet7_2MyTrue_bufchan_buf;
  assign lizzieLet7_2MyTrue_bufchan_r = (! lizzieLet7_2MyTrue_bufchan_buf[0]);
  assign lizzieLet7_2MyTrue_1_argbuf_d = (lizzieLet7_2MyTrue_bufchan_buf[0] ? lizzieLet7_2MyTrue_bufchan_buf :
                                          lizzieLet7_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet7_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet7_2MyTrue_1_argbuf_r && lizzieLet7_2MyTrue_bufchan_buf[0]))
        lizzieLet7_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet7_2MyTrue_1_argbuf_r) && (! lizzieLet7_2MyTrue_bufchan_buf[0])))
        lizzieLet7_2MyTrue_bufchan_buf <= lizzieLet7_2MyTrue_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1ae6_goMux_mux,Pointer_QTree_Int) > (m1ae6_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1ae6_goMux_mux_bufchan_d;
  logic m1ae6_goMux_mux_bufchan_r;
  assign m1ae6_goMux_mux_r = ((! m1ae6_goMux_mux_bufchan_d[0]) || m1ae6_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae6_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1ae6_goMux_mux_r)
        m1ae6_goMux_mux_bufchan_d <= m1ae6_goMux_mux_d;
  Pointer_QTree_Int_t m1ae6_goMux_mux_bufchan_buf;
  assign m1ae6_goMux_mux_bufchan_r = (! m1ae6_goMux_mux_bufchan_buf[0]);
  assign m1ae6_1_argbuf_d = (m1ae6_goMux_mux_bufchan_buf[0] ? m1ae6_goMux_mux_bufchan_buf :
                             m1ae6_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae6_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1ae6_1_argbuf_r && m1ae6_goMux_mux_bufchan_buf[0]))
        m1ae6_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1ae6_1_argbuf_r) && (! m1ae6_goMux_mux_bufchan_buf[0])))
        m1ae6_goMux_mux_bufchan_buf <= m1ae6_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2ae7_goMux_mux,Pointer_QTree_Int) > (m2ae7_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ae7_goMux_mux_bufchan_d;
  logic m2ae7_goMux_mux_bufchan_r;
  assign m2ae7_goMux_mux_r = ((! m2ae7_goMux_mux_bufchan_d[0]) || m2ae7_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae7_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2ae7_goMux_mux_r)
        m2ae7_goMux_mux_bufchan_d <= m2ae7_goMux_mux_d;
  Pointer_QTree_Int_t m2ae7_goMux_mux_bufchan_buf;
  assign m2ae7_goMux_mux_bufchan_r = (! m2ae7_goMux_mux_bufchan_buf[0]);
  assign m2ae7_1_argbuf_d = (m2ae7_goMux_mux_bufchan_buf[0] ? m2ae7_goMux_mux_bufchan_buf :
                             m2ae7_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae7_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ae7_1_argbuf_r && m2ae7_goMux_mux_bufchan_buf[0]))
        m2ae7_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ae7_1_argbuf_r) && (! m2ae7_goMux_mux_bufchan_buf[0])))
        m2ae7_goMux_mux_bufchan_buf <= m2ae7_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a84_destruct,Pointer_QTree_Bool) > (q1a84_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a84_destruct_bufchan_d;
  logic q1a84_destruct_bufchan_r;
  assign q1a84_destruct_r = ((! q1a84_destruct_bufchan_d[0]) || q1a84_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a84_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a84_destruct_r) q1a84_destruct_bufchan_d <= q1a84_destruct_d;
  Pointer_QTree_Bool_t q1a84_destruct_bufchan_buf;
  assign q1a84_destruct_bufchan_r = (! q1a84_destruct_bufchan_buf[0]);
  assign q1a84_1_argbuf_d = (q1a84_destruct_bufchan_buf[0] ? q1a84_destruct_bufchan_buf :
                             q1a84_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a84_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a84_1_argbuf_r && q1a84_destruct_bufchan_buf[0]))
        q1a84_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a84_1_argbuf_r) && (! q1a84_destruct_bufchan_buf[0])))
        q1a84_destruct_bufchan_buf <= q1a84_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1aen_3_destruct,Pointer_QTree_Int) > (q1aen_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1aen_3_destruct_bufchan_d;
  logic q1aen_3_destruct_bufchan_r;
  assign q1aen_3_destruct_r = ((! q1aen_3_destruct_bufchan_d[0]) || q1aen_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aen_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1aen_3_destruct_r)
        q1aen_3_destruct_bufchan_d <= q1aen_3_destruct_d;
  Pointer_QTree_Int_t q1aen_3_destruct_bufchan_buf;
  assign q1aen_3_destruct_bufchan_r = (! q1aen_3_destruct_bufchan_buf[0]);
  assign q1aen_3_1_argbuf_d = (q1aen_3_destruct_bufchan_buf[0] ? q1aen_3_destruct_bufchan_buf :
                               q1aen_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aen_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1aen_3_1_argbuf_r && q1aen_3_destruct_bufchan_buf[0]))
        q1aen_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1aen_3_1_argbuf_r) && (! q1aen_3_destruct_bufchan_buf[0])))
        q1aen_3_destruct_bufchan_buf <= q1aen_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a85_1_destruct,Pointer_QTree_Bool) > (q2a85_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a85_1_destruct_bufchan_d;
  logic q2a85_1_destruct_bufchan_r;
  assign q2a85_1_destruct_r = ((! q2a85_1_destruct_bufchan_d[0]) || q2a85_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a85_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a85_1_destruct_r)
        q2a85_1_destruct_bufchan_d <= q2a85_1_destruct_d;
  Pointer_QTree_Bool_t q2a85_1_destruct_bufchan_buf;
  assign q2a85_1_destruct_bufchan_r = (! q2a85_1_destruct_bufchan_buf[0]);
  assign q2a85_1_1_argbuf_d = (q2a85_1_destruct_bufchan_buf[0] ? q2a85_1_destruct_bufchan_buf :
                               q2a85_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a85_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a85_1_1_argbuf_r && q2a85_1_destruct_bufchan_buf[0]))
        q2a85_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a85_1_1_argbuf_r) && (! q2a85_1_destruct_bufchan_buf[0])))
        q2a85_1_destruct_bufchan_buf <= q2a85_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2aeo_2_destruct,Pointer_QTree_Int) > (q2aeo_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2aeo_2_destruct_bufchan_d;
  logic q2aeo_2_destruct_bufchan_r;
  assign q2aeo_2_destruct_r = ((! q2aeo_2_destruct_bufchan_d[0]) || q2aeo_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aeo_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2aeo_2_destruct_r)
        q2aeo_2_destruct_bufchan_d <= q2aeo_2_destruct_d;
  Pointer_QTree_Int_t q2aeo_2_destruct_bufchan_buf;
  assign q2aeo_2_destruct_bufchan_r = (! q2aeo_2_destruct_bufchan_buf[0]);
  assign q2aeo_2_1_argbuf_d = (q2aeo_2_destruct_bufchan_buf[0] ? q2aeo_2_destruct_bufchan_buf :
                               q2aeo_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aeo_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2aeo_2_1_argbuf_r && q2aeo_2_destruct_bufchan_buf[0]))
        q2aeo_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2aeo_2_1_argbuf_r) && (! q2aeo_2_destruct_bufchan_buf[0])))
        q2aeo_2_destruct_bufchan_buf <= q2aeo_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a86_2_destruct,Pointer_QTree_Bool) > (q3a86_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a86_2_destruct_bufchan_d;
  logic q3a86_2_destruct_bufchan_r;
  assign q3a86_2_destruct_r = ((! q3a86_2_destruct_bufchan_d[0]) || q3a86_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a86_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a86_2_destruct_r)
        q3a86_2_destruct_bufchan_d <= q3a86_2_destruct_d;
  Pointer_QTree_Bool_t q3a86_2_destruct_bufchan_buf;
  assign q3a86_2_destruct_bufchan_r = (! q3a86_2_destruct_bufchan_buf[0]);
  assign q3a86_2_1_argbuf_d = (q3a86_2_destruct_bufchan_buf[0] ? q3a86_2_destruct_bufchan_buf :
                               q3a86_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a86_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a86_2_1_argbuf_r && q3a86_2_destruct_bufchan_buf[0]))
        q3a86_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a86_2_1_argbuf_r) && (! q3a86_2_destruct_bufchan_buf[0])))
        q3a86_2_destruct_bufchan_buf <= q3a86_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3aep_1_destruct,Pointer_QTree_Int) > (q3aep_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3aep_1_destruct_bufchan_d;
  logic q3aep_1_destruct_bufchan_r;
  assign q3aep_1_destruct_r = ((! q3aep_1_destruct_bufchan_d[0]) || q3aep_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aep_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aep_1_destruct_r)
        q3aep_1_destruct_bufchan_d <= q3aep_1_destruct_d;
  Pointer_QTree_Int_t q3aep_1_destruct_bufchan_buf;
  assign q3aep_1_destruct_bufchan_r = (! q3aep_1_destruct_bufchan_buf[0]);
  assign q3aep_1_1_argbuf_d = (q3aep_1_destruct_bufchan_buf[0] ? q3aep_1_destruct_bufchan_buf :
                               q3aep_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aep_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aep_1_1_argbuf_r && q3aep_1_destruct_bufchan_buf[0]))
        q3aep_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aep_1_1_argbuf_r) && (! q3aep_1_destruct_bufchan_buf[0])))
        q3aep_1_destruct_bufchan_buf <= q3aep_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4a87_3_destruct,Pointer_QTree_Bool) > (q4a87_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4a87_3_destruct_bufchan_d;
  logic q4a87_3_destruct_bufchan_r;
  assign q4a87_3_destruct_r = ((! q4a87_3_destruct_bufchan_d[0]) || q4a87_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a87_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a87_3_destruct_r)
        q4a87_3_destruct_bufchan_d <= q4a87_3_destruct_d;
  Pointer_QTree_Bool_t q4a87_3_destruct_bufchan_buf;
  assign q4a87_3_destruct_bufchan_r = (! q4a87_3_destruct_bufchan_buf[0]);
  assign q4a87_3_1_argbuf_d = (q4a87_3_destruct_bufchan_buf[0] ? q4a87_3_destruct_bufchan_buf :
                               q4a87_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a87_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a87_3_1_argbuf_r && q4a87_3_destruct_bufchan_buf[0]))
        q4a87_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a87_3_1_argbuf_r) && (! q4a87_3_destruct_bufchan_buf[0])))
        q4a87_3_destruct_bufchan_buf <= q4a87_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a8u_goMux_mux,Pointer_QTree_Int) > (q4a8u_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a8u_goMux_mux_bufchan_d;
  logic q4a8u_goMux_mux_bufchan_r;
  assign q4a8u_goMux_mux_r = ((! q4a8u_goMux_mux_bufchan_d[0]) || q4a8u_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8u_goMux_mux_r)
        q4a8u_goMux_mux_bufchan_d <= q4a8u_goMux_mux_d;
  Pointer_QTree_Int_t q4a8u_goMux_mux_bufchan_buf;
  assign q4a8u_goMux_mux_bufchan_r = (! q4a8u_goMux_mux_bufchan_buf[0]);
  assign q4a8u_1_argbuf_d = (q4a8u_goMux_mux_bufchan_buf[0] ? q4a8u_goMux_mux_bufchan_buf :
                             q4a8u_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8u_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8u_1_argbuf_r && q4a8u_goMux_mux_bufchan_buf[0]))
        q4a8u_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8u_1_argbuf_r) && (! q4a8u_goMux_mux_bufchan_buf[0])))
        q4a8u_goMux_mux_bufchan_buf <= q4a8u_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf,CT$wnnz) > (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) */
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= {115'd0, 1'd0};
    else
      if (readPointer_CT$wnnzscfarg_0_1_argbuf_r)
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnzscfarg_0_1_argbuf_d;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf :
                                                       readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
      else if (((! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnzscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb,CT$wnnz) > [(lizzieLet44_1,CT$wnnz),
                                                                          (lizzieLet44_2,CT$wnnz),
                                                                          (lizzieLet44_3,CT$wnnz),
                                                                          (lizzieLet44_4,CT$wnnz)] */
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet44_1_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet44_2_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet44_3_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet44_4_d = {readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet44_4_d[0],
                                                                                                               lizzieLet44_3_d[0],
                                                                                                               lizzieLet44_2_d[0],
                                                                                                               lizzieLet44_1_d[0]} & {lizzieLet44_4_r,
                                                                                                                                      lizzieLet44_3_r,
                                                                                                                                      lizzieLet44_2_r,
                                                                                                                                      lizzieLet44_1_r}));
  assign readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_CT$wnnzscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTf''''''''_f'''''''') : (readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf,CTf''''''''_f'''''''') > (readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb,CTf''''''''_f'''''''') */
  \CTf''''''''_f''''''''_t  \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d  <= {67'd0,
                                                                           1'd0};
    else
      if (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_r )
        \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_d ;
  \CTf''''''''_f''''''''_t  \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf  :
                                                                         \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                             1'd0};
    else
      if ((\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                               1'd0};
      else if (((! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf''''''''_f'''''''') : (readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb,CTf''''''''_f'''''''') > [(lizzieLet48_1,CTf''''''''_f''''''''),
                                                                                                                      (lizzieLet48_2,CTf''''''''_f''''''''),
                                                                                                                      (lizzieLet48_3,CTf''''''''_f''''''''),
                                                                                                                      (lizzieLet48_4,CTf''''''''_f'''''''')] */
  logic [3:0] \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet48_1_d = {\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet48_2_d = {\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet48_3_d = {\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet48_4_d = {\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet48_4_d[0],
                                                                                                                                                   lizzieLet48_3_d[0],
                                                                                                                                                   lizzieLet48_2_d[0],
                                                                                                                                                   lizzieLet48_1_d[0]} & {lizzieLet48_4_r,
                                                                                                                                                                          lizzieLet48_3_r,
                                                                                                                                                                          lizzieLet48_2_r,
                                                                                                                                                                          lizzieLet48_1_r}));
  assign \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                             \readPointer_CTf''''''''_f''''''''scfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf_f) : (readPointer_CTf_fscfarg_0_2_1_argbuf,CTf_f) > (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb,CTf_f) */
  CTf_f_t readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_r = ((! readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d <= {115'd0, 1'd0};
    else
      if (readPointer_CTf_fscfarg_0_2_1_argbuf_r)
        readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTf_fscfarg_0_2_1_argbuf_d;
  CTf_f_t readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf :
                                                       readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_r && readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf <= {115'd0, 1'd0};
      else if (((! readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTf_fscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf_f) : (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb,CTf_f) > [(lizzieLet53_1,CTf_f),
                                                                      (lizzieLet53_2,CTf_f),
                                                                      (lizzieLet53_3,CTf_f),
                                                                      (lizzieLet53_4,CTf_f)] */
  logic [3:0] readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet53_1_d = {readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet53_2_d = {readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet53_3_d = {readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet53_4_d = {readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[115:1],
                            (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet53_4_d[0],
                                                                                                               lizzieLet53_3_d[0],
                                                                                                               lizzieLet53_2_d[0],
                                                                                                               lizzieLet53_1_d[0]} & {lizzieLet53_4_r,
                                                                                                                                      lizzieLet53_3_r,
                                                                                                                                      lizzieLet53_2_r,
                                                                                                                                      lizzieLet53_1_r}));
  assign readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_CTf_fscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_BoolwspF_1_1_argbuf,QTree_Bool) > (readPointer_QTree_BoolwspF_1_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_BoolwspF_1_1_argbuf_r = ((! readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_BoolwspF_1_1_argbuf_r)
        readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d <= readPointer_QTree_BoolwspF_1_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_r = (! readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d = (readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_BoolwspF_1_1_argbuf_rwb_r && readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_BoolwspF_1_1_argbuf_rwb_r) && (! readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_buf <= readPointer_QTree_BoolwspF_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_BoolwspF_1_1_argbuf_rwb,QTree_Bool) > [(lizzieLet1_1,QTree_Bool),
                                                                                 (lizzieLet1_2,QTree_Bool),
                                                                                 (lizzieLet1_3,QTree_Bool),
                                                                                 (lizzieLet1_4,QTree_Bool)] */
  logic [3:0] readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_BoolwspF_1_1_argbuf_rwb_done;
  assign lizzieLet1_1_d = {readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet1_2_d = {readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet1_3_d = {readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet1_4_d = {readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_BoolwspF_1_1_argbuf_rwb_done = (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted | ({lizzieLet1_4_d[0],
                                                                                                                 lizzieLet1_3_d[0],
                                                                                                                 lizzieLet1_2_d[0],
                                                                                                                 lizzieLet1_1_d[0]} & {lizzieLet1_4_r,
                                                                                                                                       lizzieLet1_3_r,
                                                                                                                                       lizzieLet1_2_r,
                                                                                                                                       lizzieLet1_1_r}));
  assign readPointer_QTree_BoolwspF_1_1_argbuf_rwb_r = (& readPointer_QTree_BoolwspF_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_BoolwspF_1_1_argbuf_rwb_emitted <= (readPointer_QTree_BoolwspF_1_1_argbuf_rwb_r ? 4'd0 :
                                                            readPointer_QTree_BoolwspF_1_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1ae6_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1ae6_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1ae6_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1ae6_1_argbuf_r = ((! readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1ae6_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1ae6_1_argbuf_r)
        readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d <= readPointer_QTree_Intm1ae6_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1ae6_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1ae6_1_argbuf_rwb_d = (readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1ae6_1_argbuf_rwb_r && readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1ae6_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1ae6_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1ae6_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1ae6_1_argbuf_rwb,QTree_Int) > [(lizzieLet12_1,QTree_Int),
                                                                             (lizzieLet12_2,QTree_Int),
                                                                             (lizzieLet12_3,QTree_Int),
                                                                             (lizzieLet12_4,QTree_Int),
                                                                             (lizzieLet12_5,QTree_Int)] */
  logic [4:0] readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted;
  logic [4:0] readPointer_QTree_Intm1ae6_1_argbuf_rwb_done;
  assign lizzieLet12_1_d = {readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet12_2_d = {readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet12_3_d = {readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet12_4_d = {readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet12_5_d = {readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm1ae6_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted[4]))};
  assign readPointer_QTree_Intm1ae6_1_argbuf_rwb_done = (readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted | ({lizzieLet12_5_d[0],
                                                                                                             lizzieLet12_4_d[0],
                                                                                                             lizzieLet12_3_d[0],
                                                                                                             lizzieLet12_2_d[0],
                                                                                                             lizzieLet12_1_d[0]} & {lizzieLet12_5_r,
                                                                                                                                    lizzieLet12_4_r,
                                                                                                                                    lizzieLet12_3_r,
                                                                                                                                    lizzieLet12_2_r,
                                                                                                                                    lizzieLet12_1_r}));
  assign readPointer_QTree_Intm1ae6_1_argbuf_rwb_r = (& readPointer_QTree_Intm1ae6_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted <= 5'd0;
    else
      readPointer_QTree_Intm1ae6_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1ae6_1_argbuf_rwb_r ? 5'd0 :
                                                          readPointer_QTree_Intm1ae6_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2ae7_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2ae7_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2ae7_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2ae7_1_argbuf_r = ((! readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2ae7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2ae7_1_argbuf_r)
        readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d <= readPointer_QTree_Intm2ae7_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2ae7_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2ae7_1_argbuf_rwb_d = (readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2ae7_1_argbuf_rwb_r && readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2ae7_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2ae7_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2ae7_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intq4a8u_1_argbuf,QTree_Int) > (readPointer_QTree_Intq4a8u_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intq4a8u_1_argbuf_r = ((! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intq4a8u_1_argbuf_r)
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d <= readPointer_QTree_Intq4a8u_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intq4a8u_1_argbuf_bufchan_r = (! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_d = (readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intq4a8u_1_argbuf_rwb_r && readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intq4a8u_1_argbuf_rwb_r) && (! readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intq4a8u_1_argbuf_bufchan_buf <= readPointer_QTree_Intq4a8u_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intq4a8u_1_argbuf_rwb,QTree_Int) > [(lizzieLet3_1,QTree_Int),
                                                                             (lizzieLet3_2,QTree_Int),
                                                                             (lizzieLet3_3,QTree_Int),
                                                                             (lizzieLet3_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_Intq4a8u_1_argbuf_rwb_done;
  assign lizzieLet3_1_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet3_2_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet3_3_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet3_4_d = {readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intq4a8u_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_done = (readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted | ({lizzieLet3_4_d[0],
                                                                                                             lizzieLet3_3_d[0],
                                                                                                             lizzieLet3_2_d[0],
                                                                                                             lizzieLet3_1_d[0]} & {lizzieLet3_4_r,
                                                                                                                                   lizzieLet3_3_r,
                                                                                                                                   lizzieLet3_2_r,
                                                                                                                                   lizzieLet3_1_r}));
  assign readPointer_QTree_Intq4a8u_1_argbuf_rwb_r = (& readPointer_QTree_Intq4a8u_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_Intq4a8u_1_argbuf_rwb_emitted <= (readPointer_QTree_Intq4a8u_1_argbuf_rwb_r ? 4'd0 :
                                                          readPointer_QTree_Intq4a8u_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (sc_0_10_destruct,Pointer_CTf''''''''_f'''''''') > (sc_0_10_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTf''''''''_f''''''''_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (sc_0_14_destruct,Pointer_CTf_f) > (sc_0_14_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  Pointer_CTf_f_t sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (sc_0_6_destruct,Pointer_CT$wnnz) > (sc_0_6_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wnnz_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (scfarg_0_1_goMux_mux,Pointer_CTf''''''''_f'''''''') > (scfarg_0_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf''''''''_f''''''''_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (scfarg_0_2_goMux_mux,Pointer_CTf_f) > (scfarg_0_2_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTf_f_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (scfarg_0_goMux_mux,Pointer_CT$wnnz) > (scfarg_0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aes_3_destruct,Pointer_QTree_Int) > (t1aes_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aes_3_destruct_bufchan_d;
  logic t1aes_3_destruct_bufchan_r;
  assign t1aes_3_destruct_r = ((! t1aes_3_destruct_bufchan_d[0]) || t1aes_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aes_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aes_3_destruct_r)
        t1aes_3_destruct_bufchan_d <= t1aes_3_destruct_d;
  Pointer_QTree_Int_t t1aes_3_destruct_bufchan_buf;
  assign t1aes_3_destruct_bufchan_r = (! t1aes_3_destruct_bufchan_buf[0]);
  assign t1aes_3_1_argbuf_d = (t1aes_3_destruct_bufchan_buf[0] ? t1aes_3_destruct_bufchan_buf :
                               t1aes_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aes_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aes_3_1_argbuf_r && t1aes_3_destruct_bufchan_buf[0]))
        t1aes_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aes_3_1_argbuf_r) && (! t1aes_3_destruct_bufchan_buf[0])))
        t1aes_3_destruct_bufchan_buf <= t1aes_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aet_2_destruct,Pointer_QTree_Int) > (t2aet_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aet_2_destruct_bufchan_d;
  logic t2aet_2_destruct_bufchan_r;
  assign t2aet_2_destruct_r = ((! t2aet_2_destruct_bufchan_d[0]) || t2aet_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aet_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aet_2_destruct_r)
        t2aet_2_destruct_bufchan_d <= t2aet_2_destruct_d;
  Pointer_QTree_Int_t t2aet_2_destruct_bufchan_buf;
  assign t2aet_2_destruct_bufchan_r = (! t2aet_2_destruct_bufchan_buf[0]);
  assign t2aet_2_1_argbuf_d = (t2aet_2_destruct_bufchan_buf[0] ? t2aet_2_destruct_bufchan_buf :
                               t2aet_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aet_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aet_2_1_argbuf_r && t2aet_2_destruct_bufchan_buf[0]))
        t2aet_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aet_2_1_argbuf_r) && (! t2aet_2_destruct_bufchan_buf[0])))
        t2aet_2_destruct_bufchan_buf <= t2aet_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aeu_1_destruct,Pointer_QTree_Int) > (t3aeu_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aeu_1_destruct_bufchan_d;
  logic t3aeu_1_destruct_bufchan_r;
  assign t3aeu_1_destruct_r = ((! t3aeu_1_destruct_bufchan_d[0]) || t3aeu_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeu_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aeu_1_destruct_r)
        t3aeu_1_destruct_bufchan_d <= t3aeu_1_destruct_d;
  Pointer_QTree_Int_t t3aeu_1_destruct_bufchan_buf;
  assign t3aeu_1_destruct_bufchan_r = (! t3aeu_1_destruct_bufchan_buf[0]);
  assign t3aeu_1_1_argbuf_d = (t3aeu_1_destruct_bufchan_buf[0] ? t3aeu_1_destruct_bufchan_buf :
                               t3aeu_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeu_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aeu_1_1_argbuf_r && t3aeu_1_destruct_bufchan_buf[0]))
        t3aeu_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aeu_1_1_argbuf_r) && (! t3aeu_1_destruct_bufchan_buf[0])))
        t3aeu_1_destruct_bufchan_buf <= t3aeu_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aev_destruct,Pointer_QTree_Int) > (t4aev_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aev_destruct_bufchan_d;
  logic t4aev_destruct_bufchan_r;
  assign t4aev_destruct_r = ((! t4aev_destruct_bufchan_d[0]) || t4aev_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aev_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aev_destruct_r) t4aev_destruct_bufchan_d <= t4aev_destruct_d;
  Pointer_QTree_Int_t t4aev_destruct_bufchan_buf;
  assign t4aev_destruct_bufchan_r = (! t4aev_destruct_bufchan_buf[0]);
  assign t4aev_1_argbuf_d = (t4aev_destruct_bufchan_buf[0] ? t4aev_destruct_bufchan_buf :
                             t4aev_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aev_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aev_1_argbuf_r && t4aev_destruct_bufchan_buf[0]))
        t4aev_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aev_1_argbuf_r) && (! t4aev_destruct_bufchan_buf[0])))
        t4aev_destruct_bufchan_buf <= t4aev_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tlae2_3_destruct,Pointer_QTree_Int) > (tlae2_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tlae2_3_destruct_bufchan_d;
  logic tlae2_3_destruct_bufchan_r;
  assign tlae2_3_destruct_r = ((! tlae2_3_destruct_bufchan_d[0]) || tlae2_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tlae2_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tlae2_3_destruct_r)
        tlae2_3_destruct_bufchan_d <= tlae2_3_destruct_d;
  Pointer_QTree_Int_t tlae2_3_destruct_bufchan_buf;
  assign tlae2_3_destruct_bufchan_r = (! tlae2_3_destruct_bufchan_buf[0]);
  assign tlae2_3_1_argbuf_d = (tlae2_3_destruct_bufchan_buf[0] ? tlae2_3_destruct_bufchan_buf :
                               tlae2_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tlae2_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tlae2_3_1_argbuf_r && tlae2_3_destruct_bufchan_buf[0]))
        tlae2_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tlae2_3_1_argbuf_r) && (! tlae2_3_destruct_bufchan_buf[0])))
        tlae2_3_destruct_bufchan_buf <= tlae2_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (tlaea_destruct,Pointer_QTree_Int) > (tlaea_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t tlaea_destruct_bufchan_d;
  logic tlaea_destruct_bufchan_r;
  assign tlaea_destruct_r = ((! tlaea_destruct_bufchan_d[0]) || tlaea_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tlaea_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (tlaea_destruct_r) tlaea_destruct_bufchan_d <= tlaea_destruct_d;
  Pointer_QTree_Int_t tlaea_destruct_bufchan_buf;
  assign tlaea_destruct_bufchan_r = (! tlaea_destruct_bufchan_buf[0]);
  assign tlaea_1_argbuf_d = (tlaea_destruct_bufchan_buf[0] ? tlaea_destruct_bufchan_buf :
                             tlaea_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) tlaea_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((tlaea_1_argbuf_r && tlaea_destruct_bufchan_buf[0]))
        tlaea_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! tlaea_1_argbuf_r) && (! tlaea_destruct_bufchan_buf[0])))
        tlaea_destruct_bufchan_buf <= tlaea_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (trae3_2_destruct,Pointer_QTree_Int) > (trae3_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t trae3_2_destruct_bufchan_d;
  logic trae3_2_destruct_bufchan_r;
  assign trae3_2_destruct_r = ((! trae3_2_destruct_bufchan_d[0]) || trae3_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) trae3_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (trae3_2_destruct_r)
        trae3_2_destruct_bufchan_d <= trae3_2_destruct_d;
  Pointer_QTree_Int_t trae3_2_destruct_bufchan_buf;
  assign trae3_2_destruct_bufchan_r = (! trae3_2_destruct_bufchan_buf[0]);
  assign trae3_2_1_argbuf_d = (trae3_2_destruct_bufchan_buf[0] ? trae3_2_destruct_bufchan_buf :
                               trae3_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) trae3_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((trae3_2_1_argbuf_r && trae3_2_destruct_bufchan_buf[0]))
        trae3_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! trae3_2_1_argbuf_r) && (! trae3_2_destruct_bufchan_buf[0])))
        trae3_2_destruct_bufchan_buf <= trae3_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (traeb_destruct,Pointer_QTree_Int) > (traeb_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t traeb_destruct_bufchan_d;
  logic traeb_destruct_bufchan_r;
  assign traeb_destruct_r = ((! traeb_destruct_bufchan_d[0]) || traeb_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) traeb_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (traeb_destruct_r) traeb_destruct_bufchan_d <= traeb_destruct_d;
  Pointer_QTree_Int_t traeb_destruct_bufchan_buf;
  assign traeb_destruct_bufchan_r = (! traeb_destruct_bufchan_buf[0]);
  assign traeb_1_argbuf_d = (traeb_destruct_bufchan_buf[0] ? traeb_destruct_bufchan_buf :
                             traeb_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) traeb_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((traeb_1_argbuf_r && traeb_destruct_bufchan_buf[0]))
        traeb_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! traeb_1_argbuf_r) && (! traeb_destruct_bufchan_buf[0])))
        traeb_destruct_bufchan_buf <= traeb_destruct_bufchan_d;
  
  /* destruct (Ty Int,Dcon I#) : (va8v_1I#,Int) > [(xakK_destruct,Int#)] */
  assign xakK_destruct_d = {\va8v_1I#_d [32:1], \va8v_1I#_d [0]};
  assign \va8v_1I#_r  = xakK_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (va8v_2,Int) (va8v_1,Int) > [(va8v_1I#,Int)] */
  assign \va8v_1I#_d  = {va8v_1_d[32:1],
                         (va8v_2_d[0] && va8v_1_d[0])};
  assign va8v_1_r = (\va8v_1I#_r  && (va8v_2_d[0] && va8v_1_d[0]));
  assign va8v_2_r = (\va8v_1I#_r  && (va8v_2_d[0] && va8v_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (va8v_3,Int) (lizzieLet3_3QVal_Int,Go) > [(va8v_3I#,Go)] */
  assign \va8v_3I#_d  = (va8v_3_d[0] && lizzieLet3_3QVal_Int_d[0]);
  assign lizzieLet3_3QVal_Int_r = (\va8v_3I#_r  && (va8v_3_d[0] && lizzieLet3_3QVal_Int_d[0]));
  assign va8v_3_r = (\va8v_3I#_r  && (va8v_3_d[0] && lizzieLet3_3QVal_Int_d[0]));
  
  /* fork (Ty Go) : (va8v_3I#,Go) > [(va8v_3I#_1,Go),
                                (va8v_3I#_2,Go),
                                (va8v_3I#_3,Go)] */
  logic [2:0] \va8v_3I#_emitted ;
  logic [2:0] \va8v_3I#_done ;
  assign \va8v_3I#_1_d  = (\va8v_3I#_d [0] && (! \va8v_3I#_emitted [0]));
  assign \va8v_3I#_2_d  = (\va8v_3I#_d [0] && (! \va8v_3I#_emitted [1]));
  assign \va8v_3I#_3_d  = (\va8v_3I#_d [0] && (! \va8v_3I#_emitted [2]));
  assign \va8v_3I#_done  = (\va8v_3I#_emitted  | ({\va8v_3I#_3_d [0],
                                                   \va8v_3I#_2_d [0],
                                                   \va8v_3I#_1_d [0]} & {\va8v_3I#_3_r ,
                                                                         \va8v_3I#_2_r ,
                                                                         \va8v_3I#_1_r }));
  assign \va8v_3I#_r  = (& \va8v_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \va8v_3I#_emitted  <= 3'd0;
    else
      \va8v_3I#_emitted  <= (\va8v_3I#_r  ? 3'd0 :
                             \va8v_3I#_done );
  
  /* buf (Ty Go) : (va8v_3I#_1,Go) > (va8v_3I#_1_argbuf,Go) */
  Go_t \va8v_3I#_1_bufchan_d ;
  logic \va8v_3I#_1_bufchan_r ;
  assign \va8v_3I#_1_r  = ((! \va8v_3I#_1_bufchan_d [0]) || \va8v_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \va8v_3I#_1_bufchan_d  <= 1'd0;
    else if (\va8v_3I#_1_r ) \va8v_3I#_1_bufchan_d  <= \va8v_3I#_1_d ;
  Go_t \va8v_3I#_1_bufchan_buf ;
  assign \va8v_3I#_1_bufchan_r  = (! \va8v_3I#_1_bufchan_buf [0]);
  assign \va8v_3I#_1_argbuf_d  = (\va8v_3I#_1_bufchan_buf [0] ? \va8v_3I#_1_bufchan_buf  :
                                  \va8v_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \va8v_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\va8v_3I#_1_argbuf_r  && \va8v_3I#_1_bufchan_buf [0]))
        \va8v_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \va8v_3I#_1_argbuf_r ) && (! \va8v_3I#_1_bufchan_buf [0])))
        \va8v_3I#_1_bufchan_buf  <= \va8v_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (va8v_3I#_1_argbuf,Go) > (va8v_3I#_1_argbuf_0,Int#) */
  assign \va8v_3I#_1_argbuf_0_d  = {32'd0, \va8v_3I#_1_argbuf_d [0]};
  assign \va8v_3I#_1_argbuf_r  = \va8v_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (va8v_3I#_1_argbuf_0,Int#) (xakK_destruct,Int#) > (lizzieLet5_1wild2XE_1_Eq,Bool) */
  assign lizzieLet5_1wild2XE_1_Eq_d = {(\va8v_3I#_1_argbuf_0_d [32:1] == xakK_destruct_d[32:1]),
                                       (\va8v_3I#_1_argbuf_0_d [0] && xakK_destruct_d[0])};
  assign {\va8v_3I#_1_argbuf_0_r ,
          xakK_destruct_r} = {2 {(lizzieLet5_1wild2XE_1_Eq_r && lizzieLet5_1wild2XE_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (va8v_3I#_2,Go) > (va8v_3I#_2_argbuf,Go) */
  Go_t \va8v_3I#_2_bufchan_d ;
  logic \va8v_3I#_2_bufchan_r ;
  assign \va8v_3I#_2_r  = ((! \va8v_3I#_2_bufchan_d [0]) || \va8v_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \va8v_3I#_2_bufchan_d  <= 1'd0;
    else if (\va8v_3I#_2_r ) \va8v_3I#_2_bufchan_d  <= \va8v_3I#_2_d ;
  Go_t \va8v_3I#_2_bufchan_buf ;
  assign \va8v_3I#_2_bufchan_r  = (! \va8v_3I#_2_bufchan_buf [0]);
  assign \va8v_3I#_2_argbuf_d  = (\va8v_3I#_2_bufchan_buf [0] ? \va8v_3I#_2_bufchan_buf  :
                                  \va8v_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \va8v_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\va8v_3I#_2_argbuf_r  && \va8v_3I#_2_bufchan_buf [0]))
        \va8v_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \va8v_3I#_2_argbuf_r ) && (! \va8v_3I#_2_bufchan_buf [0])))
        \va8v_3I#_2_bufchan_buf  <= \va8v_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,Dcon TupGo___Bool) : [(va8v_3I#_2_argbuf,Go),
                                            (lizzieLet6_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\va8v_3I#_2_argbuf_d [0],
                                                             lizzieLet6_1_argbuf_d[0]}), \va8v_3I#_2_argbuf_d , lizzieLet6_1_argbuf_d);
  assign {\va8v_3I#_2_argbuf_r ,
          lizzieLet6_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* demux (Ty Int,
       Ty Pointer_CTf''''''''_f'''''''') : (va8v_4,Int) (lizzieLet3_4QVal_Int,Pointer_CTf''''''''_f'''''''') > [(va8v_4I#,Pointer_CTf''''''''_f'''''''')] */
  assign \va8v_4I#_d  = {lizzieLet3_4QVal_Int_d[16:1],
                         (va8v_4_d[0] && lizzieLet3_4QVal_Int_d[0])};
  assign lizzieLet3_4QVal_Int_r = (\va8v_4I#_r  && (va8v_4_d[0] && lizzieLet3_4QVal_Int_d[0]));
  assign va8v_4_r = (\va8v_4I#_r  && (va8v_4_d[0] && lizzieLet3_4QVal_Int_d[0]));
  
  /* fork (Ty Int) : (va8v_destruct,Int) > [(va8v_1,Int),
                                       (va8v_2,Int),
                                       (va8v_3,Int),
                                       (va8v_4,Int)] */
  logic [3:0] va8v_destruct_emitted;
  logic [3:0] va8v_destruct_done;
  assign va8v_1_d = {va8v_destruct_d[32:1],
                     (va8v_destruct_d[0] && (! va8v_destruct_emitted[0]))};
  assign va8v_2_d = {va8v_destruct_d[32:1],
                     (va8v_destruct_d[0] && (! va8v_destruct_emitted[1]))};
  assign va8v_3_d = {va8v_destruct_d[32:1],
                     (va8v_destruct_d[0] && (! va8v_destruct_emitted[2]))};
  assign va8v_4_d = {va8v_destruct_d[32:1],
                     (va8v_destruct_d[0] && (! va8v_destruct_emitted[3]))};
  assign va8v_destruct_done = (va8v_destruct_emitted | ({va8v_4_d[0],
                                                         va8v_3_d[0],
                                                         va8v_2_d[0],
                                                         va8v_1_d[0]} & {va8v_4_r,
                                                                         va8v_3_r,
                                                                         va8v_2_r,
                                                                         va8v_1_r}));
  assign va8v_destruct_r = (& va8v_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8v_destruct_emitted <= 4'd0;
    else
      va8v_destruct_emitted <= (va8v_destruct_r ? 4'd0 :
                                va8v_destruct_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (vae8_1I#,Int) > [(xakK_1_destruct,Int#)] */
  assign xakK_1_destruct_d = {\vae8_1I#_d [32:1], \vae8_1I#_d [0]};
  assign \vae8_1I#_r  = xakK_1_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (vae8_2,Int) (vae8_1,Int) > [(vae8_1I#,Int)] */
  assign \vae8_1I#_d  = {vae8_1_d[32:1],
                         (vae8_2_d[0] && vae8_1_d[0])};
  assign vae8_1_r = (\vae8_1I#_r  && (vae8_2_d[0] && vae8_1_d[0]));
  assign vae8_2_r = (\vae8_1I#_r  && (vae8_2_d[0] && vae8_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (vae8_3,Int) (lizzieLet12_4QNone_Int_3QVal_Int,Go) > [(vae8_3I#,Go)] */
  assign \vae8_3I#_d  = (vae8_3_d[0] && lizzieLet12_4QNone_Int_3QVal_Int_d[0]);
  assign lizzieLet12_4QNone_Int_3QVal_Int_r = (\vae8_3I#_r  && (vae8_3_d[0] && lizzieLet12_4QNone_Int_3QVal_Int_d[0]));
  assign vae8_3_r = (\vae8_3I#_r  && (vae8_3_d[0] && lizzieLet12_4QNone_Int_3QVal_Int_d[0]));
  
  /* fork (Ty Go) : (vae8_3I#,Go) > [(vae8_3I#_1,Go),
                                (vae8_3I#_2,Go),
                                (vae8_3I#_3,Go)] */
  logic [2:0] \vae8_3I#_emitted ;
  logic [2:0] \vae8_3I#_done ;
  assign \vae8_3I#_1_d  = (\vae8_3I#_d [0] && (! \vae8_3I#_emitted [0]));
  assign \vae8_3I#_2_d  = (\vae8_3I#_d [0] && (! \vae8_3I#_emitted [1]));
  assign \vae8_3I#_3_d  = (\vae8_3I#_d [0] && (! \vae8_3I#_emitted [2]));
  assign \vae8_3I#_done  = (\vae8_3I#_emitted  | ({\vae8_3I#_3_d [0],
                                                   \vae8_3I#_2_d [0],
                                                   \vae8_3I#_1_d [0]} & {\vae8_3I#_3_r ,
                                                                         \vae8_3I#_2_r ,
                                                                         \vae8_3I#_1_r }));
  assign \vae8_3I#_r  = (& \vae8_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \vae8_3I#_emitted  <= 3'd0;
    else
      \vae8_3I#_emitted  <= (\vae8_3I#_r  ? 3'd0 :
                             \vae8_3I#_done );
  
  /* buf (Ty Go) : (vae8_3I#_1,Go) > (vae8_3I#_1_argbuf,Go) */
  Go_t \vae8_3I#_1_bufchan_d ;
  logic \vae8_3I#_1_bufchan_r ;
  assign \vae8_3I#_1_r  = ((! \vae8_3I#_1_bufchan_d [0]) || \vae8_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \vae8_3I#_1_bufchan_d  <= 1'd0;
    else if (\vae8_3I#_1_r ) \vae8_3I#_1_bufchan_d  <= \vae8_3I#_1_d ;
  Go_t \vae8_3I#_1_bufchan_buf ;
  assign \vae8_3I#_1_bufchan_r  = (! \vae8_3I#_1_bufchan_buf [0]);
  assign \vae8_3I#_1_argbuf_d  = (\vae8_3I#_1_bufchan_buf [0] ? \vae8_3I#_1_bufchan_buf  :
                                  \vae8_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \vae8_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\vae8_3I#_1_argbuf_r  && \vae8_3I#_1_bufchan_buf [0]))
        \vae8_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \vae8_3I#_1_argbuf_r ) && (! \vae8_3I#_1_bufchan_buf [0])))
        \vae8_3I#_1_bufchan_buf  <= \vae8_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (vae8_3I#_1_argbuf,Go) > (vae8_3I#_1_argbuf_0,Int#) */
  assign \vae8_3I#_1_argbuf_0_d  = {32'd0, \vae8_3I#_1_argbuf_d [0]};
  assign \vae8_3I#_1_argbuf_r  = \vae8_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (vae8_3I#_1_argbuf_0,Int#) (xakK_1_destruct,Int#) > (lizzieLet15_1wild3XR_1_Eq,Bool) */
  assign lizzieLet15_1wild3XR_1_Eq_d = {(\vae8_3I#_1_argbuf_0_d [32:1] == xakK_1_destruct_d[32:1]),
                                        (\vae8_3I#_1_argbuf_0_d [0] && xakK_1_destruct_d[0])};
  assign {\vae8_3I#_1_argbuf_0_r ,
          xakK_1_destruct_r} = {2 {(lizzieLet15_1wild3XR_1_Eq_r && lizzieLet15_1wild3XR_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (vae8_3I#_2,Go) > (vae8_3I#_2_argbuf,Go) */
  Go_t \vae8_3I#_2_bufchan_d ;
  logic \vae8_3I#_2_bufchan_r ;
  assign \vae8_3I#_2_r  = ((! \vae8_3I#_2_bufchan_d [0]) || \vae8_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \vae8_3I#_2_bufchan_d  <= 1'd0;
    else if (\vae8_3I#_2_r ) \vae8_3I#_2_bufchan_d  <= \vae8_3I#_2_d ;
  Go_t \vae8_3I#_2_bufchan_buf ;
  assign \vae8_3I#_2_bufchan_r  = (! \vae8_3I#_2_bufchan_buf [0]);
  assign \vae8_3I#_2_argbuf_d  = (\vae8_3I#_2_bufchan_buf [0] ? \vae8_3I#_2_bufchan_buf  :
                                  \vae8_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \vae8_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\vae8_3I#_2_argbuf_r  && \vae8_3I#_2_bufchan_buf [0]))
        \vae8_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \vae8_3I#_2_argbuf_r ) && (! \vae8_3I#_2_bufchan_buf [0])))
        \vae8_3I#_2_bufchan_buf  <= \vae8_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,Dcon TupGo___Bool) : [(vae8_3I#_2_argbuf,Go),
                                            (lizzieLet16_1_argbuf,Bool)] > (boolConvert_2TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_2TupGo___Bool_1_d = TupGo___Bool_dc((& {\vae8_3I#_2_argbuf_d [0],
                                                             lizzieLet16_1_argbuf_d[0]}), \vae8_3I#_2_argbuf_d , lizzieLet16_1_argbuf_d);
  assign {\vae8_3I#_2_argbuf_r ,
          lizzieLet16_1_argbuf_r} = {2 {(boolConvert_2TupGo___Bool_1_r && boolConvert_2TupGo___Bool_1_d[0])}};
  
  /* demux (Ty Int,
       Ty Pointer_CTf_f) : (vae8_4,Int) (lizzieLet12_4QNone_Int_4QVal_Int,Pointer_CTf_f) > [(vae8_4I#,Pointer_CTf_f)] */
  assign \vae8_4I#_d  = {lizzieLet12_4QNone_Int_4QVal_Int_d[16:1],
                         (vae8_4_d[0] && lizzieLet12_4QNone_Int_4QVal_Int_d[0])};
  assign lizzieLet12_4QNone_Int_4QVal_Int_r = (\vae8_4I#_r  && (vae8_4_d[0] && lizzieLet12_4QNone_Int_4QVal_Int_d[0]));
  assign vae8_4_r = (\vae8_4I#_r  && (vae8_4_d[0] && lizzieLet12_4QNone_Int_4QVal_Int_d[0]));
  
  /* fork (Ty Int) : (vae8_destruct,Int) > [(vae8_1,Int),
                                       (vae8_2,Int),
                                       (vae8_3,Int),
                                       (vae8_4,Int)] */
  logic [3:0] vae8_destruct_emitted;
  logic [3:0] vae8_destruct_done;
  assign vae8_1_d = {vae8_destruct_d[32:1],
                     (vae8_destruct_d[0] && (! vae8_destruct_emitted[0]))};
  assign vae8_2_d = {vae8_destruct_d[32:1],
                     (vae8_destruct_d[0] && (! vae8_destruct_emitted[1]))};
  assign vae8_3_d = {vae8_destruct_d[32:1],
                     (vae8_destruct_d[0] && (! vae8_destruct_emitted[2]))};
  assign vae8_4_d = {vae8_destruct_d[32:1],
                     (vae8_destruct_d[0] && (! vae8_destruct_emitted[3]))};
  assign vae8_destruct_done = (vae8_destruct_emitted | ({vae8_4_d[0],
                                                         vae8_3_d[0],
                                                         vae8_2_d[0],
                                                         vae8_1_d[0]} & {vae8_4_r,
                                                                         vae8_3_r,
                                                                         vae8_2_r,
                                                                         vae8_1_r}));
  assign vae8_destruct_r = (& vae8_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vae8_destruct_emitted <= 4'd0;
    else
      vae8_destruct_emitted <= (vae8_destruct_r ? 4'd0 :
                                vae8_destruct_done);
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_r)
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet0_1_argbuf_rwb_r && writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz) > (lizzieLet20_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet2_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet2_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet2_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet2_1_argbuf_r = ((! writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet2_1_argbuf_r)
        writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet2_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet2_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet2_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet2_1_argbuf_rwb_r && writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet2_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet2_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet2_1_argbuf_rwb,Pointer_CT$wnnz) > (sca3_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet2_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet2_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet2_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet45_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet45_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet45_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet45_1_argbuf_r = ((! writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet45_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet45_1_argbuf_r)
        writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet45_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet45_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet45_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet45_1_argbuf_rwb_r && writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet45_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet45_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet45_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet45_1_argbuf_rwb,Pointer_CT$wnnz) > (sca2_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet45_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet45_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet45_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet45_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet46_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet46_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet46_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet46_1_argbuf_r = ((! writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet46_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet46_1_argbuf_r)
        writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet46_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet46_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet46_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet46_1_argbuf_rwb_r && writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet46_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet46_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet46_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet46_1_argbuf_rwb,Pointer_CT$wnnz) > (sca1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet46_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet46_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet46_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet46_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet47_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet47_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet47_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet47_1_argbuf_r = ((! writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet47_1_argbuf_r)
        writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet47_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet47_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet47_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet47_1_argbuf_rwb_r && writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet47_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet47_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet47_1_argbuf_rwb,Pointer_CT$wnnz) > (sca0_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet47_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet47_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet47_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet10_1_argbuf,Pointer_CTf''''''''_f'''''''') > (writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d  <= {16'd0,
                                                                     1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_r )
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf  :
                                                                   \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
    else
      if ((\writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
      else if (((! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') > (sca3_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet10_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet42_1_argbuf,Pointer_CTf''''''''_f'''''''') > (writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d  <= {16'd0,
                                                                     1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_r )
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf  :
                                                                   \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
    else
      if ((\writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
      else if (((! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') > (lizzieLet4_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet4_1_1_argbuf_d = (\writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet42_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet49_1_argbuf,Pointer_CTf''''''''_f'''''''') > (writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d  <= {16'd0,
                                                                     1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_r )
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf  :
                                                                   \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
    else
      if ((\writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
      else if (((! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') > (sca2_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet49_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet50_1_argbuf,Pointer_CTf''''''''_f'''''''') > (writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d  <= {16'd0,
                                                                     1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_r )
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf  :
                                                                   \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
    else
      if ((\writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
      else if (((! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') > (sca1_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet50_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet51_1_argbuf,Pointer_CTf''''''''_f'''''''') > (writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_r  = ((! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d  <= {16'd0,
                                                                     1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_r )
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf [0]);
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_d  = (\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf  :
                                                                   \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf  <= {16'd0,
                                                                       1'd0};
    else
      if ((\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_r  && \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
      else if (((! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_r ) && (! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf''''''''_f'''''''') : (writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb,Pointer_CTf''''''''_f'''''''') > (sca0_1_1_argbuf,Pointer_CTf''''''''_f'''''''') */
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_r  = ((! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d [0]) || \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_r )
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d  <= \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_d ;
  \Pointer_CTf''''''''_f''''''''_t  \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_r  = (! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_buf  <= \writeCTf''''''''_f''''''''lizzieLet51_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet38_1_argbuf,Pointer_CTf_f) > (writeCTf_flizzieLet38_1_argbuf_rwb,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_bufchan_d;
  logic writeCTf_flizzieLet38_1_argbuf_bufchan_r;
  assign writeCTf_flizzieLet38_1_argbuf_r = ((! writeCTf_flizzieLet38_1_argbuf_bufchan_d[0]) || writeCTf_flizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet38_1_argbuf_r)
        writeCTf_flizzieLet38_1_argbuf_bufchan_d <= writeCTf_flizzieLet38_1_argbuf_d;
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_bufchan_buf;
  assign writeCTf_flizzieLet38_1_argbuf_bufchan_r = (! writeCTf_flizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeCTf_flizzieLet38_1_argbuf_rwb_d = (writeCTf_flizzieLet38_1_argbuf_bufchan_buf[0] ? writeCTf_flizzieLet38_1_argbuf_bufchan_buf :
                                                 writeCTf_flizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_flizzieLet38_1_argbuf_rwb_r && writeCTf_flizzieLet38_1_argbuf_bufchan_buf[0]))
        writeCTf_flizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_flizzieLet38_1_argbuf_rwb_r) && (! writeCTf_flizzieLet38_1_argbuf_bufchan_buf[0])))
        writeCTf_flizzieLet38_1_argbuf_bufchan_buf <= writeCTf_flizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet38_1_argbuf_rwb,Pointer_CTf_f) > (sca3_2_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeCTf_flizzieLet38_1_argbuf_rwb_r = ((! writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet38_1_argbuf_rwb_r)
        writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d <= writeCTf_flizzieLet38_1_argbuf_rwb_d;
  Pointer_CTf_f_t writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_r = (! writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf :
                              writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_buf <= writeCTf_flizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet43_1_argbuf,Pointer_CTf_f) > (writeCTf_flizzieLet43_1_argbuf_rwb,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_bufchan_d;
  logic writeCTf_flizzieLet43_1_argbuf_bufchan_r;
  assign writeCTf_flizzieLet43_1_argbuf_r = ((! writeCTf_flizzieLet43_1_argbuf_bufchan_d[0]) || writeCTf_flizzieLet43_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet43_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet43_1_argbuf_r)
        writeCTf_flizzieLet43_1_argbuf_bufchan_d <= writeCTf_flizzieLet43_1_argbuf_d;
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_bufchan_buf;
  assign writeCTf_flizzieLet43_1_argbuf_bufchan_r = (! writeCTf_flizzieLet43_1_argbuf_bufchan_buf[0]);
  assign writeCTf_flizzieLet43_1_argbuf_rwb_d = (writeCTf_flizzieLet43_1_argbuf_bufchan_buf[0] ? writeCTf_flizzieLet43_1_argbuf_bufchan_buf :
                                                 writeCTf_flizzieLet43_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_flizzieLet43_1_argbuf_rwb_r && writeCTf_flizzieLet43_1_argbuf_bufchan_buf[0]))
        writeCTf_flizzieLet43_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_flizzieLet43_1_argbuf_rwb_r) && (! writeCTf_flizzieLet43_1_argbuf_bufchan_buf[0])))
        writeCTf_flizzieLet43_1_argbuf_bufchan_buf <= writeCTf_flizzieLet43_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet43_1_argbuf_rwb,Pointer_CTf_f) > (lizzieLet17_1_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d;
  logic writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_r;
  assign writeCTf_flizzieLet43_1_argbuf_rwb_r = ((! writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d[0]) || writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet43_1_argbuf_rwb_r)
        writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d <= writeCTf_flizzieLet43_1_argbuf_rwb_d;
  Pointer_CTf_f_t writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_r = (! writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf :
                                     writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_buf <= writeCTf_flizzieLet43_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet54_1_argbuf,Pointer_CTf_f) > (writeCTf_flizzieLet54_1_argbuf_rwb,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_bufchan_d;
  logic writeCTf_flizzieLet54_1_argbuf_bufchan_r;
  assign writeCTf_flizzieLet54_1_argbuf_r = ((! writeCTf_flizzieLet54_1_argbuf_bufchan_d[0]) || writeCTf_flizzieLet54_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet54_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet54_1_argbuf_r)
        writeCTf_flizzieLet54_1_argbuf_bufchan_d <= writeCTf_flizzieLet54_1_argbuf_d;
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_bufchan_buf;
  assign writeCTf_flizzieLet54_1_argbuf_bufchan_r = (! writeCTf_flizzieLet54_1_argbuf_bufchan_buf[0]);
  assign writeCTf_flizzieLet54_1_argbuf_rwb_d = (writeCTf_flizzieLet54_1_argbuf_bufchan_buf[0] ? writeCTf_flizzieLet54_1_argbuf_bufchan_buf :
                                                 writeCTf_flizzieLet54_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_flizzieLet54_1_argbuf_rwb_r && writeCTf_flizzieLet54_1_argbuf_bufchan_buf[0]))
        writeCTf_flizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_flizzieLet54_1_argbuf_rwb_r) && (! writeCTf_flizzieLet54_1_argbuf_bufchan_buf[0])))
        writeCTf_flizzieLet54_1_argbuf_bufchan_buf <= writeCTf_flizzieLet54_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet54_1_argbuf_rwb,Pointer_CTf_f) > (sca2_2_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d;
  logic writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_r;
  assign writeCTf_flizzieLet54_1_argbuf_rwb_r = ((! writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d[0]) || writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet54_1_argbuf_rwb_r)
        writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d <= writeCTf_flizzieLet54_1_argbuf_rwb_d;
  Pointer_CTf_f_t writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_r = (! writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf :
                              writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_buf <= writeCTf_flizzieLet54_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet55_1_argbuf,Pointer_CTf_f) > (writeCTf_flizzieLet55_1_argbuf_rwb,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_bufchan_d;
  logic writeCTf_flizzieLet55_1_argbuf_bufchan_r;
  assign writeCTf_flizzieLet55_1_argbuf_r = ((! writeCTf_flizzieLet55_1_argbuf_bufchan_d[0]) || writeCTf_flizzieLet55_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet55_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet55_1_argbuf_r)
        writeCTf_flizzieLet55_1_argbuf_bufchan_d <= writeCTf_flizzieLet55_1_argbuf_d;
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_bufchan_buf;
  assign writeCTf_flizzieLet55_1_argbuf_bufchan_r = (! writeCTf_flizzieLet55_1_argbuf_bufchan_buf[0]);
  assign writeCTf_flizzieLet55_1_argbuf_rwb_d = (writeCTf_flizzieLet55_1_argbuf_bufchan_buf[0] ? writeCTf_flizzieLet55_1_argbuf_bufchan_buf :
                                                 writeCTf_flizzieLet55_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_flizzieLet55_1_argbuf_rwb_r && writeCTf_flizzieLet55_1_argbuf_bufchan_buf[0]))
        writeCTf_flizzieLet55_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_flizzieLet55_1_argbuf_rwb_r) && (! writeCTf_flizzieLet55_1_argbuf_bufchan_buf[0])))
        writeCTf_flizzieLet55_1_argbuf_bufchan_buf <= writeCTf_flizzieLet55_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet55_1_argbuf_rwb,Pointer_CTf_f) > (sca1_2_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d;
  logic writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_r;
  assign writeCTf_flizzieLet55_1_argbuf_rwb_r = ((! writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d[0]) || writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet55_1_argbuf_rwb_r)
        writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d <= writeCTf_flizzieLet55_1_argbuf_rwb_d;
  Pointer_CTf_f_t writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_r = (! writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf :
                              writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_buf <= writeCTf_flizzieLet55_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet56_1_argbuf,Pointer_CTf_f) > (writeCTf_flizzieLet56_1_argbuf_rwb,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_bufchan_d;
  logic writeCTf_flizzieLet56_1_argbuf_bufchan_r;
  assign writeCTf_flizzieLet56_1_argbuf_r = ((! writeCTf_flizzieLet56_1_argbuf_bufchan_d[0]) || writeCTf_flizzieLet56_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet56_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet56_1_argbuf_r)
        writeCTf_flizzieLet56_1_argbuf_bufchan_d <= writeCTf_flizzieLet56_1_argbuf_d;
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_bufchan_buf;
  assign writeCTf_flizzieLet56_1_argbuf_bufchan_r = (! writeCTf_flizzieLet56_1_argbuf_bufchan_buf[0]);
  assign writeCTf_flizzieLet56_1_argbuf_rwb_d = (writeCTf_flizzieLet56_1_argbuf_bufchan_buf[0] ? writeCTf_flizzieLet56_1_argbuf_bufchan_buf :
                                                 writeCTf_flizzieLet56_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet56_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_flizzieLet56_1_argbuf_rwb_r && writeCTf_flizzieLet56_1_argbuf_bufchan_buf[0]))
        writeCTf_flizzieLet56_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_flizzieLet56_1_argbuf_rwb_r) && (! writeCTf_flizzieLet56_1_argbuf_bufchan_buf[0])))
        writeCTf_flizzieLet56_1_argbuf_bufchan_buf <= writeCTf_flizzieLet56_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f) : (writeCTf_flizzieLet56_1_argbuf_rwb,Pointer_CTf_f) > (sca0_2_1_argbuf,Pointer_CTf_f) */
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d;
  logic writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_r;
  assign writeCTf_flizzieLet56_1_argbuf_rwb_r = ((! writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d[0]) || writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_flizzieLet56_1_argbuf_rwb_r)
        writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d <= writeCTf_flizzieLet56_1_argbuf_rwb_d;
  Pointer_CTf_f_t writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_r = (! writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf :
                              writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_buf <= writeCTf_flizzieLet56_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet11_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_argbuf_r = ((! writeQTree_BoollizzieLet11_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_argbuf_r)
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet11_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_d = (writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet11_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet11_1_argbuf_rwb_r && writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet11_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet11_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet11_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet11_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet11_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet11_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_r = ((! writeQTree_BoollizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_r)
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_d = (writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet14_1_argbuf_rwb_r && writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet14_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet19_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_1_argbuf_r = ((! writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_1_argbuf_r)
        writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet19_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet19_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet19_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet19_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet19_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet19_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet19_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet20_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet20_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet20_1_1_argbuf_r = ((! writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet20_1_1_argbuf_r)
        writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet20_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet20_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet20_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet20_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet20_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet20_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet20_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet20_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet20_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet20_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet21_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet21_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet21_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet21_1_argbuf_r = ((! writeQTree_BoollizzieLet21_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet21_1_argbuf_r)
        writeQTree_BoollizzieLet21_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet21_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet21_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet21_1_argbuf_rwb_d = (writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet21_1_argbuf_rwb_r && writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet21_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet21_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet21_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet21_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet21_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet21_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet27_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet27_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet27_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet27_1_argbuf_r = ((! writeQTree_BoollizzieLet27_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet27_1_argbuf_r)
        writeQTree_BoollizzieLet27_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet27_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet27_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet27_1_argbuf_rwb_d = (writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet27_1_argbuf_rwb_r && writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet27_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet27_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet27_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet27_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet27_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet27_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet32_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet32_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet32_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet32_1_argbuf_r = ((! writeQTree_BoollizzieLet32_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet32_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet32_1_argbuf_r)
        writeQTree_BoollizzieLet32_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet32_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet32_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet32_1_argbuf_rwb_d = (writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet32_1_argbuf_rwb_r && writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet32_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet32_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet32_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet10_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet32_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet32_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet32_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet33_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet33_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet33_1_argbuf_r = ((! writeQTree_BoollizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet33_1_argbuf_r)
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet33_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet33_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_d = (writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet33_1_argbuf_rwb_r && writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet33_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet33_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet33_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet11_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet33_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_r = ((! writeQTree_BoollizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_r)
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_d = (writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet34_1_argbuf_rwb_r && writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet34_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet34_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet12_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet34_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_r = ((! writeQTree_BoollizzieLet36_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_r)
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_d = (writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet36_1_argbuf_rwb_r && writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet36_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet36_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet13_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet36_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet36_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_r = ((! writeQTree_BoollizzieLet37_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_r)
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_d = (writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet37_1_argbuf_rwb_r && writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet37_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet14_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet39_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet39_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet39_1_argbuf_r = ((! writeQTree_BoollizzieLet39_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet39_1_argbuf_r)
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet39_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet39_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_d = (writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet39_1_argbuf_rwb_r && writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet39_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet39_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet39_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet39_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet15_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet39_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet39_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet39_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet40_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet40_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet40_1_argbuf_r = ((! writeQTree_BoollizzieLet40_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet40_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet40_1_argbuf_r)
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet40_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet40_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_d = (writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet40_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet40_1_argbuf_rwb_r && writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet40_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet40_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet40_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet40_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet16_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet40_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet40_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet40_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet41_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet41_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet41_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet41_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet41_1_argbuf_r = ((! writeQTree_BoollizzieLet41_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet41_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet41_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet41_1_argbuf_r)
        writeQTree_BoollizzieLet41_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet41_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet41_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet41_1_argbuf_rwb_d = (writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet41_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet41_1_argbuf_rwb_r && writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet41_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet41_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet41_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_r = ((! writeQTree_BoollizzieLet4_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_r)
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_d = (writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet4_1_argbuf_rwb_r && writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet4_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet52_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet52_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet52_1_argbuf_r = ((! writeQTree_BoollizzieLet52_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet52_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet52_1_argbuf_r)
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet52_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet52_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_d = (writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet52_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet52_1_argbuf_rwb_r && writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet52_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet52_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet52_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet52_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet52_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet52_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet52_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet57_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet57_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet57_1_argbuf_r = ((! writeQTree_BoollizzieLet57_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet57_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet57_1_argbuf_r)
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet57_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet57_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_d = (writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet57_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet57_1_argbuf_rwb_r && writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet57_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet57_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet57_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet57_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet57_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet57_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet57_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet9_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_argbuf_r = ((! writeQTree_BoollizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_argbuf_r)
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet9_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_d = (writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet9_1_argbuf_rwb_r && writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet9_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (wspF_1_goMux_mux,Pointer_QTree_Bool) > (wspF_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t wspF_1_goMux_mux_bufchan_d;
  logic wspF_1_goMux_mux_bufchan_r;
  assign wspF_1_goMux_mux_r = ((! wspF_1_goMux_mux_bufchan_d[0]) || wspF_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wspF_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wspF_1_goMux_mux_r)
        wspF_1_goMux_mux_bufchan_d <= wspF_1_goMux_mux_d;
  Pointer_QTree_Bool_t wspF_1_goMux_mux_bufchan_buf;
  assign wspF_1_goMux_mux_bufchan_r = (! wspF_1_goMux_mux_bufchan_buf[0]);
  assign wspF_1_1_argbuf_d = (wspF_1_goMux_mux_bufchan_buf[0] ? wspF_1_goMux_mux_bufchan_buf :
                              wspF_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wspF_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wspF_1_1_argbuf_r && wspF_1_goMux_mux_bufchan_buf[0]))
        wspF_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wspF_1_1_argbuf_r) && (! wspF_1_goMux_mux_bufchan_buf[0])))
        wspF_1_goMux_mux_bufchan_buf <= wspF_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1,CT$wnnz) > (lizzieLet46_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d;
  logic wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r;
  assign wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r = ((! wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d[0]) || wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r)
        wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d <= wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d;
  CT$wnnz_t wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf;
  assign wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_r = (! wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet46_1_argbuf_d = (wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0] ? wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf :
                                   wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet46_1_argbuf_r && wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0]))
        wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet46_1_argbuf_r) && (! wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf[0])))
        wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_buf <= wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz1) : [(wwspI_2_destruct,Int#),
                                       (lizzieLet44_4Lcall_$wnnz2,Int#),
                                       (sc_0_4_destruct,Pointer_CT$wnnz),
                                       (q4a87_2_destruct,Pointer_QTree_Bool)] > (wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1,CT$wnnz) */
  assign wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d = Lcall_$wnnz1_dc((& {wwspI_2_destruct_d[0],
                                                                                                   lizzieLet44_4Lcall_$wnnz2_d[0],
                                                                                                   sc_0_4_destruct_d[0],
                                                                                                   q4a87_2_destruct_d[0]}), wwspI_2_destruct_d, lizzieLet44_4Lcall_$wnnz2_d, sc_0_4_destruct_d, q4a87_2_destruct_d);
  assign {wwspI_2_destruct_r,
          lizzieLet44_4Lcall_$wnnz2_r,
          sc_0_4_destruct_r,
          q4a87_2_destruct_r} = {4 {(wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_r && wwspI_2_1lizzieLet44_4Lcall_$wnnz2_1sc_0_4_1q4a87_2_1Lcall_$wnnz1_d[0])}};
  
  /* buf (Ty CT$wnnz) : (wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) > (lizzieLet47_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  logic wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r;
  assign wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r = ((! wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d[0]) || wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= {115'd0,
                                                                                       1'd0};
    else
      if (wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r)
        wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d <= wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d;
  CT$wnnz_t wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf;
  assign wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_r = (! wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0] ? wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf :
                                   wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0]))
        wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                           1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf[0])))
        wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_buf <= wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz0) : [(wwspI_3_destruct,Int#),
                                       (ww1Xqr_1_destruct,Int#),
                                       (lizzieLet44_4Lcall_$wnnz1,Int#),
                                       (sc_0_5_destruct,Pointer_CT$wnnz)] > (wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0,CT$wnnz) */
  assign wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d = Lcall_$wnnz0_dc((& {wwspI_3_destruct_d[0],
                                                                                                    ww1Xqr_1_destruct_d[0],
                                                                                                    lizzieLet44_4Lcall_$wnnz1_d[0],
                                                                                                    sc_0_5_destruct_d[0]}), wwspI_3_destruct_d, ww1Xqr_1_destruct_d, lizzieLet44_4Lcall_$wnnz1_d, sc_0_5_destruct_d);
  assign {wwspI_3_destruct_r,
          ww1Xqr_1_destruct_r,
          lizzieLet44_4Lcall_$wnnz1_r,
          sc_0_5_destruct_r} = {4 {(wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_r && wwspI_3_1ww1Xqr_1_1lizzieLet44_4Lcall_$wnnz1_1sc_0_5_1Lcall_$wnnz0_d[0])}};
  
  /* op_add (Ty Int#) : (wwspI_4_1ww1Xqr_2_1_Add32,Int#) (ww2Xqu_1_destruct,Int#) > (es_6_1_1ww2Xqu_1_1_Add32,Int#) */
  assign es_6_1_1ww2Xqu_1_1_Add32_d = {(wwspI_4_1ww1Xqr_2_1_Add32_d[32:1] + ww2Xqu_1_destruct_d[32:1]),
                                       (wwspI_4_1ww1Xqr_2_1_Add32_d[0] && ww2Xqu_1_destruct_d[0])};
  assign {wwspI_4_1ww1Xqr_2_1_Add32_r,
          ww2Xqu_1_destruct_r} = {2 {(es_6_1_1ww2Xqu_1_1_Add32_r && es_6_1_1ww2Xqu_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwspI_4_destruct,Int#) (ww1Xqr_2_destruct,Int#) > (wwspI_4_1ww1Xqr_2_1_Add32,Int#) */
  assign wwspI_4_1ww1Xqr_2_1_Add32_d = {(wwspI_4_destruct_d[32:1] + ww1Xqr_2_destruct_d[32:1]),
                                        (wwspI_4_destruct_d[0] && ww1Xqr_2_destruct_d[0])};
  assign {wwspI_4_destruct_r,
          ww1Xqr_2_destruct_r} = {2 {(wwspI_4_1ww1Xqr_2_1_Add32_r && wwspI_4_1ww1Xqr_2_1_Add32_d[0])}};
endmodule