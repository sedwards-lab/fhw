`timescale 1ns/1ns
import mMaskAdd_package::*;

module mMaskAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1a8v_0_d,
  output logic m1a8v_0_r,
  input Pointer_QTree_Int_t m2a8w_1_d,
  output logic m2a8w_1_r,
  input Pointer_QTree_Int_t m3a8x_2_d,
  output logic m3a8x_2_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Int_t \es_6_1I#_dout ,
  input logic \es_6_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1a8v_0, 16, 65536, Pointer_MaskQTree), (m2a8w_1, 16, 65536, Pointer_QTree_Int), (m3a8x_2, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (es_6_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTf__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
CTf__027_f__027_Int 16 3 (0,[0]) (1,[16p,16p,16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,0,0,16p,16p]) (3,[16p,16p,16p,16p,16p,0,0]) (4,[16p,16p,16p,16p])
CTf_f_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p,0,0,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,16p,16p,16p,0,0]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf__027__027__027__027__027__027__027__027__027_f__027__027__027__027__027__027__027__027__027_Int 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf__027_f__027_Int 16 0 (0,[0,16p,16p,0,0,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int 16 0 (0,[0,16p,16p,16p,0,0,16p])
TupGo___Pointer_MaskQTree___Pointer_QTree_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int 16 0 (0,[0,16p,16p,0,0])
TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int 16 0 (0,[0,16p,16p,16p,0,0])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  Go_t go__11_d;
  logic go__11_r;
  Go_t go__12_d;
  logic go__12_r;
  \Word16#_t  initHP_CT$wnnz_Int_d;
  logic initHP_CT$wnnz_Int_r;
  \Word16#_t  incrHP_CT$wnnz_Int_d;
  logic incrHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_d;
  logic incrHP_mergeCT$wnnz_Int_r;
  Go_t incrHP_CT$wnnz_Int1_d;
  logic incrHP_CT$wnnz_Int1_r;
  Go_t incrHP_CT$wnnz_Int2_d;
  logic incrHP_CT$wnnz_Int2_r;
  \Word16#_t  addHP_CT$wnnz_Int_d;
  logic addHP_CT$wnnz_Int_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_d;
  logic mergeHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_buf_d;
  logic incrHP_mergeCT$wnnz_Int_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_buf_d;
  logic mergeHP_CT$wnnz_Int_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_Int_d;
  logic forkHP1_CT$wnnz_Int_r;
  \Word16#_t  forkHP1_CT$wnnz_In2_d;
  logic forkHP1_CT$wnnz_In2_r;
  \Word16#_t  forkHP1_CT$wnnz_In3_d;
  logic forkHP1_CT$wnnz_In3_r;
  C2_t memMergeChoice_CT$wnnz_Int_d;
  logic memMergeChoice_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_d;
  logic memMergeIn_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_d;
  logic memOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memReadOut_CT$wnnz_Int_d;
  logic memReadOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memWriteOut_CT$wnnz_Int_d;
  logic memWriteOut_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_dbuf_d;
  logic memMergeIn_CT$wnnz_Int_dbuf_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_rbuf_d;
  logic memMergeIn_CT$wnnz_Int_rbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_dbuf_d;
  logic memOut_CT$wnnz_Int_dbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_rbuf_d;
  logic memOut_CT$wnnz_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_Int_d;
  logic destructReadIn_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t dconReadIn_CT$wnnz_Int_d;
  logic dconReadIn_CT$wnnz_Int_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_Int_d;
  logic writeMerge_choice_CT$wnnz_Int_r;
  CT$wnnz_Int_t writeMerge_data_CT$wnnz_Int_d;
  logic writeMerge_data_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet47_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet48_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet49_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_r;
  MemIn_CT$wnnz_Int_t dconWriteIn_CT$wnnz_Int_d;
  logic dconWriteIn_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t dconPtr_CT$wnnz_Int_d;
  logic dconPtr_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t _171_d;
  logic _171_r;
  assign _171_r = 1'd1;
  Pointer_CT$wnnz_Int_t demuxWriteResult_CT$wnnz_Int_d;
  logic demuxWriteResult_CT$wnnz_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C6_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm2ae4_1_argbuf_d;
  logic readPointer_QTree_Intm2ae4_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm2aeH_1_argbuf_d;
  logic readPointer_QTree_Intm2aeH_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm3ae5_1_argbuf_d;
  logic readPointer_QTree_Intm3ae5_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm3aeI_1_argbuf_d;
  logic readPointer_QTree_Intm3aeI_1_argbuf_r;
  QTree_Int_t \readPointer_QTree_Intq4'aex_1_argbuf_d ;
  logic \readPointer_QTree_Intq4'aex_1_argbuf_r ;
  QTree_Int_t readPointer_QTree_IntwsjQ_1_1_argbuf_d;
  logic readPointer_QTree_IntwsjQ_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C29_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_d;
  logic writeQTree_IntlizzieLet12_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_d;
  logic writeQTree_IntlizzieLet28_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet29_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet30_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet33_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_d;
  logic writeQTree_IntlizzieLet59_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_d;
  logic writeQTree_IntlizzieLet64_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _170_d;
  logic _170_r;
  assign _170_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  \initHP_CTf'''''''''_f'''''''''_Int_d ;
  logic \initHP_CTf'''''''''_f'''''''''_Int_r ;
  \Word16#_t  \incrHP_CTf'''''''''_f'''''''''_Int_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Int_r ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Int_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Int_r ;
  Go_t \incrHP_CTf'''''''''_f'''''''''_Int1_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Int1_r ;
  Go_t \incrHP_CTf'''''''''_f'''''''''_Int2_d ;
  logic \incrHP_CTf'''''''''_f'''''''''_Int2_r ;
  \Word16#_t  \addHP_CTf'''''''''_f'''''''''_Int_d ;
  logic \addHP_CTf'''''''''_f'''''''''_Int_r ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Int_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Int_r ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_r ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Int_buf_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Int_buf_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_Int_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_Int_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_In2_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_In2_r ;
  \Word16#_t  \forkHP1_CTf'''''''''_f'''''''''_In3_d ;
  logic \forkHP1_CTf'''''''''_f'''''''''_In3_r ;
  C2_t \memMergeChoice_CTf'''''''''_f'''''''''_Int_d ;
  logic \memMergeChoice_CTf'''''''''_f'''''''''_Int_r ;
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \memMergeIn_CTf'''''''''_f'''''''''_Int_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Int_r ;
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memOut_CTf'''''''''_f'''''''''_Int_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Int_r ;
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memReadOut_CTf'''''''''_f'''''''''_Int_d ;
  logic \memReadOut_CTf'''''''''_f'''''''''_Int_r ;
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memWriteOut_CTf'''''''''_f'''''''''_Int_d ;
  logic \memWriteOut_CTf'''''''''_f'''''''''_Int_r ;
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_r ;
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_d ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_r ;
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memOut_CTf'''''''''_f'''''''''_Int_dbuf_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Int_dbuf_r ;
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memOut_CTf'''''''''_f'''''''''_Int_rbuf_d ;
  logic \memOut_CTf'''''''''_f'''''''''_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf'''''''''_f'''''''''_Int_d ;
  logic \destructReadIn_CTf'''''''''_f'''''''''_Int_r ;
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \dconReadIn_CTf'''''''''_f'''''''''_Int_d ;
  logic \dconReadIn_CTf'''''''''_f'''''''''_Int_r ;
  \CTf'''''''''_f'''''''''_Int_t  \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf'''''''''_f'''''''''_Int_d ;
  logic \writeMerge_choice_CTf'''''''''_f'''''''''_Int_r ;
  \CTf'''''''''_f'''''''''_Int_t  \writeMerge_data_CTf'''''''''_f'''''''''_Int_d ;
  logic \writeMerge_data_CTf'''''''''_f'''''''''_Int_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_r ;
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \dconWriteIn_CTf'''''''''_f'''''''''_Int_d ;
  logic \dconWriteIn_CTf'''''''''_f'''''''''_Int_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \dconPtr_CTf'''''''''_f'''''''''_Int_d ;
  logic \dconPtr_CTf'''''''''_f'''''''''_Int_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  _169_d;
  logic _169_r;
  assign _169_r = 1'd1;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \demuxWriteResult_CTf'''''''''_f'''''''''_Int_d ;
  logic \demuxWriteResult_CTf'''''''''_f'''''''''_Int_r ;
  \Word16#_t  \initHP_CTf'_f'_Int_d ;
  logic \initHP_CTf'_f'_Int_r ;
  \Word16#_t  \incrHP_CTf'_f'_Int_d ;
  logic \incrHP_CTf'_f'_Int_r ;
  Go_t \incrHP_mergeCTf'_f'_Int_d ;
  logic \incrHP_mergeCTf'_f'_Int_r ;
  Go_t \incrHP_CTf'_f'_Int1_d ;
  logic \incrHP_CTf'_f'_Int1_r ;
  Go_t \incrHP_CTf'_f'_Int2_d ;
  logic \incrHP_CTf'_f'_Int2_r ;
  \Word16#_t  \addHP_CTf'_f'_Int_d ;
  logic \addHP_CTf'_f'_Int_r ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_d ;
  logic \mergeHP_CTf'_f'_Int_r ;
  Go_t \incrHP_mergeCTf'_f'_Int_buf_d ;
  logic \incrHP_mergeCTf'_f'_Int_buf_r ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_buf_d ;
  logic \mergeHP_CTf'_f'_Int_buf_r ;
  \Word16#_t  \forkHP1_CTf'_f'_Int_d ;
  logic \forkHP1_CTf'_f'_Int_r ;
  \Word16#_t  \forkHP1_CTf'_f'_In2_d ;
  logic \forkHP1_CTf'_f'_In2_r ;
  \Word16#_t  \forkHP1_CTf'_f'_In3_d ;
  logic \forkHP1_CTf'_f'_In3_r ;
  C2_t \memMergeChoice_CTf'_f'_Int_d ;
  logic \memMergeChoice_CTf'_f'_Int_r ;
  \MemIn_CTf'_f'_Int_t  \memMergeIn_CTf'_f'_Int_d ;
  logic \memMergeIn_CTf'_f'_Int_r ;
  \MemOut_CTf'_f'_Int_t  \memOut_CTf'_f'_Int_d ;
  logic \memOut_CTf'_f'_Int_r ;
  \MemOut_CTf'_f'_Int_t  \memReadOut_CTf'_f'_Int_d ;
  logic \memReadOut_CTf'_f'_Int_r ;
  \MemOut_CTf'_f'_Int_t  \memWriteOut_CTf'_f'_Int_d ;
  logic \memWriteOut_CTf'_f'_Int_r ;
  \MemIn_CTf'_f'_Int_t  \memMergeIn_CTf'_f'_Int_dbuf_d ;
  logic \memMergeIn_CTf'_f'_Int_dbuf_r ;
  \MemIn_CTf'_f'_Int_t  \memMergeIn_CTf'_f'_Int_rbuf_d ;
  logic \memMergeIn_CTf'_f'_Int_rbuf_r ;
  \MemOut_CTf'_f'_Int_t  \memOut_CTf'_f'_Int_dbuf_d ;
  logic \memOut_CTf'_f'_Int_dbuf_r ;
  \MemOut_CTf'_f'_Int_t  \memOut_CTf'_f'_Int_rbuf_d ;
  logic \memOut_CTf'_f'_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf'_f'_Int_d ;
  logic \destructReadIn_CTf'_f'_Int_r ;
  \MemIn_CTf'_f'_Int_t  \dconReadIn_CTf'_f'_Int_d ;
  logic \dconReadIn_CTf'_f'_Int_r ;
  \CTf'_f'_Int_t  \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf'_f'_Int_d ;
  logic \writeMerge_choice_CTf'_f'_Int_r ;
  \CTf'_f'_Int_t  \writeMerge_data_CTf'_f'_Int_d ;
  logic \writeMerge_data_CTf'_f'_Int_r ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_d ;
  logic \writeCTf'_f'_IntlizzieLet21_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_d ;
  logic \writeCTf'_f'_IntlizzieLet44_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_d ;
  logic \writeCTf'_f'_IntlizzieLet56_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_d ;
  logic \writeCTf'_f'_IntlizzieLet57_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_d ;
  logic \writeCTf'_f'_IntlizzieLet58_1_argbuf_r ;
  \MemIn_CTf'_f'_Int_t  \dconWriteIn_CTf'_f'_Int_d ;
  logic \dconWriteIn_CTf'_f'_Int_r ;
  \Pointer_CTf'_f'_Int_t  \dconPtr_CTf'_f'_Int_d ;
  logic \dconPtr_CTf'_f'_Int_r ;
  \Pointer_CTf'_f'_Int_t  _168_d;
  logic _168_r;
  assign _168_r = 1'd1;
  \Pointer_CTf'_f'_Int_t  \demuxWriteResult_CTf'_f'_Int_d ;
  logic \demuxWriteResult_CTf'_f'_Int_r ;
  \Word16#_t  initHP_CTf_f_Int_d;
  logic initHP_CTf_f_Int_r;
  \Word16#_t  incrHP_CTf_f_Int_d;
  logic incrHP_CTf_f_Int_r;
  Go_t incrHP_mergeCTf_f_Int_d;
  logic incrHP_mergeCTf_f_Int_r;
  Go_t incrHP_CTf_f_Int1_d;
  logic incrHP_CTf_f_Int1_r;
  Go_t incrHP_CTf_f_Int2_d;
  logic incrHP_CTf_f_Int2_r;
  \Word16#_t  addHP_CTf_f_Int_d;
  logic addHP_CTf_f_Int_r;
  \Word16#_t  mergeHP_CTf_f_Int_d;
  logic mergeHP_CTf_f_Int_r;
  Go_t incrHP_mergeCTf_f_Int_buf_d;
  logic incrHP_mergeCTf_f_Int_buf_r;
  \Word16#_t  mergeHP_CTf_f_Int_buf_d;
  logic mergeHP_CTf_f_Int_buf_r;
  \Word16#_t  forkHP1_CTf_f_Int_d;
  logic forkHP1_CTf_f_Int_r;
  \Word16#_t  forkHP1_CTf_f_In2_d;
  logic forkHP1_CTf_f_In2_r;
  \Word16#_t  forkHP1_CTf_f_In3_d;
  logic forkHP1_CTf_f_In3_r;
  C2_t memMergeChoice_CTf_f_Int_d;
  logic memMergeChoice_CTf_f_Int_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_d;
  logic memMergeIn_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_d;
  logic memOut_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memReadOut_CTf_f_Int_d;
  logic memReadOut_CTf_f_Int_r;
  MemOut_CTf_f_Int_t memWriteOut_CTf_f_Int_d;
  logic memWriteOut_CTf_f_Int_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_dbuf_d;
  logic memMergeIn_CTf_f_Int_dbuf_r;
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_rbuf_d;
  logic memMergeIn_CTf_f_Int_rbuf_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_dbuf_d;
  logic memOut_CTf_f_Int_dbuf_r;
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_rbuf_d;
  logic memOut_CTf_f_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTf_f_Int_d;
  logic destructReadIn_CTf_f_Int_r;
  MemIn_CTf_f_Int_t dconReadIn_CTf_f_Int_d;
  logic dconReadIn_CTf_f_Int_r;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_3_1_argbuf_d;
  logic readPointer_CTf_f_Intscfarg_0_3_1_argbuf_r;
  C5_t writeMerge_choice_CTf_f_Int_d;
  logic writeMerge_choice_CTf_f_Int_r;
  CTf_f_Int_t writeMerge_data_CTf_f_Int_d;
  logic writeMerge_data_CTf_f_Int_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet40_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet45_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet61_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet62_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_d;
  logic writeCTf_f_IntlizzieLet63_1_argbuf_r;
  MemIn_CTf_f_Int_t dconWriteIn_CTf_f_Int_d;
  logic dconWriteIn_CTf_f_Int_r;
  Pointer_CTf_f_Int_t dconPtr_CTf_f_Int_d;
  logic dconPtr_CTf_f_Int_r;
  Pointer_CTf_f_Int_t _167_d;
  logic _167_r;
  assign _167_r = 1'd1;
  Pointer_CTf_f_Int_t demuxWriteResult_CTf_f_Int_d;
  logic demuxWriteResult_CTf_f_Int_r;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  C2_t readMerge_choice_MaskQTree_d;
  logic readMerge_choice_MaskQTree_r;
  Pointer_MaskQTree_t readMerge_data_MaskQTree_d;
  logic readMerge_data_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreem1ae3_1_argbuf_d;
  logic readPointer_MaskQTreem1ae3_1_argbuf_r;
  MaskQTree_t readPointer_MaskQTreeq4aew_1_argbuf_d;
  logic readPointer_MaskQTreeq4aew_1_argbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t destructReadOut_MaskQTree_d;
  logic destructReadOut_MaskQTree_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _166_d;
  logic _166_r;
  assign _166_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_r ;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Int_t wsjQ_1_argbuf_d;
  logic wsjQ_1_argbuf_r;
  Int_t \es_6_1I#_d ;
  logic \es_6_1I#_r ;
  C2_t applyfnInt_Bool_5_choice_d;
  logic applyfnInt_Bool_5_choice_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5_data_d;
  logic applyfnInt_Bool_5_data_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t applyfnInt_Bool_5_2_argbuf_d;
  logic applyfnInt_Bool_5_2_argbuf_r;
  MyBool_t es_6_1_1_d;
  logic es_6_1_1_r;
  MyBool_t es_6_1_2_d;
  logic es_6_1_2_r;
  MyBool_t applyfnInt_Bool_5_1_d;
  logic applyfnInt_Bool_5_1_r;
  MyBool_t applyfnInt_Bool_5_2_d;
  logic applyfnInt_Bool_5_2_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyBool_t es_2_1_d;
  logic es_2_1_r;
  MyBool_t es_2_2_d;
  logic es_2_2_r;
  MyBool_t es_2_3_d;
  logic es_2_3_r;
  MyBool_t es_2_4_d;
  logic es_2_4_r;
  MyBool_t es_2_5_d;
  logic es_2_5_r;
  C3_t applyfnInt_Int_Int_5_choice_d;
  logic applyfnInt_Int_Int_5_choice_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5_data_d;
  logic applyfnInt_Int_Int_5_data_r;
  MyDTInt_Int_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Int_t applyfnInt_Int_Int_5_2_argbuf_d;
  logic applyfnInt_Int_Int_5_2_argbuf_r;
  QTree_Int_t es_3_1QVal_Int_d;
  logic es_3_1QVal_Int_r;
  Int_t applyfnInt_Int_Int_5_3_argbuf_d;
  logic applyfnInt_Int_Int_5_3_argbuf_r;
  Int_t es_5_1_1_argbuf_d;
  logic es_5_1_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_1_d;
  logic applyfnInt_Int_Int_5_1_r;
  Int_t applyfnInt_Int_Int_5_2_d;
  logic applyfnInt_Int_Int_5_2_r;
  Int_t applyfnInt_Int_Int_5_3_d;
  logic applyfnInt_Int_Int_5_3_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r;
  Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Int_t arg0_1Dcon_main1_d;
  logic arg0_1Dcon_main1_r;
  Int_t arg0_1Dcon_main1_1_d;
  logic arg0_1Dcon_main1_1_r;
  Int_t arg0_1Dcon_main1_2_d;
  logic arg0_1Dcon_main1_2_r;
  Int_t arg0_1Dcon_main1_3_d;
  logic arg0_1Dcon_main1_3_r;
  Int_t arg0_1Dcon_main1_4_d;
  logic arg0_1Dcon_main1_4_r;
  \Int#_t  xahT_destruct_d;
  logic xahT_destruct_r;
  Int_t \arg0_1Dcon_main1_1I#_d ;
  logic \arg0_1Dcon_main1_1I#_r ;
  Go_t \arg0_1Dcon_main1_3I#_d ;
  logic \arg0_1Dcon_main1_3I#_r ;
  Go_t \arg0_1Dcon_main1_3I#_1_d ;
  logic \arg0_1Dcon_main1_3I#_1_r ;
  Go_t \arg0_1Dcon_main1_3I#_2_d ;
  logic \arg0_1Dcon_main1_3I#_2_r ;
  Go_t \arg0_1Dcon_main1_3I#_3_d ;
  logic \arg0_1Dcon_main1_3I#_3_r ;
  Go_t \arg0_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_main1_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_main1_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1Xt_1_Eq_d;
  logic lizzieLet1_1wild1Xt_1_Eq_r;
  Go_t \arg0_1Dcon_main1_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_main1_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_main1_d;
  logic arg0_2Dcon_main1_r;
  Int_t \arg0_2_1Dcon_$fNumInt_$c+_d ;
  logic \arg0_2_1Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_4_r ;
  \Int#_t  xa1lV_destruct_d;
  logic xa1lV_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_1I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r ;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r ;
  \Int#_t  ya1lW_destruct_d;
  logic ya1lW_destruct_r;
  Int_t \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r ;
  \Int#_t  \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d ;
  logic \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r ;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  Int_t \es_0_1_1I#_mux_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r;
  Pointer_QTree_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r;
  Go_t call_$wnnz_Int_initBufi_d;
  logic call_$wnnz_Int_initBufi_r;
  C5_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t call_$wnnz_Int_unlockFork1_d;
  logic call_$wnnz_Int_unlockFork1_r;
  Go_t call_$wnnz_Int_unlockFork2_d;
  logic call_$wnnz_Int_unlockFork2_r;
  Go_t call_$wnnz_Int_unlockFork3_d;
  logic call_$wnnz_Int_unlockFork3_r;
  Go_t call_$wnnz_Int_initBuf_d;
  logic call_$wnnz_Int_initBuf_r;
  Go_t call_$wnnz_Int_goMux1_d;
  logic call_$wnnz_Int_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_Int_goMux2_d;
  logic call_$wnnz_Int_goMux2_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_Int_goMux3_d;
  logic call_$wnnz_Int_goMux3_r;
  Go_t \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d ;
  logic \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_r ;
  Pointer_MaskQTree_t \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d ;
  logic \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_r ;
  Pointer_QTree_Int_t \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d ;
  logic \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d ;
  logic \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_initBufi_d ;
  logic \call_f'''''''''_f'''''''''_Int_initBufi_r ;
  C5_t go_9_goMux_choice_d;
  logic go_9_goMux_choice_r;
  Go_t go_9_goMux_data_d;
  logic go_9_goMux_data_r;
  Go_t \call_f'''''''''_f'''''''''_Int_unlockFork1_d ;
  logic \call_f'''''''''_f'''''''''_Int_unlockFork1_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_unlockFork2_d ;
  logic \call_f'''''''''_f'''''''''_Int_unlockFork2_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_unlockFork3_d ;
  logic \call_f'''''''''_f'''''''''_Int_unlockFork3_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_unlockFork4_d ;
  logic \call_f'''''''''_f'''''''''_Int_unlockFork4_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_initBuf_d ;
  logic \call_f'''''''''_f'''''''''_Int_initBuf_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_goMux1_d ;
  logic \call_f'''''''''_f'''''''''_Int_goMux1_r ;
  Pointer_MaskQTree_t \call_f'''''''''_f'''''''''_Int_goMux2_d ;
  logic \call_f'''''''''_f'''''''''_Int_goMux2_r ;
  Pointer_QTree_Int_t \call_f'''''''''_f'''''''''_Int_goMux3_d ;
  logic \call_f'''''''''_f'''''''''_Int_goMux3_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \call_f'''''''''_f'''''''''_Int_goMux4_d ;
  logic \call_f'''''''''_f'''''''''_Int_goMux4_r ;
  Go_t \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_r ;
  Pointer_QTree_Int_t \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_r ;
  Pointer_QTree_Int_t \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_r ;
  MyDTInt_Bool_t \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_r ;
  MyDTInt_Int_Int_t \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_r ;
  \Pointer_CTf'_f'_Int_t  \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_r ;
  Go_t \call_f'_f'_Int_initBufi_d ;
  logic \call_f'_f'_Int_initBufi_r ;
  C5_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t \call_f'_f'_Int_unlockFork1_d ;
  logic \call_f'_f'_Int_unlockFork1_r ;
  Go_t \call_f'_f'_Int_unlockFork2_d ;
  logic \call_f'_f'_Int_unlockFork2_r ;
  Go_t \call_f'_f'_Int_unlockFork3_d ;
  logic \call_f'_f'_Int_unlockFork3_r ;
  Go_t \call_f'_f'_Int_unlockFork4_d ;
  logic \call_f'_f'_Int_unlockFork4_r ;
  Go_t \call_f'_f'_Int_unlockFork5_d ;
  logic \call_f'_f'_Int_unlockFork5_r ;
  Go_t \call_f'_f'_Int_unlockFork6_d ;
  logic \call_f'_f'_Int_unlockFork6_r ;
  Go_t \call_f'_f'_Int_initBuf_d ;
  logic \call_f'_f'_Int_initBuf_r ;
  Go_t \call_f'_f'_Int_goMux1_d ;
  logic \call_f'_f'_Int_goMux1_r ;
  Pointer_QTree_Int_t \call_f'_f'_Int_goMux2_d ;
  logic \call_f'_f'_Int_goMux2_r ;
  Pointer_QTree_Int_t \call_f'_f'_Int_goMux3_d ;
  logic \call_f'_f'_Int_goMux3_r ;
  MyDTInt_Bool_t \call_f'_f'_Int_goMux4_d ;
  logic \call_f'_f'_Int_goMux4_r ;
  MyDTInt_Int_Int_t \call_f'_f'_Int_goMux5_d ;
  logic \call_f'_f'_Int_goMux5_r ;
  \Pointer_CTf'_f'_Int_t  \call_f'_f'_Int_goMux6_d ;
  logic \call_f'_f'_Int_goMux6_r ;
  Go_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_r;
  Pointer_MaskQTree_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_r;
  Pointer_QTree_Int_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_r;
  Pointer_QTree_Int_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_r;
  MyDTInt_Bool_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_r;
  MyDTInt_Int_Int_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_r;
  Pointer_CTf_f_Int_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_r;
  Go_t call_f_f_Int_initBufi_d;
  logic call_f_f_Int_initBufi_r;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t call_f_f_Int_unlockFork1_d;
  logic call_f_f_Int_unlockFork1_r;
  Go_t call_f_f_Int_unlockFork2_d;
  logic call_f_f_Int_unlockFork2_r;
  Go_t call_f_f_Int_unlockFork3_d;
  logic call_f_f_Int_unlockFork3_r;
  Go_t call_f_f_Int_unlockFork4_d;
  logic call_f_f_Int_unlockFork4_r;
  Go_t call_f_f_Int_unlockFork5_d;
  logic call_f_f_Int_unlockFork5_r;
  Go_t call_f_f_Int_unlockFork6_d;
  logic call_f_f_Int_unlockFork6_r;
  Go_t call_f_f_Int_unlockFork7_d;
  logic call_f_f_Int_unlockFork7_r;
  Go_t call_f_f_Int_initBuf_d;
  logic call_f_f_Int_initBuf_r;
  Go_t call_f_f_Int_goMux1_d;
  logic call_f_f_Int_goMux1_r;
  Pointer_MaskQTree_t call_f_f_Int_goMux2_d;
  logic call_f_f_Int_goMux2_r;
  Pointer_QTree_Int_t call_f_f_Int_goMux3_d;
  logic call_f_f_Int_goMux3_r;
  Pointer_QTree_Int_t call_f_f_Int_goMux4_d;
  logic call_f_f_Int_goMux4_r;
  MyDTInt_Bool_t call_f_f_Int_goMux5_d;
  logic call_f_f_Int_goMux5_r;
  MyDTInt_Int_Int_t call_f_f_Int_goMux6_d;
  logic call_f_f_Int_goMux6_r;
  Pointer_CTf_f_Int_t call_f_f_Int_goMux7_d;
  logic call_f_f_Int_goMux7_r;
  QTree_Int_t lizzieLet30_1_1_argbuf_d;
  logic lizzieLet30_1_1_argbuf_r;
  Go_t es_2_1MyFalse_d;
  logic es_2_1MyFalse_r;
  Go_t es_2_1MyTrue_d;
  logic es_2_1MyTrue_r;
  Go_t es_2_1MyFalse_1_argbuf_d;
  logic es_2_1MyFalse_1_argbuf_r;
  Go_t es_2_1MyTrue_1_d;
  logic es_2_1MyTrue_1_r;
  Go_t es_2_1MyTrue_2_d;
  logic es_2_1MyTrue_2_r;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_d;
  logic es_2_1MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t es_2_1MyTrue_2_argbuf_d;
  logic es_2_1MyTrue_2_argbuf_r;
  MyDTInt_Int_Int_t es_2_2MyFalse_d;
  logic es_2_2MyFalse_r;
  MyDTInt_Int_Int_t _165_d;
  logic _165_r;
  assign _165_r = 1'd1;
  MyDTInt_Int_Int_t es_2_2MyFalse_1_argbuf_d;
  logic es_2_2MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r;
  \Pointer_CTf'_f'_Int_t  es_2_3MyFalse_d;
  logic es_2_3MyFalse_r;
  \Pointer_CTf'_f'_Int_t  es_2_3MyTrue_d;
  logic es_2_3MyTrue_r;
  \Pointer_CTf'_f'_Int_t  es_2_3MyFalse_1_argbuf_d;
  logic es_2_3MyFalse_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  es_2_3MyTrue_1_argbuf_d;
  logic es_2_3MyTrue_1_argbuf_r;
  Int_t es_2_4MyFalse_d;
  logic es_2_4MyFalse_r;
  Int_t _164_d;
  logic _164_r;
  assign _164_r = 1'd1;
  Int_t es_2_4MyFalse_1_argbuf_d;
  logic es_2_4MyFalse_1_argbuf_r;
  Int_t es_2_5MyFalse_d;
  logic es_2_5MyFalse_r;
  Int_t _163_d;
  logic _163_r;
  assign _163_r = 1'd1;
  Int_t es_2_5MyFalse_1_argbuf_d;
  logic es_2_5MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_CTf_f_Int_t es_6_1_1MyFalse_d;
  logic es_6_1_1MyFalse_r;
  Pointer_CTf_f_Int_t es_6_1_1MyTrue_d;
  logic es_6_1_1MyTrue_r;
  Pointer_CTf_f_Int_t es_6_1_1MyFalse_1_argbuf_d;
  logic es_6_1_1MyFalse_1_argbuf_r;
  Pointer_CTf_f_Int_t es_6_1_1MyTrue_1_argbuf_d;
  logic es_6_1_1MyTrue_1_argbuf_r;
  Go_t es_6_1_2MyFalse_d;
  logic es_6_1_2MyFalse_r;
  Go_t es_6_1_2MyTrue_d;
  logic es_6_1_2MyTrue_r;
  Go_t es_6_1_2MyFalse_1_d;
  logic es_6_1_2MyFalse_1_r;
  Go_t es_6_1_2MyFalse_2_d;
  logic es_6_1_2MyFalse_2_r;
  QTree_Int_t es_6_1_2MyFalse_1QError_Int_d;
  logic es_6_1_2MyFalse_1QError_Int_r;
  QTree_Int_t lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Go_t es_6_1_2MyFalse_2_argbuf_d;
  logic es_6_1_2MyFalse_2_argbuf_r;
  Go_t es_6_1_2MyTrue_1_d;
  logic es_6_1_2MyTrue_1_r;
  Go_t es_6_1_2MyTrue_2_d;
  logic es_6_1_2MyTrue_2_r;
  QTree_Int_t es_6_1_2MyTrue_1QNone_Int_d;
  logic es_6_1_2MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  Go_t es_6_1_2MyTrue_2_argbuf_d;
  logic es_6_1_2MyTrue_2_argbuf_r;
  \Int#_t  es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_d;
  logic es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_r;
  QTree_Int_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  C8_t \f'''''''''_f'''''''''_Int_choice_d ;
  logic \f'''''''''_f'''''''''_Int_choice_r ;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_data_d ;
  logic \f'''''''''_f'''''''''_Int_data_r ;
  Go_t go_12_1_d;
  logic go_12_1_r;
  Go_t go_12_2_d;
  logic go_12_2_r;
  Pointer_QTree_Int_t \q4'aex_1_1_argbuf_d ;
  logic \q4'aex_1_1_argbuf_r ;
  Pointer_MaskQTree_t q4aew_1_1_argbuf_d;
  logic q4aew_1_1_argbuf_r;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_resbuf_d ;
  logic \f'''''''''_f'''''''''_Int_resbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_2_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_2_argbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_3_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_3_argbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_4_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_4_argbuf_r ;
  QTree_Int_t es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_d;
  logic es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_r;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_5_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_5_argbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_6_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_6_argbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_7_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_7_argbuf_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_8_argbuf_d ;
  logic \f'''''''''_f'''''''''_Int_8_argbuf_r ;
  QTree_Int_t es_7_1es_8_1es_9_1es_10_1QNode_Int_d;
  logic es_7_1es_8_1es_9_1es_10_1QNode_Int_r;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_1_d ;
  logic \f'''''''''_f'''''''''_Int_1_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_2_d ;
  logic \f'''''''''_f'''''''''_Int_2_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_3_d ;
  logic \f'''''''''_f'''''''''_Int_3_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_4_d ;
  logic \f'''''''''_f'''''''''_Int_4_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_5_d ;
  logic \f'''''''''_f'''''''''_Int_5_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_6_d ;
  logic \f'''''''''_f'''''''''_Int_6_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_7_d ;
  logic \f'''''''''_f'''''''''_Int_7_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_8_d ;
  logic \f'''''''''_f'''''''''_Int_8_r ;
  Go_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_r ;
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_r ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_r ;
  Go_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_r ;
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_r ;
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_r ;
  MyDTInt_Bool_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_r ;
  MyDTInt_Int_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_r ;
  Go_t go_13_1_d;
  logic go_13_1_r;
  Go_t go_13_2_d;
  logic go_13_2_r;
  MyDTInt_Bool_t is_zaeJ_1_1_argbuf_d;
  logic is_zaeJ_1_1_argbuf_r;
  Pointer_QTree_Int_t m2aeH_1_1_argbuf_d;
  logic m2aeH_1_1_argbuf_r;
  Pointer_QTree_Int_t m3aeI_1_1_argbuf_d;
  logic m3aeI_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_addaeK_1_1_argbuf_d;
  logic op_addaeK_1_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Go_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r;
  Pointer_MaskQTree_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_r;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_r;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_r;
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_r;
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_r;
  Go_t go_14_1_d;
  logic go_14_1_r;
  Go_t go_14_2_d;
  logic go_14_2_r;
  MyDTInt_Bool_t is_zae6_1_1_argbuf_d;
  logic is_zae6_1_1_argbuf_r;
  Pointer_MaskQTree_t m1ae3_1_1_argbuf_d;
  logic m1ae3_1_1_argbuf_r;
  Pointer_QTree_Int_t m2ae4_1_1_argbuf_d;
  logic m2ae4_1_1_argbuf_r;
  Pointer_QTree_Int_t m3ae5_1_1_argbuf_d;
  logic m3ae5_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_addae7_1_1_argbuf_d;
  logic op_addae7_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_d ;
  logic \go_1Dcon_$fNumInt_$c+_r ;
  C5_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C5_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  C5_t go_10_goMux_choice_3_d;
  logic go_10_goMux_choice_3_r;
  C5_t go_10_goMux_choice_4_d;
  logic go_10_goMux_choice_4_r;
  C5_t go_10_goMux_choice_5_d;
  logic go_10_goMux_choice_5_r;
  Pointer_QTree_Int_t m2aeH_goMux_mux_d;
  logic m2aeH_goMux_mux_r;
  Pointer_QTree_Int_t m3aeI_goMux_mux_d;
  logic m3aeI_goMux_mux_r;
  MyDTInt_Bool_t is_zaeJ_goMux_mux_d;
  logic is_zaeJ_goMux_mux_r;
  MyDTInt_Int_Int_t op_addaeK_goMux_mux_d;
  logic op_addaeK_goMux_mux_r;
  \Pointer_CTf'_f'_Int_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  C5_t go_11_goMux_choice_3_d;
  logic go_11_goMux_choice_3_r;
  C5_t go_11_goMux_choice_4_d;
  logic go_11_goMux_choice_4_r;
  C5_t go_11_goMux_choice_5_d;
  logic go_11_goMux_choice_5_r;
  C5_t go_11_goMux_choice_6_d;
  logic go_11_goMux_choice_6_r;
  Pointer_MaskQTree_t m1ae3_goMux_mux_d;
  logic m1ae3_goMux_mux_r;
  Pointer_QTree_Int_t m2ae4_goMux_mux_d;
  logic m2ae4_goMux_mux_r;
  Pointer_QTree_Int_t m3ae5_goMux_mux_d;
  logic m3ae5_goMux_mux_r;
  MyDTInt_Bool_t is_zae6_goMux_mux_d;
  logic is_zae6_goMux_mux_r;
  MyDTInt_Int_Int_t op_addae7_goMux_mux_d;
  logic op_addae7_goMux_mux_r;
  Pointer_CTf_f_Int_t sc_0_3_goMux_mux_d;
  logic sc_0_3_goMux_mux_r;
  \CTf'''''''''_f'''''''''_Int_t  \go_12_1Lf'''''''''_f'''''''''_Intsbos_d ;
  logic \go_12_1Lf'''''''''_f'''''''''_Intsbos_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet43_1_argbuf_d;
  logic lizzieLet43_1_argbuf_r;
  Go_t go_12_2_argbuf_d;
  logic go_12_2_argbuf_r;
  \TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_t  \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d ;
  logic \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_r ;
  \CTf'_f'_Int_t  \go_13_1Lf'_f'_Intsbos_d ;
  logic \go_13_1Lf'_f'_Intsbos_r ;
  \CTf'_f'_Int_t  lizzieLet44_1_argbuf_d;
  logic lizzieLet44_1_argbuf_r;
  Go_t go_13_2_argbuf_d;
  logic go_13_2_argbuf_r;
  \TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_t  \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d ;
  logic \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_r ;
  CTf_f_Int_t go_14_1Lf_f_Intsbos_d;
  logic go_14_1Lf_f_Intsbos_r;
  CTf_f_Int_t lizzieLet45_1_argbuf_d;
  logic lizzieLet45_1_argbuf_r;
  Go_t go_14_2_argbuf_d;
  logic go_14_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_t call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d;
  logic call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r;
  C4_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C4_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C6_t go_16_goMux_choice_1_d;
  logic go_16_goMux_choice_1_r;
  C6_t go_16_goMux_choice_2_d;
  logic go_16_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C11_t go_17_goMux_choice_1_d;
  logic go_17_goMux_choice_1_r;
  C11_t go_17_goMux_choice_2_d;
  logic go_17_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTf'_f'_Int_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  C16_t go_18_goMux_choice_1_d;
  logic go_18_goMux_choice_1_r;
  C16_t go_18_goMux_choice_2_d;
  logic go_18_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_3_goMux_mux_d;
  logic srtarg_0_3_goMux_mux_r;
  Pointer_CTf_f_Int_t scfarg_0_3_goMux_mux_d;
  logic scfarg_0_3_goMux_mux_r;
  MyDTInt_Int_Int_t es_5_1_argbuf_d;
  logic es_5_1_argbuf_r;
  MyDTInt_Bool_t go_2Dcon_main1_d;
  logic go_2Dcon_main1_r;
  MyDTInt_Bool_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r;
  Go_t go_4_argbuf_d;
  logic go_4_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_d;
  logic go_6_1L$wnnz_Intsbos_r;
  CT$wnnz_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r;
  C5_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C5_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  Pointer_QTree_Int_t wsjQ_1_goMux_mux_d;
  logic wsjQ_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_9_goMux_choice_1_d;
  logic go_9_goMux_choice_1_r;
  C5_t go_9_goMux_choice_2_d;
  logic go_9_goMux_choice_2_r;
  C5_t go_9_goMux_choice_3_d;
  logic go_9_goMux_choice_3_r;
  Pointer_MaskQTree_t q4aew_goMux_mux_d;
  logic q4aew_goMux_mux_r;
  Pointer_QTree_Int_t \q4'aex_goMux_mux_d ;
  logic \q4'aex_goMux_mux_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  MyDTInt_Bool_t is_zae6_2_2_argbuf_d;
  logic is_zae6_2_2_argbuf_r;
  MyDTInt_Bool_t is_zae6_2_1_d;
  logic is_zae6_2_1_r;
  MyDTInt_Bool_t is_zae6_2_2_d;
  logic is_zae6_2_2_r;
  MyDTInt_Bool_t is_zae6_3_2_argbuf_d;
  logic is_zae6_3_2_argbuf_r;
  MyDTInt_Bool_t is_zae6_3_1_d;
  logic is_zae6_3_1_r;
  MyDTInt_Bool_t is_zae6_3_2_d;
  logic is_zae6_3_2_r;
  MyDTInt_Bool_t is_zae6_4_1_argbuf_d;
  logic is_zae6_4_1_argbuf_r;
  MyDTInt_Bool_t is_zaeJ_2_2_argbuf_d;
  logic is_zaeJ_2_2_argbuf_r;
  MyDTInt_Bool_t is_zaeJ_2_1_d;
  logic is_zaeJ_2_1_r;
  MyDTInt_Bool_t is_zaeJ_2_2_d;
  logic is_zaeJ_2_2_r;
  MyDTInt_Bool_t is_zaeJ_3_2_argbuf_d;
  logic is_zaeJ_3_2_argbuf_r;
  MyDTInt_Bool_t is_zaeJ_3_1_d;
  logic is_zaeJ_3_1_r;
  MyDTInt_Bool_t is_zaeJ_3_2_d;
  logic is_zaeJ_3_2_r;
  MyDTInt_Bool_t is_zaeJ_4_1_argbuf_d;
  logic is_zaeJ_4_1_argbuf_r;
  Pointer_QTree_Int_t q1aeR_destruct_d;
  logic q1aeR_destruct_r;
  Pointer_QTree_Int_t q2aeS_destruct_d;
  logic q2aeS_destruct_r;
  Pointer_QTree_Int_t q3aeT_destruct_d;
  logic q3aeT_destruct_r;
  Pointer_QTree_Int_t q4aeU_destruct_d;
  logic q4aeU_destruct_r;
  Int_t v1aeL_destruct_d;
  logic v1aeL_destruct_r;
  QTree_Int_t _162_d;
  logic _162_r;
  assign _162_r = 1'd1;
  QTree_Int_t lizzieLet13_1QVal_Int_d;
  logic lizzieLet13_1QVal_Int_r;
  QTree_Int_t lizzieLet13_1QNode_Int_d;
  logic lizzieLet13_1QNode_Int_r;
  QTree_Int_t _161_d;
  logic _161_r;
  assign _161_r = 1'd1;
  Go_t lizzieLet13_3QNone_Int_d;
  logic lizzieLet13_3QNone_Int_r;
  Go_t lizzieLet13_3QVal_Int_d;
  logic lizzieLet13_3QVal_Int_r;
  Go_t lizzieLet13_3QNode_Int_d;
  logic lizzieLet13_3QNode_Int_r;
  Go_t lizzieLet13_3QError_Int_d;
  logic lizzieLet13_3QError_Int_r;
  Go_t lizzieLet13_3QError_Int_1_d;
  logic lizzieLet13_3QError_Int_1_r;
  Go_t lizzieLet13_3QError_Int_2_d;
  logic lizzieLet13_3QError_Int_2_r;
  QTree_Int_t lizzieLet13_3QError_Int_1QError_Int_d;
  logic lizzieLet13_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t lizzieLet13_3QError_Int_2_argbuf_d;
  logic lizzieLet13_3QError_Int_2_argbuf_r;
  Go_t lizzieLet13_3QNone_Int_1_argbuf_d;
  logic lizzieLet13_3QNone_Int_1_argbuf_r;
  C11_t go_17_goMux_choice_d;
  logic go_17_goMux_choice_r;
  Go_t go_17_goMux_data_d;
  logic go_17_goMux_data_r;
  MyDTInt_Bool_t _160_d;
  logic _160_r;
  assign _160_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_4QVal_Int_d;
  logic lizzieLet13_4QVal_Int_r;
  MyDTInt_Bool_t lizzieLet13_4QNode_Int_d;
  logic lizzieLet13_4QNode_Int_r;
  MyDTInt_Bool_t _159_d;
  logic _159_r;
  assign _159_r = 1'd1;
  QTree_Int_t _158_d;
  logic _158_r;
  assign _158_r = 1'd1;
  QTree_Int_t lizzieLet13_5QVal_Int_d;
  logic lizzieLet13_5QVal_Int_r;
  QTree_Int_t lizzieLet13_5QNode_Int_d;
  logic lizzieLet13_5QNode_Int_r;
  QTree_Int_t _157_d;
  logic _157_r;
  assign _157_r = 1'd1;
  QTree_Int_t lizzieLet13_5QNode_Int_1_d;
  logic lizzieLet13_5QNode_Int_1_r;
  QTree_Int_t lizzieLet13_5QNode_Int_2_d;
  logic lizzieLet13_5QNode_Int_2_r;
  QTree_Int_t lizzieLet13_5QNode_Int_3_d;
  logic lizzieLet13_5QNode_Int_3_r;
  QTree_Int_t lizzieLet13_5QNode_Int_4_d;
  logic lizzieLet13_5QNode_Int_4_r;
  QTree_Int_t lizzieLet13_5QNode_Int_5_d;
  logic lizzieLet13_5QNode_Int_5_r;
  QTree_Int_t lizzieLet13_5QNode_Int_6_d;
  logic lizzieLet13_5QNode_Int_6_r;
  QTree_Int_t lizzieLet13_5QNode_Int_7_d;
  logic lizzieLet13_5QNode_Int_7_r;
  QTree_Int_t lizzieLet13_5QNode_Int_8_d;
  logic lizzieLet13_5QNode_Int_8_r;
  QTree_Int_t lizzieLet13_5QNode_Int_9_d;
  logic lizzieLet13_5QNode_Int_9_r;
  QTree_Int_t lizzieLet13_5QNode_Int_10_d;
  logic lizzieLet13_5QNode_Int_10_r;
  QTree_Int_t lizzieLet13_5QNode_Int_11_d;
  logic lizzieLet13_5QNode_Int_11_r;
  Pointer_QTree_Int_t _156_d;
  logic _156_r;
  assign _156_r = 1'd1;
  Pointer_QTree_Int_t _155_d;
  logic _155_r;
  assign _155_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_10QNode_Int_d;
  logic lizzieLet13_5QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _154_d;
  logic _154_r;
  assign _154_r = 1'd1;
  Pointer_QTree_Int_t _153_d;
  logic _153_r;
  assign _153_r = 1'd1;
  Pointer_QTree_Int_t _152_d;
  logic _152_r;
  assign _152_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_11QNode_Int_d;
  logic lizzieLet13_5QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _151_d;
  logic _151_r;
  assign _151_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1aeW_destruct_d;
  logic t1aeW_destruct_r;
  Pointer_QTree_Int_t t2aeX_destruct_d;
  logic t2aeX_destruct_r;
  Pointer_QTree_Int_t t3aeY_destruct_d;
  logic t3aeY_destruct_r;
  Pointer_QTree_Int_t t4aeZ_destruct_d;
  logic t4aeZ_destruct_r;
  QTree_Int_t _150_d;
  logic _150_r;
  assign _150_r = 1'd1;
  QTree_Int_t _149_d;
  logic _149_r;
  assign _149_r = 1'd1;
  QTree_Int_t lizzieLet13_5QNode_Int_1QNode_Int_d;
  logic lizzieLet13_5QNode_Int_1QNode_Int_r;
  QTree_Int_t _148_d;
  logic _148_r;
  assign _148_r = 1'd1;
  Go_t lizzieLet13_5QNode_Int_3QNone_Int_d;
  logic lizzieLet13_5QNode_Int_3QNone_Int_r;
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_r;
  Go_t lizzieLet13_5QNode_Int_3QNode_Int_d;
  logic lizzieLet13_5QNode_Int_3QNode_Int_r;
  Go_t lizzieLet13_5QNode_Int_3QError_Int_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_r;
  Go_t lizzieLet13_5QNode_Int_3QError_Int_1_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet13_5QNode_Int_3QError_Int_2_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_1_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_2_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_2_r;
  QTree_Int_t lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _147_d;
  logic _147_r;
  assign _147_r = 1'd1;
  MyDTInt_Bool_t _146_d;
  logic _146_r;
  assign _146_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_d;
  logic lizzieLet13_5QNode_Int_4QNode_Int_r;
  MyDTInt_Bool_t _145_d;
  logic _145_r;
  assign _145_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_1_d;
  logic lizzieLet13_5QNode_Int_4QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_2_d;
  logic lizzieLet13_5QNode_Int_4QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_d;
  logic lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_5QNone_Int_d;
  logic lizzieLet13_5QNode_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _144_d;
  logic _144_r;
  assign _144_r = 1'd1;
  Pointer_QTree_Int_t _143_d;
  logic _143_r;
  assign _143_r = 1'd1;
  Pointer_QTree_Int_t _142_d;
  logic _142_r;
  assign _142_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _141_d;
  logic _141_r;
  assign _141_r = 1'd1;
  MyDTInt_Int_Int_t _140_d;
  logic _140_r;
  assign _140_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_d;
  logic lizzieLet13_5QNode_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _139_d;
  logic _139_r;
  assign _139_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_1_d;
  logic lizzieLet13_5QNode_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_2_d;
  logic lizzieLet13_5QNode_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QNone_Int_d;
  logic lizzieLet13_5QNode_Int_7QNone_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QVal_Int_d;
  logic lizzieLet13_5QNode_Int_7QVal_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QNode_Int_d;
  logic lizzieLet13_5QNode_Int_7QNode_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QError_Int_d;
  logic lizzieLet13_5QNode_Int_7QError_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_r;
  \CTf'_f'_Int_t  \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_d ;
  logic \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_r ;
  \CTf'_f'_Int_t  lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _138_d;
  logic _138_r;
  assign _138_r = 1'd1;
  Pointer_QTree_Int_t _137_d;
  logic _137_r;
  assign _137_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_8QNode_Int_d;
  logic lizzieLet13_5QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _136_d;
  logic _136_r;
  assign _136_r = 1'd1;
  Pointer_QTree_Int_t _135_d;
  logic _135_r;
  assign _135_r = 1'd1;
  Pointer_QTree_Int_t _134_d;
  logic _134_r;
  assign _134_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_9QNode_Int_d;
  logic lizzieLet13_5QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _133_d;
  logic _133_r;
  assign _133_r = 1'd1;
  QTree_Int_t lizzieLet13_5QVal_Int_1_d;
  logic lizzieLet13_5QVal_Int_1_r;
  QTree_Int_t lizzieLet13_5QVal_Int_2_d;
  logic lizzieLet13_5QVal_Int_2_r;
  QTree_Int_t lizzieLet13_5QVal_Int_3_d;
  logic lizzieLet13_5QVal_Int_3_r;
  QTree_Int_t lizzieLet13_5QVal_Int_4_d;
  logic lizzieLet13_5QVal_Int_4_r;
  QTree_Int_t lizzieLet13_5QVal_Int_5_d;
  logic lizzieLet13_5QVal_Int_5_r;
  QTree_Int_t lizzieLet13_5QVal_Int_6_d;
  logic lizzieLet13_5QVal_Int_6_r;
  QTree_Int_t lizzieLet13_5QVal_Int_7_d;
  logic lizzieLet13_5QVal_Int_7_r;
  QTree_Int_t lizzieLet13_5QVal_Int_8_d;
  logic lizzieLet13_5QVal_Int_8_r;
  Int_t vaeM_destruct_d;
  logic vaeM_destruct_r;
  QTree_Int_t _132_d;
  logic _132_r;
  assign _132_r = 1'd1;
  QTree_Int_t lizzieLet13_5QVal_Int_1QVal_Int_d;
  logic lizzieLet13_5QVal_Int_1QVal_Int_r;
  QTree_Int_t _131_d;
  logic _131_r;
  assign _131_r = 1'd1;
  QTree_Int_t _130_d;
  logic _130_r;
  assign _130_r = 1'd1;
  Go_t lizzieLet13_5QVal_Int_3QNone_Int_d;
  logic lizzieLet13_5QVal_Int_3QNone_Int_r;
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_d;
  logic lizzieLet13_5QVal_Int_3QVal_Int_r;
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_r;
  Go_t lizzieLet13_5QVal_Int_3QError_Int_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_r;
  Go_t lizzieLet13_5QVal_Int_3QError_Int_1_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet13_5QVal_Int_3QError_Int_2_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_1_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_2_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_2_r;
  QTree_Int_t lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_1_d;
  logic lizzieLet13_5QVal_Int_3QVal_Int_1_r;
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_2_d;
  logic lizzieLet13_5QVal_Int_3QVal_Int_2_r;
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _129_d;
  logic _129_r;
  assign _129_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_5QVal_Int_4QVal_Int_d;
  logic lizzieLet13_5QVal_Int_4QVal_Int_r;
  MyDTInt_Bool_t _128_d;
  logic _128_r;
  assign _128_r = 1'd1;
  MyDTInt_Bool_t _127_d;
  logic _127_r;
  assign _127_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet13_5QVal_Int_5QNone_Int_d;
  logic lizzieLet13_5QVal_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _126_d;
  logic _126_r;
  assign _126_r = 1'd1;
  Pointer_QTree_Int_t _125_d;
  logic _125_r;
  assign _125_r = 1'd1;
  Pointer_QTree_Int_t _124_d;
  logic _124_r;
  assign _124_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _123_d;
  logic _123_r;
  assign _123_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_d;
  logic lizzieLet13_5QVal_Int_6QVal_Int_r;
  MyDTInt_Int_Int_t _122_d;
  logic _122_r;
  assign _122_r = 1'd1;
  MyDTInt_Int_Int_t _121_d;
  logic _121_r;
  assign _121_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_1_d;
  logic lizzieLet13_5QVal_Int_6QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_2_d;
  logic lizzieLet13_5QVal_Int_6QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNone_Int_d;
  logic lizzieLet13_5QVal_Int_7QNone_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QVal_Int_d;
  logic lizzieLet13_5QVal_Int_7QVal_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNode_Int_d;
  logic lizzieLet13_5QVal_Int_7QNode_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QError_Int_d;
  logic lizzieLet13_5QVal_Int_7QError_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_r;
  Int_t _120_d;
  logic _120_r;
  assign _120_r = 1'd1;
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_d;
  logic lizzieLet13_5QVal_Int_8QVal_Int_r;
  Int_t _119_d;
  logic _119_r;
  assign _119_r = 1'd1;
  Int_t _118_d;
  logic _118_r;
  assign _118_r = 1'd1;
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_1_d;
  logic lizzieLet13_5QVal_Int_8QVal_Int_1_r;
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_2_d;
  logic lizzieLet13_5QVal_Int_8QVal_Int_2_r;
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_d;
  logic lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _117_d;
  logic _117_r;
  assign _117_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_6QVal_Int_d;
  logic lizzieLet13_6QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet13_6QNode_Int_d;
  logic lizzieLet13_6QNode_Int_r;
  Pointer_QTree_Int_t _116_d;
  logic _116_r;
  assign _116_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_7QNone_Int_d;
  logic lizzieLet13_7QNone_Int_r;
  Pointer_QTree_Int_t _115_d;
  logic _115_r;
  assign _115_r = 1'd1;
  Pointer_QTree_Int_t _114_d;
  logic _114_r;
  assign _114_r = 1'd1;
  Pointer_QTree_Int_t _113_d;
  logic _113_r;
  assign _113_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_7QNone_Int_1_argbuf_d;
  logic lizzieLet13_7QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _112_d;
  logic _112_r;
  assign _112_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_8QVal_Int_d;
  logic lizzieLet13_8QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet13_8QNode_Int_d;
  logic lizzieLet13_8QNode_Int_r;
  MyDTInt_Int_Int_t _111_d;
  logic _111_r;
  assign _111_r = 1'd1;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QNone_Int_d;
  logic lizzieLet13_9QNone_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QVal_Int_d;
  logic lizzieLet13_9QVal_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QNode_Int_d;
  logic lizzieLet13_9QNode_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QError_Int_d;
  logic lizzieLet13_9QError_Int_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QError_Int_1_argbuf_d;
  logic lizzieLet13_9QError_Int_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QNone_Int_1_argbuf_d;
  logic lizzieLet13_9QNone_Int_1_argbuf_r;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_10MQNone_d;
  logic lizzieLet24_10MQNone_r;
  Pointer_CTf_f_Int_t lizzieLet24_10MQVal_d;
  logic lizzieLet24_10MQVal_r;
  Pointer_CTf_f_Int_t lizzieLet24_10MQNode_d;
  logic lizzieLet24_10MQNode_r;
  Pointer_CTf_f_Int_t lizzieLet24_10MQNone_1_argbuf_d;
  logic lizzieLet24_10MQNone_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_10MQVal_1_argbuf_d;
  logic lizzieLet24_10MQVal_1_argbuf_r;
  Pointer_MaskQTree_t q1ae8_destruct_d;
  logic q1ae8_destruct_r;
  Pointer_MaskQTree_t q2ae9_destruct_d;
  logic q2ae9_destruct_r;
  Pointer_MaskQTree_t q3aea_destruct_d;
  logic q3aea_destruct_r;
  Pointer_MaskQTree_t q4aeb_destruct_d;
  logic q4aeb_destruct_r;
  MaskQTree_t _110_d;
  logic _110_r;
  assign _110_r = 1'd1;
  MaskQTree_t _109_d;
  logic _109_r;
  assign _109_r = 1'd1;
  MaskQTree_t lizzieLet24_1MQNode_d;
  logic lizzieLet24_1MQNode_r;
  Go_t lizzieLet24_3MQNone_d;
  logic lizzieLet24_3MQNone_r;
  Go_t lizzieLet24_3MQVal_d;
  logic lizzieLet24_3MQVal_r;
  Go_t lizzieLet24_3MQNode_d;
  logic lizzieLet24_3MQNode_r;
  Go_t lizzieLet24_3MQNone_1_d;
  logic lizzieLet24_3MQNone_1_r;
  Go_t lizzieLet24_3MQNone_2_d;
  logic lizzieLet24_3MQNone_2_r;
  QTree_Int_t lizzieLet24_3MQNone_1QNone_Int_d;
  logic lizzieLet24_3MQNone_1QNone_Int_r;
  QTree_Int_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Go_t lizzieLet24_3MQNone_2_argbuf_d;
  logic lizzieLet24_3MQNone_2_argbuf_r;
  C16_t go_18_goMux_choice_d;
  logic go_18_goMux_choice_r;
  Go_t go_18_goMux_data_d;
  logic go_18_goMux_data_r;
  Go_t lizzieLet24_3MQVal_1_d;
  logic lizzieLet24_3MQVal_1_r;
  Go_t lizzieLet24_3MQVal_2_d;
  logic lizzieLet24_3MQVal_2_r;
  Go_t lizzieLet24_3MQVal_1_argbuf_d;
  logic lizzieLet24_3MQVal_1_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r ;
  Go_t lizzieLet24_3MQVal_2_argbuf_d;
  logic lizzieLet24_3MQVal_2_argbuf_r;
  MyDTInt_Bool_t _108_d;
  logic _108_r;
  assign _108_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_4MQVal_d;
  logic lizzieLet24_4MQVal_r;
  MyDTInt_Bool_t lizzieLet24_4MQNode_d;
  logic lizzieLet24_4MQNode_r;
  MyDTInt_Bool_t lizzieLet24_4MQVal_1_argbuf_d;
  logic lizzieLet24_4MQVal_1_argbuf_r;
  QTree_Int_t _107_d;
  logic _107_r;
  assign _107_r = 1'd1;
  QTree_Int_t _106_d;
  logic _106_r;
  assign _106_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_d;
  logic lizzieLet24_5MQNode_r;
  QTree_Int_t lizzieLet24_5MQNode_1_d;
  logic lizzieLet24_5MQNode_1_r;
  QTree_Int_t lizzieLet24_5MQNode_2_d;
  logic lizzieLet24_5MQNode_2_r;
  QTree_Int_t lizzieLet24_5MQNode_3_d;
  logic lizzieLet24_5MQNode_3_r;
  QTree_Int_t lizzieLet24_5MQNode_4_d;
  logic lizzieLet24_5MQNode_4_r;
  QTree_Int_t lizzieLet24_5MQNode_5_d;
  logic lizzieLet24_5MQNode_5_r;
  QTree_Int_t lizzieLet24_5MQNode_6_d;
  logic lizzieLet24_5MQNode_6_r;
  QTree_Int_t lizzieLet24_5MQNode_7_d;
  logic lizzieLet24_5MQNode_7_r;
  QTree_Int_t lizzieLet24_5MQNode_8_d;
  logic lizzieLet24_5MQNode_8_r;
  QTree_Int_t lizzieLet24_5MQNode_9_d;
  logic lizzieLet24_5MQNode_9_r;
  QTree_Int_t lizzieLet24_5MQNode_10_d;
  logic lizzieLet24_5MQNode_10_r;
  QTree_Int_t lizzieLet24_5MQNode_11_d;
  logic lizzieLet24_5MQNode_11_r;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_10QNone_Int_d;
  logic lizzieLet24_5MQNode_10QNone_Int_r;
  Pointer_MaskQTree_t _105_d;
  logic _105_r;
  assign _105_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_10QNode_Int_d;
  logic lizzieLet24_5MQNode_10QNode_Int_r;
  Pointer_MaskQTree_t _104_d;
  logic _104_r;
  assign _104_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_11QNone_Int_d;
  logic lizzieLet24_5MQNode_11QNone_Int_r;
  Pointer_MaskQTree_t _103_d;
  logic _103_r;
  assign _103_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_11QNode_Int_d;
  logic lizzieLet24_5MQNode_11QNode_Int_r;
  Pointer_MaskQTree_t _102_d;
  logic _102_r;
  assign _102_r = 1'd1;
  Pointer_QTree_Int_t \q1'aen_destruct_d ;
  logic \q1'aen_destruct_r ;
  Pointer_QTree_Int_t \q2'aeo_destruct_d ;
  logic \q2'aeo_destruct_r ;
  Pointer_QTree_Int_t \q3'aep_destruct_d ;
  logic \q3'aep_destruct_r ;
  Pointer_QTree_Int_t \q4'aeq_destruct_d ;
  logic \q4'aeq_destruct_r ;
  Int_t v1aeh_destruct_d;
  logic v1aeh_destruct_r;
  QTree_Int_t _101_d;
  logic _101_r;
  assign _101_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_1QVal_Int_d;
  logic lizzieLet24_5MQNode_1QVal_Int_r;
  QTree_Int_t lizzieLet24_5MQNode_1QNode_Int_d;
  logic lizzieLet24_5MQNode_1QNode_Int_r;
  QTree_Int_t _100_d;
  logic _100_r;
  assign _100_r = 1'd1;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QNone_Int_d;
  logic lizzieLet24_5MQNode_3QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QVal_Int_d;
  logic lizzieLet24_5MQNode_3QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QNode_Int_d;
  logic lizzieLet24_5MQNode_3QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QError_Int_d;
  logic lizzieLet24_5MQNode_3QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QError_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_3QError_Int_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_4QNone_Int_d;
  logic lizzieLet24_5MQNode_4QNone_Int_r;
  Go_t lizzieLet24_5MQNode_4QVal_Int_d;
  logic lizzieLet24_5MQNode_4QVal_Int_r;
  Go_t lizzieLet24_5MQNode_4QNode_Int_d;
  logic lizzieLet24_5MQNode_4QNode_Int_r;
  Go_t lizzieLet24_5MQNode_4QError_Int_d;
  logic lizzieLet24_5MQNode_4QError_Int_r;
  Go_t lizzieLet24_5MQNode_4QError_Int_1_d;
  logic lizzieLet24_5MQNode_4QError_Int_1_r;
  Go_t lizzieLet24_5MQNode_4QError_Int_2_d;
  logic lizzieLet24_5MQNode_4QError_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_4QError_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet42_1_argbuf_d;
  logic lizzieLet42_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_4QError_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_4QError_Int_2_argbuf_r;
  MyDTInt_Bool_t _99_d;
  logic _99_r;
  assign _99_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_5MQNode_5QVal_Int_d;
  logic lizzieLet24_5MQNode_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet24_5MQNode_5QNode_Int_d;
  logic lizzieLet24_5MQNode_5QNode_Int_r;
  MyDTInt_Bool_t _98_d;
  logic _98_r;
  assign _98_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_r;
  QTree_Int_t _97_d;
  logic _97_r;
  assign _97_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_1_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_3_d;
  logic lizzieLet24_5MQNode_6QNode_Int_3_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_4_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_5_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_7_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_8_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_9_d;
  logic lizzieLet24_5MQNode_6QNode_Int_9_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_10_d;
  logic lizzieLet24_5MQNode_6QNode_Int_10_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11_d;
  logic lizzieLet24_5MQNode_6QNode_Int_11_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12_d;
  logic lizzieLet24_5MQNode_6QNode_Int_12_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13_d;
  logic lizzieLet24_5MQNode_6QNode_Int_13_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14_r;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_r;
  Pointer_MaskQTree_t _96_d;
  logic _96_r;
  assign _96_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_r;
  Pointer_MaskQTree_t _95_d;
  logic _95_r;
  assign _95_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_r;
  Pointer_QTree_Int_t _94_d;
  logic _94_r;
  assign _94_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_r;
  Pointer_QTree_Int_t _93_d;
  logic _93_r;
  assign _93_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_r;
  Pointer_QTree_Int_t _92_d;
  logic _92_r;
  assign _92_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_r;
  Pointer_QTree_Int_t _91_d;
  logic _91_r;
  assign _91_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_r;
  Pointer_QTree_Int_t _90_d;
  logic _90_r;
  assign _90_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_r;
  Pointer_QTree_Int_t _89_d;
  logic _89_r;
  assign _89_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_r;
  Pointer_QTree_Int_t _88_d;
  logic _88_r;
  assign _88_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_r;
  Pointer_QTree_Int_t _87_d;
  logic _87_r;
  assign _87_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1aes_destruct_d;
  logic t1aes_destruct_r;
  Pointer_QTree_Int_t t2aet_destruct_d;
  logic t2aet_destruct_r;
  Pointer_QTree_Int_t t3aeu_destruct_d;
  logic t3aeu_destruct_r;
  Pointer_QTree_Int_t t4aev_destruct_d;
  logic t4aev_destruct_r;
  QTree_Int_t _86_d;
  logic _86_r;
  assign _86_r = 1'd1;
  QTree_Int_t _85_d;
  logic _85_r;
  assign _85_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_r;
  QTree_Int_t _84_d;
  logic _84_r;
  assign _84_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_r;
  Pointer_MaskQTree_t _83_d;
  logic _83_r;
  assign _83_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_r;
  Pointer_MaskQTree_t _82_d;
  logic _82_r;
  assign _82_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_r;
  Pointer_MaskQTree_t _81_d;
  logic _81_r;
  assign _81_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_r;
  Pointer_MaskQTree_t _80_d;
  logic _80_r;
  assign _80_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_r;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QError_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_r;
  CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_r;
  CTf_f_Int_t lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet41_1_argbuf_d;
  logic lizzieLet41_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_r ;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_r ;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_r ;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_r ;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _79_d;
  logic _79_r;
  assign _79_r = 1'd1;
  MyDTInt_Bool_t _78_d;
  logic _78_r;
  assign _78_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_r;
  MyDTInt_Bool_t _77_d;
  logic _77_r;
  assign _77_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t _76_d;
  logic _76_r;
  assign _76_r = 1'd1;
  MyDTInt_Int_Int_t _75_d;
  logic _75_r;
  assign _75_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_r;
  MyDTInt_Int_Int_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_r;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_r;
  Pointer_MaskQTree_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_r;
  Pointer_MaskQTree_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_1_d;
  logic lizzieLet24_5MQNode_6QNone_Int_1_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_2_d;
  logic lizzieLet24_5MQNode_6QNone_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_3_d;
  logic lizzieLet24_5MQNode_6QNone_Int_3_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_4_d;
  logic lizzieLet24_5MQNode_6QNone_Int_4_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_5_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_7_d;
  logic lizzieLet24_5MQNode_6QNone_Int_7_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_8_d;
  logic lizzieLet24_5MQNode_6QNone_Int_8_r;
  Pointer_QTree_Int_t t1aed_destruct_d;
  logic t1aed_destruct_r;
  Pointer_QTree_Int_t t2aee_destruct_d;
  logic t2aee_destruct_r;
  Pointer_QTree_Int_t t3aef_destruct_d;
  logic t3aef_destruct_r;
  Pointer_QTree_Int_t t4aeg_destruct_d;
  logic t4aeg_destruct_r;
  QTree_Int_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  QTree_Int_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_r;
  QTree_Int_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  Pointer_MaskQTree_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  Pointer_MaskQTree_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_r;
  Pointer_MaskQTree_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_r;
  Pointer_MaskQTree_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  Pointer_MaskQTree_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_r;
  Pointer_MaskQTree_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QError_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_r ;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_r ;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_r ;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_r;
  TupGo___Pointer_MaskQTree___Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_r ;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet28_2_1_argbuf_d;
  logic lizzieLet28_2_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet29_1_1_argbuf_d;
  logic lizzieLet29_1_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_r;
  Pointer_MaskQTree_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Pointer_MaskQTree_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_r;
  Pointer_MaskQTree_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_r;
  Pointer_MaskQTree_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  Pointer_MaskQTree_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_d;
  logic lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_r;
  Pointer_MaskQTree_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_1_d;
  logic lizzieLet24_5MQNode_6QVal_Int_1_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_2_d;
  logic lizzieLet24_5MQNode_6QVal_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_3_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_5_d;
  logic lizzieLet24_5MQNode_6QVal_Int_5_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_6_d;
  logic lizzieLet24_5MQNode_6QVal_Int_6_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_7_d;
  logic lizzieLet24_5MQNode_6QVal_Int_7_r;
  Int_t vaei_destruct_d;
  logic vaei_destruct_r;
  QTree_Int_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_r;
  QTree_Int_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  QTree_Int_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QError_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QError_Int_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_r;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet33_1_1_argbuf_d;
  logic lizzieLet33_1_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_r;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_r;
  QTree_Int_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_r;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r;
  MyDTInt_Bool_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_r;
  MyDTInt_Bool_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  MyDTInt_Bool_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_r;
  MyDTInt_Int_Int_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  MyDTInt_Int_Int_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r;
  Int_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  Int_t lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_d;
  logic lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_r;
  Int_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  Int_t lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_7QVal_Int_d;
  logic lizzieLet24_5MQNode_7QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_7QNode_Int_d;
  logic lizzieLet24_5MQNode_7QNode_Int_r;
  MyDTInt_Int_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_8QNone_Int_d;
  logic lizzieLet24_5MQNode_8QNone_Int_r;
  Pointer_MaskQTree_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_8QNode_Int_d;
  logic lizzieLet24_5MQNode_8QNode_Int_r;
  Pointer_MaskQTree_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_9QNone_Int_d;
  logic lizzieLet24_5MQNode_9QNone_Int_r;
  Pointer_MaskQTree_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_9QNode_Int_d;
  logic lizzieLet24_5MQNode_9QNode_Int_r;
  Pointer_MaskQTree_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  QTree_Int_t lizzieLet24_6MQNode_d;
  logic lizzieLet24_6MQNode_r;
  Pointer_QTree_Int_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_7MQVal_d;
  logic lizzieLet24_7MQVal_r;
  Pointer_QTree_Int_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_7MQVal_1_argbuf_d;
  logic lizzieLet24_7MQVal_1_argbuf_r;
  Pointer_QTree_Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_8MQVal_d;
  logic lizzieLet24_8MQVal_r;
  Pointer_QTree_Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet24_8MQVal_1_argbuf_d;
  logic lizzieLet24_8MQVal_1_argbuf_r;
  MyDTInt_Int_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet24_9MQVal_d;
  logic lizzieLet24_9MQVal_r;
  MyDTInt_Int_Int_t lizzieLet24_9MQNode_d;
  logic lizzieLet24_9MQNode_r;
  MyDTInt_Int_Int_t lizzieLet24_9MQVal_1_argbuf_d;
  logic lizzieLet24_9MQVal_1_argbuf_r;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  \Int#_t  wwsjT_4_destruct_d;
  logic wwsjT_4_destruct_r;
  \Int#_t  ww1Xkr_2_destruct_d;
  logic ww1Xkr_2_destruct_r;
  \Int#_t  ww2Xku_1_destruct_d;
  logic ww2Xku_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  \Int#_t  wwsjT_3_destruct_d;
  logic wwsjT_3_destruct_r;
  \Int#_t  ww1Xkr_1_destruct_d;
  logic ww1Xkr_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Int_t q4a88_3_destruct_d;
  logic q4a88_3_destruct_r;
  \Int#_t  wwsjT_2_destruct_d;
  logic wwsjT_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4a88_2_destruct_d;
  logic q4a88_2_destruct_r;
  Pointer_QTree_Int_t q3a87_2_destruct_d;
  logic q3a87_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4a88_1_destruct_d;
  logic q4a88_1_destruct_r;
  Pointer_QTree_Int_t q3a87_1_destruct_d;
  logic q3a87_1_destruct_r;
  Pointer_QTree_Int_t q2a86_1_destruct_d;
  logic q2a86_1_destruct_r;
  CT$wnnz_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  CT$wnnz_Int_t lizzieLet46_1Lcall_$wnnz_Int3_d;
  logic lizzieLet46_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet46_1Lcall_$wnnz_Int2_d;
  logic lizzieLet46_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet46_1Lcall_$wnnz_Int1_d;
  logic lizzieLet46_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet46_1Lcall_$wnnz_Int0_d;
  logic lizzieLet46_1Lcall_$wnnz_Int0_r;
  Go_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  Go_t lizzieLet46_3Lcall_$wnnz_Int3_d;
  logic lizzieLet46_3Lcall_$wnnz_Int3_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int2_d;
  logic lizzieLet46_3Lcall_$wnnz_Int2_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int1_d;
  logic lizzieLet46_3Lcall_$wnnz_Int1_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int0_d;
  logic lizzieLet46_3Lcall_$wnnz_Int0_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_d;
  logic lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_d;
  logic lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_d;
  logic lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_r;
  Go_t lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_d;
  logic lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_r;
  \Int#_t  lizzieLet46_4L$wnnz_Intsbos_d;
  logic lizzieLet46_4L$wnnz_Intsbos_r;
  \Int#_t  lizzieLet46_4Lcall_$wnnz_Int3_d;
  logic lizzieLet46_4Lcall_$wnnz_Int3_r;
  \Int#_t  lizzieLet46_4Lcall_$wnnz_Int2_d;
  logic lizzieLet46_4Lcall_$wnnz_Int2_r;
  \Int#_t  lizzieLet46_4Lcall_$wnnz_Int1_d;
  logic lizzieLet46_4Lcall_$wnnz_Int1_r;
  \Int#_t  lizzieLet46_4Lcall_$wnnz_Int0_d;
  logic lizzieLet46_4Lcall_$wnnz_Int0_r;
  \Int#_t  lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_Int_goConst_d;
  logic call_$wnnz_Int_goConst_r;
  \Int#_t  \$wnnz_Int_resbuf_d ;
  logic \$wnnz_Int_resbuf_r ;
  CT$wnnz_Int_t lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_d;
  logic lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet47_1_argbuf_d;
  logic lizzieLet47_1_argbuf_r;
  Pointer_QTree_Int_t q1a85_destruct_d;
  logic q1a85_destruct_r;
  Pointer_QTree_Int_t q2a86_destruct_d;
  logic q2a86_destruct_r;
  Pointer_QTree_Int_t q3a87_destruct_d;
  logic q3a87_destruct_r;
  Pointer_QTree_Int_t q4a88_destruct_d;
  logic q4a88_destruct_r;
  QTree_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  QTree_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet28_1_1_argbuf_d;
  logic lizzieLet28_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_d;
  logic lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t es_1_2_destruct_d;
  logic es_1_2_destruct_r;
  Pointer_QTree_Int_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Int_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Int_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_MaskQTree_t q1aey_3_destruct_d;
  logic q1aey_3_destruct_r;
  Pointer_QTree_Int_t t1aeD_3_destruct_d;
  logic t1aeD_3_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_MaskQTree_t q1aey_2_destruct_d;
  logic q1aey_2_destruct_r;
  Pointer_QTree_Int_t t1aeD_2_destruct_d;
  logic t1aeD_2_destruct_r;
  Pointer_MaskQTree_t q2aez_2_destruct_d;
  logic q2aez_2_destruct_r;
  Pointer_QTree_Int_t t2aeE_2_destruct_d;
  logic t2aeE_2_destruct_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_MaskQTree_t q1aey_1_destruct_d;
  logic q1aey_1_destruct_r;
  Pointer_QTree_Int_t t1aeD_1_destruct_d;
  logic t1aeD_1_destruct_r;
  Pointer_MaskQTree_t q2aez_1_destruct_d;
  logic q2aez_1_destruct_r;
  Pointer_QTree_Int_t t2aeE_1_destruct_d;
  logic t2aeE_1_destruct_r;
  Pointer_MaskQTree_t q3aeA_1_destruct_d;
  logic q3aeA_1_destruct_r;
  Pointer_QTree_Int_t t3aeF_1_destruct_d;
  logic t3aeF_1_destruct_r;
  \CTf'''''''''_f'''''''''_Int_t  _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d ;
  logic \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_r ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d ;
  logic \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_r ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d ;
  logic \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_r ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d ;
  logic \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_r ;
  Go_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_r ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d ;
  logic \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_r ;
  QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_r ;
  QTree_Int_t lizzieLet54_1_argbuf_d;
  logic lizzieLet54_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet53_1_argbuf_d;
  logic lizzieLet53_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet52_1_argbuf_d;
  logic lizzieLet52_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet51_1_argbuf_d;
  logic lizzieLet51_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f'''''''''_f'''''''''_Int_goConst_d ;
  logic \call_f'''''''''_f'''''''''_Int_goConst_r ;
  Pointer_QTree_Int_t es_5_2_destruct_d;
  logic es_5_2_destruct_r;
  Pointer_QTree_Int_t es_6_4_destruct_d;
  logic es_6_4_destruct_r;
  Pointer_QTree_Int_t es_7_3_destruct_d;
  logic es_7_3_destruct_r;
  \Pointer_CTf'_f'_Int_t  sc_0_15_destruct_d;
  logic sc_0_15_destruct_r;
  Pointer_QTree_Int_t es_6_3_destruct_d;
  logic es_6_3_destruct_r;
  Pointer_QTree_Int_t es_7_2_destruct_d;
  logic es_7_2_destruct_r;
  \Pointer_CTf'_f'_Int_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t q1aeR_3_destruct_d;
  logic q1aeR_3_destruct_r;
  Pointer_QTree_Int_t t1aeW_3_destruct_d;
  logic t1aeW_3_destruct_r;
  MyDTInt_Bool_t is_zaeJ_4_destruct_d;
  logic is_zaeJ_4_destruct_r;
  MyDTInt_Int_Int_t op_addaeK_4_destruct_d;
  logic op_addaeK_4_destruct_r;
  Pointer_QTree_Int_t es_7_1_destruct_d;
  logic es_7_1_destruct_r;
  \Pointer_CTf'_f'_Int_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t q1aeR_2_destruct_d;
  logic q1aeR_2_destruct_r;
  Pointer_QTree_Int_t t1aeW_2_destruct_d;
  logic t1aeW_2_destruct_r;
  MyDTInt_Bool_t is_zaeJ_3_destruct_d;
  logic is_zaeJ_3_destruct_r;
  MyDTInt_Int_Int_t op_addaeK_3_destruct_d;
  logic op_addaeK_3_destruct_r;
  Pointer_QTree_Int_t q2aeS_2_destruct_d;
  logic q2aeS_2_destruct_r;
  Pointer_QTree_Int_t t2aeX_2_destruct_d;
  logic t2aeX_2_destruct_r;
  \Pointer_CTf'_f'_Int_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t q1aeR_1_destruct_d;
  logic q1aeR_1_destruct_r;
  Pointer_QTree_Int_t t1aeW_1_destruct_d;
  logic t1aeW_1_destruct_r;
  MyDTInt_Bool_t is_zaeJ_2_destruct_d;
  logic is_zaeJ_2_destruct_r;
  MyDTInt_Int_Int_t op_addaeK_2_destruct_d;
  logic op_addaeK_2_destruct_r;
  Pointer_QTree_Int_t q2aeS_1_destruct_d;
  logic q2aeS_1_destruct_r;
  Pointer_QTree_Int_t t2aeX_1_destruct_d;
  logic t2aeX_1_destruct_r;
  Pointer_QTree_Int_t q3aeT_1_destruct_d;
  logic q3aeT_1_destruct_r;
  Pointer_QTree_Int_t t3aeY_1_destruct_d;
  logic t3aeY_1_destruct_r;
  \CTf'_f'_Int_t  _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  \CTf'_f'_Int_t  \lizzieLet55_1Lcall_f'_f'_Int3_d ;
  logic \lizzieLet55_1Lcall_f'_f'_Int3_r ;
  \CTf'_f'_Int_t  \lizzieLet55_1Lcall_f'_f'_Int2_d ;
  logic \lizzieLet55_1Lcall_f'_f'_Int2_r ;
  \CTf'_f'_Int_t  \lizzieLet55_1Lcall_f'_f'_Int1_d ;
  logic \lizzieLet55_1Lcall_f'_f'_Int1_r ;
  \CTf'_f'_Int_t  \lizzieLet55_1Lcall_f'_f'_Int0_d ;
  logic \lizzieLet55_1Lcall_f'_f'_Int0_r ;
  Go_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int3_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int3_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int2_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int2_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int1_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int1_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int0_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int0_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_r ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lf'_f'_Intsbos_d ;
  logic \lizzieLet55_4Lf'_f'_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int3_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int2_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int1_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int0_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int0_r ;
  QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r ;
  QTree_Int_t lizzieLet59_1_argbuf_d;
  logic lizzieLet59_1_argbuf_r;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_r ;
  \CTf'_f'_Int_t  lizzieLet58_1_argbuf_d;
  logic lizzieLet58_1_argbuf_r;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_r ;
  \CTf'_f'_Int_t  lizzieLet57_1_argbuf_d;
  logic lizzieLet57_1_argbuf_r;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_r ;
  \CTf'_f'_Int_t  lizzieLet56_1_argbuf_d;
  logic lizzieLet56_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f'_f'_Int_goConst_d ;
  logic \call_f'_f'_Int_goConst_r ;
  Pointer_QTree_Int_t \f'_f'_Int_resbuf_d ;
  logic \f'_f'_Int_resbuf_r ;
  Pointer_QTree_Int_t es_12_destruct_d;
  logic es_12_destruct_r;
  Pointer_QTree_Int_t es_13_1_destruct_d;
  logic es_13_1_destruct_r;
  Pointer_QTree_Int_t es_14_2_destruct_d;
  logic es_14_2_destruct_r;
  Pointer_CTf_f_Int_t sc_0_19_destruct_d;
  logic sc_0_19_destruct_r;
  Pointer_QTree_Int_t es_13_destruct_d;
  logic es_13_destruct_r;
  Pointer_QTree_Int_t es_14_1_destruct_d;
  logic es_14_1_destruct_r;
  Pointer_CTf_f_Int_t sc_0_18_destruct_d;
  logic sc_0_18_destruct_r;
  Pointer_MaskQTree_t q1ae8_3_destruct_d;
  logic q1ae8_3_destruct_r;
  Pointer_QTree_Int_t \q1'aen_3_destruct_d ;
  logic \q1'aen_3_destruct_r ;
  Pointer_QTree_Int_t t1aes_3_destruct_d;
  logic t1aes_3_destruct_r;
  MyDTInt_Bool_t is_zae6_4_destruct_d;
  logic is_zae6_4_destruct_r;
  MyDTInt_Int_Int_t op_addae7_4_destruct_d;
  logic op_addae7_4_destruct_r;
  Pointer_QTree_Int_t es_14_destruct_d;
  logic es_14_destruct_r;
  Pointer_CTf_f_Int_t sc_0_17_destruct_d;
  logic sc_0_17_destruct_r;
  Pointer_MaskQTree_t q1ae8_2_destruct_d;
  logic q1ae8_2_destruct_r;
  Pointer_QTree_Int_t \q1'aen_2_destruct_d ;
  logic \q1'aen_2_destruct_r ;
  Pointer_QTree_Int_t t1aes_2_destruct_d;
  logic t1aes_2_destruct_r;
  MyDTInt_Bool_t is_zae6_3_destruct_d;
  logic is_zae6_3_destruct_r;
  MyDTInt_Int_Int_t op_addae7_3_destruct_d;
  logic op_addae7_3_destruct_r;
  Pointer_MaskQTree_t q2ae9_2_destruct_d;
  logic q2ae9_2_destruct_r;
  Pointer_QTree_Int_t \q2'aeo_2_destruct_d ;
  logic \q2'aeo_2_destruct_r ;
  Pointer_QTree_Int_t t2aet_2_destruct_d;
  logic t2aet_2_destruct_r;
  Pointer_CTf_f_Int_t sc_0_16_destruct_d;
  logic sc_0_16_destruct_r;
  Pointer_MaskQTree_t q1ae8_1_destruct_d;
  logic q1ae8_1_destruct_r;
  Pointer_QTree_Int_t \q1'aen_1_destruct_d ;
  logic \q1'aen_1_destruct_r ;
  Pointer_QTree_Int_t t1aes_1_destruct_d;
  logic t1aes_1_destruct_r;
  MyDTInt_Bool_t is_zae6_2_destruct_d;
  logic is_zae6_2_destruct_r;
  MyDTInt_Int_Int_t op_addae7_2_destruct_d;
  logic op_addae7_2_destruct_r;
  Pointer_MaskQTree_t q2ae9_1_destruct_d;
  logic q2ae9_1_destruct_r;
  Pointer_QTree_Int_t \q2'aeo_1_destruct_d ;
  logic \q2'aeo_1_destruct_r ;
  Pointer_QTree_Int_t t2aet_1_destruct_d;
  logic t2aet_1_destruct_r;
  Pointer_MaskQTree_t q3aea_1_destruct_d;
  logic q3aea_1_destruct_r;
  Pointer_QTree_Int_t \q3'aep_1_destruct_d ;
  logic \q3'aep_1_destruct_r ;
  Pointer_QTree_Int_t t3aeu_1_destruct_d;
  logic t3aeu_1_destruct_r;
  CTf_f_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  CTf_f_Int_t lizzieLet60_1Lcall_f_f_Int3_d;
  logic lizzieLet60_1Lcall_f_f_Int3_r;
  CTf_f_Int_t lizzieLet60_1Lcall_f_f_Int2_d;
  logic lizzieLet60_1Lcall_f_f_Int2_r;
  CTf_f_Int_t lizzieLet60_1Lcall_f_f_Int1_d;
  logic lizzieLet60_1Lcall_f_f_Int1_r;
  CTf_f_Int_t lizzieLet60_1Lcall_f_f_Int0_d;
  logic lizzieLet60_1Lcall_f_f_Int0_r;
  Go_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Go_t lizzieLet60_3Lcall_f_f_Int3_d;
  logic lizzieLet60_3Lcall_f_f_Int3_r;
  Go_t lizzieLet60_3Lcall_f_f_Int2_d;
  logic lizzieLet60_3Lcall_f_f_Int2_r;
  Go_t lizzieLet60_3Lcall_f_f_Int1_d;
  logic lizzieLet60_3Lcall_f_f_Int1_r;
  Go_t lizzieLet60_3Lcall_f_f_Int0_d;
  logic lizzieLet60_3Lcall_f_f_Int0_r;
  Go_t lizzieLet60_3Lcall_f_f_Int0_1_argbuf_d;
  logic lizzieLet60_3Lcall_f_f_Int0_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f_f_Int1_1_argbuf_d;
  logic lizzieLet60_3Lcall_f_f_Int1_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f_f_Int2_1_argbuf_d;
  logic lizzieLet60_3Lcall_f_f_Int2_1_argbuf_r;
  Go_t lizzieLet60_3Lcall_f_f_Int3_1_argbuf_d;
  logic lizzieLet60_3Lcall_f_f_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet60_4Lf_f_Intsbos_d;
  logic lizzieLet60_4Lf_f_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet60_4Lcall_f_f_Int3_d;
  logic lizzieLet60_4Lcall_f_f_Int3_r;
  Pointer_QTree_Int_t lizzieLet60_4Lcall_f_f_Int2_d;
  logic lizzieLet60_4Lcall_f_f_Int2_r;
  Pointer_QTree_Int_t lizzieLet60_4Lcall_f_f_Int1_d;
  logic lizzieLet60_4Lcall_f_f_Int1_r;
  Pointer_QTree_Int_t lizzieLet60_4Lcall_f_f_Int0_d;
  logic lizzieLet60_4Lcall_f_f_Int0_r;
  QTree_Int_t lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d;
  logic lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r;
  QTree_Int_t lizzieLet64_1_argbuf_d;
  logic lizzieLet64_1_argbuf_r;
  CTf_f_Int_t lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_d;
  logic lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_r;
  CTf_f_Int_t lizzieLet63_1_argbuf_d;
  logic lizzieLet63_1_argbuf_r;
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_d ;
  logic \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_r ;
  CTf_f_Int_t lizzieLet62_1_argbuf_d;
  logic lizzieLet62_1_argbuf_r;
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_d ;
  logic \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_r ;
  CTf_f_Int_t lizzieLet61_1_argbuf_d;
  logic lizzieLet61_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_f_f_Int_goConst_d;
  logic call_f_f_Int_goConst_r;
  Pointer_QTree_Int_t f_f_Int_resbuf_d;
  logic f_f_Int_resbuf_r;
  Pointer_MaskQTree_t q1aey_destruct_d;
  logic q1aey_destruct_r;
  Pointer_MaskQTree_t q2aez_destruct_d;
  logic q2aez_destruct_r;
  Pointer_MaskQTree_t q3aeA_destruct_d;
  logic q3aeA_destruct_r;
  Pointer_MaskQTree_t q5aeB_destruct_d;
  logic q5aeB_destruct_r;
  MaskQTree_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  MaskQTree_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  MaskQTree_t lizzieLet6_1MQNode_d;
  logic lizzieLet6_1MQNode_r;
  Go_t lizzieLet6_3MQNone_d;
  logic lizzieLet6_3MQNone_r;
  Go_t lizzieLet6_3MQVal_d;
  logic lizzieLet6_3MQVal_r;
  Go_t lizzieLet6_3MQNode_d;
  logic lizzieLet6_3MQNode_r;
  Go_t lizzieLet6_3MQNone_1_d;
  logic lizzieLet6_3MQNone_1_r;
  Go_t lizzieLet6_3MQNone_2_d;
  logic lizzieLet6_3MQNone_2_r;
  QTree_Int_t lizzieLet6_3MQNone_1QNone_Int_d;
  logic lizzieLet6_3MQNone_1QNone_Int_r;
  QTree_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_3MQNone_2_argbuf_d;
  logic lizzieLet6_3MQNone_2_argbuf_r;
  C6_t go_16_goMux_choice_d;
  logic go_16_goMux_choice_r;
  Go_t go_16_goMux_data_d;
  logic go_16_goMux_data_r;
  Go_t lizzieLet6_3MQVal_1_argbuf_d;
  logic lizzieLet6_3MQVal_1_argbuf_r;
  QTree_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  QTree_Int_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  QTree_Int_t lizzieLet6_4MQNode_d;
  logic lizzieLet6_4MQNode_r;
  QTree_Int_t lizzieLet6_4MQNode_1_d;
  logic lizzieLet6_4MQNode_1_r;
  QTree_Int_t lizzieLet6_4MQNode_2_d;
  logic lizzieLet6_4MQNode_2_r;
  QTree_Int_t lizzieLet6_4MQNode_3_d;
  logic lizzieLet6_4MQNode_3_r;
  QTree_Int_t lizzieLet6_4MQNode_4_d;
  logic lizzieLet6_4MQNode_4_r;
  QTree_Int_t lizzieLet6_4MQNode_5_d;
  logic lizzieLet6_4MQNode_5_r;
  QTree_Int_t lizzieLet6_4MQNode_6_d;
  logic lizzieLet6_4MQNode_6_r;
  QTree_Int_t lizzieLet6_4MQNode_7_d;
  logic lizzieLet6_4MQNode_7_r;
  QTree_Int_t lizzieLet6_4MQNode_8_d;
  logic lizzieLet6_4MQNode_8_r;
  Pointer_QTree_Int_t t1aeD_destruct_d;
  logic t1aeD_destruct_r;
  Pointer_QTree_Int_t t2aeE_destruct_d;
  logic t2aeE_destruct_r;
  Pointer_QTree_Int_t t3aeF_destruct_d;
  logic t3aeF_destruct_r;
  Pointer_QTree_Int_t t4aeG_destruct_d;
  logic t4aeG_destruct_r;
  QTree_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  QTree_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  QTree_Int_t lizzieLet6_4MQNode_1QNode_Int_d;
  logic lizzieLet6_4MQNode_1QNode_Int_r;
  QTree_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  Go_t lizzieLet6_4MQNode_3QNone_Int_d;
  logic lizzieLet6_4MQNode_3QNone_Int_r;
  Go_t lizzieLet6_4MQNode_3QVal_Int_d;
  logic lizzieLet6_4MQNode_3QVal_Int_r;
  Go_t lizzieLet6_4MQNode_3QNode_Int_d;
  logic lizzieLet6_4MQNode_3QNode_Int_r;
  Go_t lizzieLet6_4MQNode_3QError_Int_d;
  logic lizzieLet6_4MQNode_3QError_Int_r;
  Go_t lizzieLet6_4MQNode_3QError_Int_1_d;
  logic lizzieLet6_4MQNode_3QError_Int_1_r;
  Go_t lizzieLet6_4MQNode_3QError_Int_2_d;
  logic lizzieLet6_4MQNode_3QError_Int_2_r;
  QTree_Int_t lizzieLet6_4MQNode_3QError_Int_1QError_Int_d;
  logic lizzieLet6_4MQNode_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QError_Int_2_argbuf_d;
  logic lizzieLet6_4MQNode_3QError_Int_2_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QNode_Int_1_argbuf_d;
  logic lizzieLet6_4MQNode_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QNone_Int_1_d;
  logic lizzieLet6_4MQNode_3QNone_Int_1_r;
  Go_t lizzieLet6_4MQNode_3QNone_Int_2_d;
  logic lizzieLet6_4MQNode_3QNone_Int_2_r;
  QTree_Int_t lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_d;
  logic lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QNone_Int_2_argbuf_d;
  logic lizzieLet6_4MQNode_3QNone_Int_2_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QVal_Int_1_d;
  logic lizzieLet6_4MQNode_3QVal_Int_1_r;
  Go_t lizzieLet6_4MQNode_3QVal_Int_2_d;
  logic lizzieLet6_4MQNode_3QVal_Int_2_r;
  QTree_Int_t lizzieLet6_4MQNode_3QVal_Int_1QError_Int_d;
  logic lizzieLet6_4MQNode_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Go_t lizzieLet6_4MQNode_3QVal_Int_2_argbuf_d;
  logic lizzieLet6_4MQNode_3QVal_Int_2_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QNone_Int_d;
  logic lizzieLet6_4MQNode_4QNone_Int_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QVal_Int_d;
  logic lizzieLet6_4MQNode_4QVal_Int_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QNode_Int_d;
  logic lizzieLet6_4MQNode_4QNode_Int_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QError_Int_d;
  logic lizzieLet6_4MQNode_4QError_Int_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QError_Int_1_argbuf_d;
  logic lizzieLet6_4MQNode_4QError_Int_1_argbuf_r;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_d ;
  logic \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QNone_Int_1_argbuf_d;
  logic lizzieLet6_4MQNode_4QNone_Int_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_4MQNode_4QVal_Int_1_argbuf_r;
  Pointer_MaskQTree_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Pointer_MaskQTree_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_5QNode_Int_d;
  logic lizzieLet6_4MQNode_5QNode_Int_r;
  Pointer_MaskQTree_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  Pointer_MaskQTree_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  Pointer_MaskQTree_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_6QNode_Int_d;
  logic lizzieLet6_4MQNode_6QNode_Int_r;
  Pointer_MaskQTree_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_MaskQTree_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Pointer_MaskQTree_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_7QNode_Int_d;
  logic lizzieLet6_4MQNode_7QNode_Int_r;
  Pointer_MaskQTree_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_MaskQTree_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_MaskQTree_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_8QNode_Int_d;
  logic lizzieLet6_4MQNode_8QNode_Int_r;
  Pointer_MaskQTree_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_8QNode_Int_1_argbuf_d;
  logic lizzieLet6_4MQNode_8QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5MQVal_d;
  logic lizzieLet6_5MQVal_r;
  Pointer_QTree_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet6_5MQVal_1_argbuf_d;
  logic lizzieLet6_5MQVal_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQNone_d;
  logic lizzieLet6_6MQNone_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQVal_d;
  logic lizzieLet6_6MQVal_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQNode_d;
  logic lizzieLet6_6MQNode_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQNone_1_argbuf_d;
  logic lizzieLet6_6MQNone_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQVal_1_argbuf_d;
  logic lizzieLet6_6MQVal_1_argbuf_r;
  Pointer_MaskQTree_t m1ae3_1_argbuf_d;
  logic m1ae3_1_argbuf_r;
  Pointer_QTree_Int_t m2ae4_1_argbuf_d;
  logic m2ae4_1_argbuf_r;
  Pointer_QTree_Int_t m2ae4_1_d;
  logic m2ae4_1_r;
  Pointer_QTree_Int_t m2ae4_2_d;
  logic m2ae4_2_r;
  Pointer_QTree_Int_t m2aeH_1_argbuf_d;
  logic m2aeH_1_argbuf_r;
  Pointer_QTree_Int_t m2aeH_1_d;
  logic m2aeH_1_r;
  Pointer_QTree_Int_t m2aeH_2_d;
  logic m2aeH_2_r;
  Pointer_QTree_Int_t m3ae5_1_argbuf_d;
  logic m3ae5_1_argbuf_r;
  Pointer_QTree_Int_t m3ae5_1_d;
  logic m3ae5_1_r;
  Pointer_QTree_Int_t m3ae5_2_d;
  logic m3ae5_2_r;
  Pointer_QTree_Int_t m3aeI_1_argbuf_d;
  logic m3aeI_1_argbuf_r;
  Pointer_QTree_Int_t m3aeI_1_d;
  logic m3aeI_1_r;
  Pointer_QTree_Int_t m3aeI_2_d;
  logic m3aeI_2_r;
  MyDTInt_Int_Int_t op_addae7_2_2_argbuf_d;
  logic op_addae7_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_addae7_2_1_d;
  logic op_addae7_2_1_r;
  MyDTInt_Int_Int_t op_addae7_2_2_d;
  logic op_addae7_2_2_r;
  MyDTInt_Int_Int_t op_addae7_3_2_argbuf_d;
  logic op_addae7_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_addae7_3_1_d;
  logic op_addae7_3_1_r;
  MyDTInt_Int_Int_t op_addae7_3_2_d;
  logic op_addae7_3_2_r;
  MyDTInt_Int_Int_t op_addae7_4_1_argbuf_d;
  logic op_addae7_4_1_argbuf_r;
  MyDTInt_Int_Int_t op_addaeK_2_2_argbuf_d;
  logic op_addaeK_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_addaeK_2_1_d;
  logic op_addaeK_2_1_r;
  MyDTInt_Int_Int_t op_addaeK_2_2_d;
  logic op_addaeK_2_2_r;
  MyDTInt_Int_Int_t op_addaeK_3_2_argbuf_d;
  logic op_addaeK_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_addaeK_3_1_d;
  logic op_addaeK_3_1_r;
  MyDTInt_Int_Int_t op_addaeK_3_2_d;
  logic op_addaeK_3_2_r;
  MyDTInt_Int_Int_t op_addaeK_4_1_argbuf_d;
  logic op_addaeK_4_1_argbuf_r;
  Pointer_QTree_Int_t \q1'aen_3_1_argbuf_d ;
  logic \q1'aen_3_1_argbuf_r ;
  Pointer_QTree_Int_t q1a85_1_argbuf_d;
  logic q1a85_1_argbuf_r;
  Pointer_MaskQTree_t q1ae8_3_1_argbuf_d;
  logic q1ae8_3_1_argbuf_r;
  Pointer_QTree_Int_t q1aeR_3_1_argbuf_d;
  logic q1aeR_3_1_argbuf_r;
  Pointer_MaskQTree_t q1aey_3_1_argbuf_d;
  logic q1aey_3_1_argbuf_r;
  Pointer_QTree_Int_t \q2'aeo_2_1_argbuf_d ;
  logic \q2'aeo_2_1_argbuf_r ;
  Pointer_QTree_Int_t q2a86_1_1_argbuf_d;
  logic q2a86_1_1_argbuf_r;
  Pointer_MaskQTree_t q2ae9_2_1_argbuf_d;
  logic q2ae9_2_1_argbuf_r;
  Pointer_QTree_Int_t q2aeS_2_1_argbuf_d;
  logic q2aeS_2_1_argbuf_r;
  Pointer_MaskQTree_t q2aez_2_1_argbuf_d;
  logic q2aez_2_1_argbuf_r;
  Pointer_QTree_Int_t \q3'aep_1_1_argbuf_d ;
  logic \q3'aep_1_1_argbuf_r ;
  Pointer_QTree_Int_t q3a87_2_1_argbuf_d;
  logic q3a87_2_1_argbuf_r;
  Pointer_MaskQTree_t q3aeA_1_1_argbuf_d;
  logic q3aeA_1_1_argbuf_r;
  Pointer_QTree_Int_t q3aeT_1_1_argbuf_d;
  logic q3aeT_1_1_argbuf_r;
  Pointer_MaskQTree_t q3aea_1_1_argbuf_d;
  logic q3aea_1_1_argbuf_r;
  Pointer_QTree_Int_t \q4'aex_1_argbuf_d ;
  logic \q4'aex_1_argbuf_r ;
  Pointer_QTree_Int_t \q4'aex_1_d ;
  logic \q4'aex_1_r ;
  Pointer_QTree_Int_t \q4'aex_2_d ;
  logic \q4'aex_2_r ;
  Pointer_QTree_Int_t q4a88_3_1_argbuf_d;
  logic q4a88_3_1_argbuf_r;
  Pointer_MaskQTree_t q4aew_1_argbuf_d;
  logic q4aew_1_argbuf_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_Int_t lizzieLet46_1_d;
  logic lizzieLet46_1_r;
  CT$wnnz_Int_t lizzieLet46_2_d;
  logic lizzieLet46_2_r;
  CT$wnnz_Int_t lizzieLet46_3_d;
  logic lizzieLet46_3_r;
  CT$wnnz_Int_t lizzieLet46_4_d;
  logic lizzieLet46_4_r;
  \CTf'''''''''_f'''''''''_Int_t  \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_r ;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet50_1_d;
  logic lizzieLet50_1_r;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet50_2_d;
  logic lizzieLet50_2_r;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet50_3_d;
  logic lizzieLet50_3_r;
  \CTf'''''''''_f'''''''''_Int_t  lizzieLet50_4_d;
  logic lizzieLet50_4_r;
  \CTf'_f'_Int_t  \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_r ;
  \CTf'_f'_Int_t  lizzieLet55_1_d;
  logic lizzieLet55_1_r;
  \CTf'_f'_Int_t  lizzieLet55_2_d;
  logic lizzieLet55_2_r;
  \CTf'_f'_Int_t  lizzieLet55_3_d;
  logic lizzieLet55_3_r;
  \CTf'_f'_Int_t  lizzieLet55_4_d;
  logic lizzieLet55_4_r;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d;
  logic readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_r;
  CTf_f_Int_t lizzieLet60_1_d;
  logic lizzieLet60_1_r;
  CTf_f_Int_t lizzieLet60_2_d;
  logic lizzieLet60_2_r;
  CTf_f_Int_t lizzieLet60_3_d;
  logic lizzieLet60_3_r;
  CTf_f_Int_t lizzieLet60_4_d;
  logic lizzieLet60_4_r;
  MaskQTree_t readPointer_MaskQTreem1ae3_1_argbuf_rwb_d;
  logic readPointer_MaskQTreem1ae3_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet24_1_d;
  logic lizzieLet24_1_r;
  MaskQTree_t lizzieLet24_2_d;
  logic lizzieLet24_2_r;
  MaskQTree_t lizzieLet24_3_d;
  logic lizzieLet24_3_r;
  MaskQTree_t lizzieLet24_4_d;
  logic lizzieLet24_4_r;
  MaskQTree_t lizzieLet24_5_d;
  logic lizzieLet24_5_r;
  MaskQTree_t lizzieLet24_6_d;
  logic lizzieLet24_6_r;
  MaskQTree_t lizzieLet24_7_d;
  logic lizzieLet24_7_r;
  MaskQTree_t lizzieLet24_8_d;
  logic lizzieLet24_8_r;
  MaskQTree_t lizzieLet24_9_d;
  logic lizzieLet24_9_r;
  MaskQTree_t lizzieLet24_10_d;
  logic lizzieLet24_10_r;
  MaskQTree_t readPointer_MaskQTreeq4aew_1_argbuf_rwb_d;
  logic readPointer_MaskQTreeq4aew_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  MaskQTree_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  MaskQTree_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  MaskQTree_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  MaskQTree_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  MaskQTree_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t readPointer_QTree_Intm2ae4_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2ae4_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intm2aeH_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2aeH_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet13_1_d;
  logic lizzieLet13_1_r;
  QTree_Int_t lizzieLet13_2_d;
  logic lizzieLet13_2_r;
  QTree_Int_t lizzieLet13_3_d;
  logic lizzieLet13_3_r;
  QTree_Int_t lizzieLet13_4_d;
  logic lizzieLet13_4_r;
  QTree_Int_t lizzieLet13_5_d;
  logic lizzieLet13_5_r;
  QTree_Int_t lizzieLet13_6_d;
  logic lizzieLet13_6_r;
  QTree_Int_t lizzieLet13_7_d;
  logic lizzieLet13_7_r;
  QTree_Int_t lizzieLet13_8_d;
  logic lizzieLet13_8_r;
  QTree_Int_t lizzieLet13_9_d;
  logic lizzieLet13_9_r;
  QTree_Int_t readPointer_QTree_Intm3ae5_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm3ae5_1_argbuf_rwb_r;
  QTree_Int_t readPointer_QTree_Intm3aeI_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm3aeI_1_argbuf_rwb_r;
  QTree_Int_t \readPointer_QTree_Intq4'aex_1_argbuf_rwb_d ;
  logic \readPointer_QTree_Intq4'aex_1_argbuf_rwb_r ;
  QTree_Int_t readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d;
  logic readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_11_1_argbuf_d;
  logic sc_0_11_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  sc_0_15_1_argbuf_d;
  logic sc_0_15_1_argbuf_r;
  Pointer_CTf_f_Int_t sc_0_19_1_argbuf_d;
  logic sc_0_19_1_argbuf_r;
  Pointer_CT$wnnz_Int_t sc_0_7_1_argbuf_d;
  logic sc_0_7_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CTf_f_Int_t scfarg_0_3_1_argbuf_d;
  logic scfarg_0_3_1_argbuf_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1aeD_3_1_argbuf_d;
  logic t1aeD_3_1_argbuf_r;
  Pointer_QTree_Int_t t1aeW_3_1_argbuf_d;
  logic t1aeW_3_1_argbuf_r;
  Pointer_QTree_Int_t t1aed_1_argbuf_d;
  logic t1aed_1_argbuf_r;
  Pointer_QTree_Int_t t1aes_3_1_argbuf_d;
  logic t1aes_3_1_argbuf_r;
  Pointer_QTree_Int_t t2aeE_2_1_argbuf_d;
  logic t2aeE_2_1_argbuf_r;
  Pointer_QTree_Int_t t2aeX_2_1_argbuf_d;
  logic t2aeX_2_1_argbuf_r;
  Pointer_QTree_Int_t t2aee_1_argbuf_d;
  logic t2aee_1_argbuf_r;
  Pointer_QTree_Int_t t2aet_2_1_argbuf_d;
  logic t2aet_2_1_argbuf_r;
  Pointer_QTree_Int_t t3aeF_1_1_argbuf_d;
  logic t3aeF_1_1_argbuf_r;
  Pointer_QTree_Int_t t3aeY_1_1_argbuf_d;
  logic t3aeY_1_1_argbuf_r;
  Pointer_QTree_Int_t t3aef_1_argbuf_d;
  logic t3aef_1_argbuf_r;
  Pointer_QTree_Int_t t3aeu_1_1_argbuf_d;
  logic t3aeu_1_1_argbuf_r;
  Pointer_QTree_Int_t t4aeG_1_argbuf_d;
  logic t4aeG_1_argbuf_r;
  Pointer_QTree_Int_t t4aeZ_1_argbuf_d;
  logic t4aeZ_1_argbuf_r;
  Pointer_QTree_Int_t t4aeg_1_argbuf_d;
  logic t4aeg_1_argbuf_r;
  Pointer_QTree_Int_t t4aev_1_argbuf_d;
  logic t4aev_1_argbuf_r;
  Int_t vaeM_1_argbuf_d;
  logic vaeM_1_argbuf_r;
  Int_t vaeM_1_d;
  logic vaeM_1_r;
  Int_t vaeM_2_d;
  logic vaeM_2_r;
  Int_t vaei_1_argbuf_d;
  logic vaei_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_r ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_t  lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet40_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca3_3_1_argbuf_d;
  logic sca3_3_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet45_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t lizzieLet27_1_1_argbuf_d;
  logic lizzieLet27_1_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet61_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca2_3_1_argbuf_d;
  logic sca2_3_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet62_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca1_3_1_argbuf_d;
  logic sca1_3_1_argbuf_r;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_rwb_d;
  logic writeCTf_f_IntlizzieLet63_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_t sca0_3_1_argbuf_d;
  logic sca0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet12_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet28_2_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet15_1_1_argbuf_d;
  logic lizzieLet15_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet29_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet16_1_1_argbuf_d;
  logic lizzieLet16_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet30_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet17_1_1_argbuf_d;
  logic lizzieLet17_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet18_1_1_argbuf_d;
  logic lizzieLet18_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet33_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet19_1_1_argbuf_d;
  logic lizzieLet19_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet20_1_1_argbuf_d;
  logic lizzieLet20_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet21_1_1_argbuf_d;
  logic lizzieLet21_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet22_1_1_argbuf_d;
  logic lizzieLet22_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet23_1_1_argbuf_d;
  logic lizzieLet23_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet24_1_1_argbuf_d;
  logic lizzieLet24_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet25_1_1_argbuf_d;
  logic lizzieLet25_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet26_1_1_argbuf_d;
  logic lizzieLet26_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet59_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet64_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_3_1_argbuf_d;
  logic contRet_0_3_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t wsjQ_1_1_argbuf_d;
  logic wsjQ_1_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet48_1_argbuf_d;
  logic lizzieLet48_1_argbuf_r;
  CT$wnnz_Int_t wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_d;
  logic wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet49_1_argbuf_d;
  logic lizzieLet49_1_argbuf_r;
  CT$wnnz_Int_t wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  logic wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r;
  \Int#_t  es_6_2_1ww2Xku_1_1_Add32_d;
  logic es_6_2_1ww2Xku_1_1_Add32_r;
  \Int#_t  wwsjT_4_1ww1Xkr_2_1_Add32_d;
  logic wwsjT_4_1ww1Xkr_2_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go),
                                (go__11,Go),
                                (go__12,Go)] */
  logic [11:0] sourceGo_emitted;
  logic [11:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign go__11_d = (sourceGo_d[0] && (! sourceGo_emitted[10]));
  assign go__12_d = (sourceGo_d[0] && (! sourceGo_emitted[11]));
  assign sourceGo_done = (sourceGo_emitted | ({go__12_d[0],
                                               go__11_d[0],
                                               go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__12_r,
                                                             go__11_r,
                                                             go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 12'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 12'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go__5,Go) > (initHP_CT$wnnz_Int,Word16#) */
  assign initHP_CT$wnnz_Int_d = {16'd0, go__5_d[0]};
  assign go__5_r = initHP_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz_Int1,Go) > (incrHP_CT$wnnz_Int,Word16#) */
  assign incrHP_CT$wnnz_Int_d = {16'd1, incrHP_CT$wnnz_Int1_d[0]};
  assign incrHP_CT$wnnz_Int1_r = incrHP_CT$wnnz_Int_r;
  
  /* merge (Ty Go) : [(go__6,Go),
                 (incrHP_CT$wnnz_Int2,Go)] > (incrHP_mergeCT$wnnz_Int,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_Int_selected;
  logic [1:0] incrHP_mergeCT$wnnz_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_Int_select))
        incrHP_mergeCT$wnnz_Int_selected = incrHP_mergeCT$wnnz_Int_select;
      else
        if (go__6_d[0]) incrHP_mergeCT$wnnz_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz_Int2_d[0])
          incrHP_mergeCT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_select <= (incrHP_mergeCT$wnnz_Int_r ? 2'd0 :
                                         incrHP_mergeCT$wnnz_Int_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_Int_selected[0])
      incrHP_mergeCT$wnnz_Int_d = go__6_d;
    else if (incrHP_mergeCT$wnnz_Int_selected[1])
      incrHP_mergeCT$wnnz_Int_d = incrHP_CT$wnnz_Int2_d;
    else incrHP_mergeCT$wnnz_Int_d = 1'd0;
  assign {incrHP_CT$wnnz_Int2_r,
          go__6_r} = (incrHP_mergeCT$wnnz_Int_r ? incrHP_mergeCT$wnnz_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_Int_buf,Go) > [(incrHP_CT$wnnz_Int1,Go),
                                                   (incrHP_CT$wnnz_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_done;
  assign incrHP_CT$wnnz_Int1_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[0]));
  assign incrHP_CT$wnnz_Int2_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_Int_buf_done = (incrHP_mergeCT$wnnz_Int_buf_emitted | ({incrHP_CT$wnnz_Int2_d[0],
                                                                                     incrHP_CT$wnnz_Int1_d[0]} & {incrHP_CT$wnnz_Int2_r,
                                                                                                                  incrHP_CT$wnnz_Int1_r}));
  assign incrHP_mergeCT$wnnz_Int_buf_r = (& incrHP_mergeCT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_buf_emitted <= (incrHP_mergeCT$wnnz_Int_buf_r ? 2'd0 :
                                              incrHP_mergeCT$wnnz_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz_Int,Word16#) (forkHP1_CT$wnnz_Int,Word16#) > (addHP_CT$wnnz_Int,Word16#) */
  assign addHP_CT$wnnz_Int_d = {(incrHP_CT$wnnz_Int_d[16:1] + forkHP1_CT$wnnz_Int_d[16:1]),
                                (incrHP_CT$wnnz_Int_d[0] && forkHP1_CT$wnnz_Int_d[0])};
  assign {incrHP_CT$wnnz_Int_r,
          forkHP1_CT$wnnz_Int_r} = {2 {(addHP_CT$wnnz_Int_r && addHP_CT$wnnz_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz_Int,Word16#),
                      (addHP_CT$wnnz_Int,Word16#)] > (mergeHP_CT$wnnz_Int,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_Int_selected;
  logic [1:0] mergeHP_CT$wnnz_Int_select;
  always_comb
    begin
      mergeHP_CT$wnnz_Int_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_Int_select))
        mergeHP_CT$wnnz_Int_selected = mergeHP_CT$wnnz_Int_select;
      else
        if (initHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_select <= 2'd0;
    else
      mergeHP_CT$wnnz_Int_select <= (mergeHP_CT$wnnz_Int_r ? 2'd0 :
                                     mergeHP_CT$wnnz_Int_selected);
  always_comb
    if (mergeHP_CT$wnnz_Int_selected[0])
      mergeHP_CT$wnnz_Int_d = initHP_CT$wnnz_Int_d;
    else if (mergeHP_CT$wnnz_Int_selected[1])
      mergeHP_CT$wnnz_Int_d = addHP_CT$wnnz_Int_d;
    else mergeHP_CT$wnnz_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_Int_r,
          initHP_CT$wnnz_Int_r} = (mergeHP_CT$wnnz_Int_r ? mergeHP_CT$wnnz_Int_selected :
                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz_Int,Go) > (incrHP_mergeCT$wnnz_Int_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_d;
  logic incrHP_mergeCT$wnnz_Int_bufchan_r;
  assign incrHP_mergeCT$wnnz_Int_r = ((! incrHP_mergeCT$wnnz_Int_bufchan_d[0]) || incrHP_mergeCT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_Int_r)
        incrHP_mergeCT$wnnz_Int_bufchan_d <= incrHP_mergeCT$wnnz_Int_d;
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_buf;
  assign incrHP_mergeCT$wnnz_Int_bufchan_r = (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_Int_buf_d = (incrHP_mergeCT$wnnz_Int_bufchan_buf[0] ? incrHP_mergeCT$wnnz_Int_bufchan_buf :
                                          incrHP_mergeCT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_Int_buf_r && incrHP_mergeCT$wnnz_Int_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_Int_buf_r) && (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= incrHP_mergeCT$wnnz_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz_Int,Word16#) > (mergeHP_CT$wnnz_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_d;
  logic mergeHP_CT$wnnz_Int_bufchan_r;
  assign mergeHP_CT$wnnz_Int_r = ((! mergeHP_CT$wnnz_Int_bufchan_d[0]) || mergeHP_CT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_Int_r)
        mergeHP_CT$wnnz_Int_bufchan_d <= mergeHP_CT$wnnz_Int_d;
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_buf;
  assign mergeHP_CT$wnnz_Int_bufchan_r = (! mergeHP_CT$wnnz_Int_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_Int_buf_d = (mergeHP_CT$wnnz_Int_bufchan_buf[0] ? mergeHP_CT$wnnz_Int_bufchan_buf :
                                      mergeHP_CT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_Int_buf_r && mergeHP_CT$wnnz_Int_bufchan_buf[0]))
        mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_Int_buf_r) && (! mergeHP_CT$wnnz_Int_bufchan_buf[0])))
        mergeHP_CT$wnnz_Int_bufchan_buf <= mergeHP_CT$wnnz_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_Int_buf,Word16#) > [(forkHP1_CT$wnnz_Int,Word16#),
                                                         (forkHP1_CT$wnnz_In2,Word16#),
                                                         (forkHP1_CT$wnnz_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_Int_buf_done;
  assign forkHP1_CT$wnnz_Int_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[0]))};
  assign forkHP1_CT$wnnz_In2_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[1]))};
  assign forkHP1_CT$wnnz_In3_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_Int_buf_done = (mergeHP_CT$wnnz_Int_buf_emitted | ({forkHP1_CT$wnnz_In3_d[0],
                                                                             forkHP1_CT$wnnz_In2_d[0],
                                                                             forkHP1_CT$wnnz_Int_d[0]} & {forkHP1_CT$wnnz_In3_r,
                                                                                                          forkHP1_CT$wnnz_In2_r,
                                                                                                          forkHP1_CT$wnnz_Int_r}));
  assign mergeHP_CT$wnnz_Int_buf_r = (& mergeHP_CT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_Int_buf_emitted <= (mergeHP_CT$wnnz_Int_buf_r ? 3'd0 :
                                          mergeHP_CT$wnnz_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz_Int) : [(dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int),
                                    (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int)] > (memMergeChoice_CT$wnnz_Int,C2) (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  logic [1:0] dconReadIn_CT$wnnz_Int_select_d;
  assign dconReadIn_CT$wnnz_Int_select_d = ((| dconReadIn_CT$wnnz_Int_select_q) ? dconReadIn_CT$wnnz_Int_select_q :
                                            (dconReadIn_CT$wnnz_Int_d[0] ? 2'd1 :
                                             (dconWriteIn_CT$wnnz_Int_d[0] ? 2'd2 :
                                              2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_select_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                          dconReadIn_CT$wnnz_Int_select_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_emit_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                        dconReadIn_CT$wnnz_Int_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_d;
  assign dconReadIn_CT$wnnz_Int_emit_d = (dconReadIn_CT$wnnz_Int_emit_q | ({memMergeChoice_CT$wnnz_Int_d[0],
                                                                            memMergeIn_CT$wnnz_Int_d[0]} & {memMergeChoice_CT$wnnz_Int_r,
                                                                                                            memMergeIn_CT$wnnz_Int_r}));
  logic dconReadIn_CT$wnnz_Int_done;
  assign dconReadIn_CT$wnnz_Int_done = (& dconReadIn_CT$wnnz_Int_emit_d);
  assign {dconWriteIn_CT$wnnz_Int_r,
          dconReadIn_CT$wnnz_Int_r} = (dconReadIn_CT$wnnz_Int_done ? dconReadIn_CT$wnnz_Int_select_d :
                                       2'd0);
  assign memMergeIn_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconReadIn_CT$wnnz_Int_d :
                                     ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconWriteIn_CT$wnnz_Int_d :
                                      {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz_Int,
      Ty MemOut_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) > (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) */
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_din;
  logic [114:0] memOut_CT$wnnz_Int_q;
  logic memOut_CT$wnnz_Int_valid;
  logic memMergeIn_CT$wnnz_Int_dbuf_we;
  logic memOut_CT$wnnz_Int_we;
  assign memMergeIn_CT$wnnz_Int_dbuf_din = memMergeIn_CT$wnnz_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_Int_dbuf_address = memMergeIn_CT$wnnz_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_Int_dbuf_we = (memMergeIn_CT$wnnz_Int_dbuf_d[1:1] && memMergeIn_CT$wnnz_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_Int_we <= 1'd0;
        memOut_CT$wnnz_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_Int_we <= memMergeIn_CT$wnnz_Int_dbuf_we;
        memOut_CT$wnnz_Int_valid <= memMergeIn_CT$wnnz_Int_dbuf_d[0];
        if (memMergeIn_CT$wnnz_Int_dbuf_we)
          begin
            memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address] <= memMergeIn_CT$wnnz_Int_dbuf_din;
            memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_din;
          end
        else
          memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address];
      end
  assign memOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_q,
                                 memOut_CT$wnnz_Int_we,
                                 memOut_CT$wnnz_Int_valid};
  assign memMergeIn_CT$wnnz_Int_dbuf_r = ((! memOut_CT$wnnz_Int_valid) || memOut_CT$wnnz_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz_Int) : (memMergeChoice_CT$wnnz_Int,C2) (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) > [(memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int),
                                                                                                                (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int)] */
  logic [1:0] memOut_CT$wnnz_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_Int_d[0] && memOut_CT$wnnz_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_Int_d[1:1])
        1'd0: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                     memOut_CT$wnnz_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                      memOut_CT$wnnz_Int_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_Int_dbuf_r = (| (memOut_CT$wnnz_Int_dbuf_onehotd & {memWriteOut_CT$wnnz_Int_r,
                                                                            memReadOut_CT$wnnz_Int_r}));
  assign memMergeChoice_CT$wnnz_Int_r = memOut_CT$wnnz_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) */
  assign memMergeIn_CT$wnnz_Int_rbuf_r = ((! memMergeIn_CT$wnnz_Int_dbuf_d[0]) || memMergeIn_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wnnz_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_Int_rbuf_r)
        memMergeIn_CT$wnnz_Int_dbuf_d <= memMergeIn_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) */
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_buf;
  assign memMergeIn_CT$wnnz_Int_r = (! memMergeIn_CT$wnnz_Int_buf[0]);
  assign memMergeIn_CT$wnnz_Int_rbuf_d = (memMergeIn_CT$wnnz_Int_buf[0] ? memMergeIn_CT$wnnz_Int_buf :
                                          memMergeIn_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_Int_rbuf_r && memMergeIn_CT$wnnz_Int_buf[0]))
        memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_Int_rbuf_r) && (! memMergeIn_CT$wnnz_Int_buf[0])))
        memMergeIn_CT$wnnz_Int_buf <= memMergeIn_CT$wnnz_Int_d;
  
  /* dbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) */
  assign memOut_CT$wnnz_Int_rbuf_r = ((! memOut_CT$wnnz_Int_dbuf_d[0]) || memOut_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_Int_rbuf_r)
        memOut_CT$wnnz_Int_dbuf_d <= memOut_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) */
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_buf;
  assign memOut_CT$wnnz_Int_r = (! memOut_CT$wnnz_Int_buf[0]);
  assign memOut_CT$wnnz_Int_rbuf_d = (memOut_CT$wnnz_Int_buf[0] ? memOut_CT$wnnz_Int_buf :
                                      memOut_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_Int_rbuf_r && memOut_CT$wnnz_Int_buf[0]))
        memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_Int_rbuf_r) && (! memOut_CT$wnnz_Int_buf[0])))
        memOut_CT$wnnz_Int_buf <= memOut_CT$wnnz_Int_d;
  
  /* destruct (Ty Pointer_CT$wnnz_Int,
          Dcon Pointer_CT$wnnz_Int) : (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) > [(destructReadIn_CT$wnnz_Int,Word16#)] */
  assign destructReadIn_CT$wnnz_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                         scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon ReadIn_CT$wnnz_Int) : [(destructReadIn_CT$wnnz_Int,Word16#)] > (dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconReadIn_CT$wnnz_Int_d = ReadIn_CT$wnnz_Int_dc((& {destructReadIn_CT$wnnz_Int_d[0]}), destructReadIn_CT$wnnz_Int_d);
  assign {destructReadIn_CT$wnnz_Int_r} = {1 {(dconReadIn_CT$wnnz_Int_r && dconReadIn_CT$wnnz_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz_Int,
          Dcon ReadOut_CT$wnnz_Int) : (memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > [(readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int)] */
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_Int_d[116:2],
                                                       memReadOut_CT$wnnz_Int_d[0]};
  assign memReadOut_CT$wnnz_Int_r = readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wnnz_Int) : [(lizzieLet0_1_argbuf,CT$wnnz_Int),
                              (lizzieLet47_1_argbuf,CT$wnnz_Int),
                              (lizzieLet48_1_argbuf,CT$wnnz_Int),
                              (lizzieLet49_1_argbuf,CT$wnnz_Int),
                              (lizzieLet5_1_argbuf,CT$wnnz_Int)] > (writeMerge_choice_CT$wnnz_Int,C5) (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet47_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet48_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet49_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet5_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_Int_d[0],
                                                                      writeMerge_data_CT$wnnz_Int_d[0]} & {writeMerge_choice_CT$wnnz_Int_r,
                                                                                                           writeMerge_data_CT$wnnz_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet5_1_argbuf_r,
          lizzieLet49_1_argbuf_r,
          lizzieLet48_1_argbuf_r,
          lizzieLet47_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                          ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet47_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet48_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet49_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                              {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                            ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz_Int) : (writeMerge_choice_CT$wnnz_Int,C5) (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet47_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet48_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet49_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int)] */
  logic [4:0] demuxWriteResult_CT$wnnz_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_Int_d[0] && demuxWriteResult_CT$wnnz_Int_d[0]))
      unique case (writeMerge_choice_CT$wnnz_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[0]};
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[1]};
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[2]};
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[3]};
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_Int_r = (| (demuxWriteResult_CT$wnnz_Int_onehotd & {writeCT$wnnz_IntlizzieLet5_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet49_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet48_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet47_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_Int_r = demuxWriteResult_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon WriteIn_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In2,Word16#),
                                   (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int)] > (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconWriteIn_CT$wnnz_Int_d = WriteIn_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In2_d[0],
                                                                writeMerge_data_CT$wnnz_Int_d[0]}), forkHP1_CT$wnnz_In2_d, writeMerge_data_CT$wnnz_Int_d);
  assign {forkHP1_CT$wnnz_In2_r,
          writeMerge_data_CT$wnnz_Int_r} = {2 {(dconWriteIn_CT$wnnz_Int_r && dconWriteIn_CT$wnnz_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz_Int,
      Dcon Pointer_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In3,Word16#)] > (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) */
  assign dconPtr_CT$wnnz_Int_d = Pointer_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In3_d[0]}), forkHP1_CT$wnnz_In3_d);
  assign {forkHP1_CT$wnnz_In3_r} = {1 {(dconPtr_CT$wnnz_Int_r && dconPtr_CT$wnnz_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz_Int,
       Ty Pointer_CT$wnnz_Int) : (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(_171,Pointer_CT$wnnz_Int),
                                                                                                                           (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int)] */
  logic [1:0] dconPtr_CT$wnnz_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_Int_d[0] && dconPtr_CT$wnnz_Int_d[0]))
      unique case (memWriteOut_CT$wnnz_Int_d[1:1])
        1'd0: dconPtr_CT$wnnz_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_Int_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_Int_onehotd = 2'd0;
  assign _171_d = {dconPtr_CT$wnnz_Int_d[16:1],
                   dconPtr_CT$wnnz_Int_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_Int_d = {dconPtr_CT$wnnz_Int_d[16:1],
                                           dconPtr_CT$wnnz_Int_onehotd[1]};
  assign dconPtr_CT$wnnz_Int_r = (| (dconPtr_CT$wnnz_Int_onehotd & {demuxWriteResult_CT$wnnz_Int_r,
                                                                    _171_r}));
  assign memWriteOut_CT$wnnz_Int_r = dconPtr_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C6,
           Ty Pointer_QTree_Int) : [(m2ae4_1_argbuf,Pointer_QTree_Int),
                                    (m2aeH_1_argbuf,Pointer_QTree_Int),
                                    (m3ae5_1_argbuf,Pointer_QTree_Int),
                                    (m3aeI_1_argbuf,Pointer_QTree_Int),
                                    (q4'aex_1_argbuf,Pointer_QTree_Int),
                                    (wsjQ_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C6) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [5:0] m2ae4_1_argbuf_select_d;
  assign m2ae4_1_argbuf_select_d = ((| m2ae4_1_argbuf_select_q) ? m2ae4_1_argbuf_select_q :
                                    (m2ae4_1_argbuf_d[0] ? 6'd1 :
                                     (m2aeH_1_argbuf_d[0] ? 6'd2 :
                                      (m3ae5_1_argbuf_d[0] ? 6'd4 :
                                       (m3aeI_1_argbuf_d[0] ? 6'd8 :
                                        (\q4'aex_1_argbuf_d [0] ? 6'd16 :
                                         (wsjQ_1_1_argbuf_d[0] ? 6'd32 :
                                          6'd0)))))));
  logic [5:0] m2ae4_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae4_1_argbuf_select_q <= 6'd0;
    else
      m2ae4_1_argbuf_select_q <= (m2ae4_1_argbuf_done ? 6'd0 :
                                  m2ae4_1_argbuf_select_d);
  logic [1:0] m2ae4_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae4_1_argbuf_emit_q <= 2'd0;
    else
      m2ae4_1_argbuf_emit_q <= (m2ae4_1_argbuf_done ? 2'd0 :
                                m2ae4_1_argbuf_emit_d);
  logic [1:0] m2ae4_1_argbuf_emit_d;
  assign m2ae4_1_argbuf_emit_d = (m2ae4_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m2ae4_1_argbuf_done;
  assign m2ae4_1_argbuf_done = (& m2ae4_1_argbuf_emit_d);
  assign {wsjQ_1_1_argbuf_r,
          \q4'aex_1_argbuf_r ,
          m3aeI_1_argbuf_r,
          m3ae5_1_argbuf_r,
          m2aeH_1_argbuf_r,
          m2ae4_1_argbuf_r} = (m2ae4_1_argbuf_done ? m2ae4_1_argbuf_select_d :
                               6'd0);
  assign readMerge_data_QTree_Int_d = ((m2ae4_1_argbuf_select_d[0] && (! m2ae4_1_argbuf_emit_q[0])) ? m2ae4_1_argbuf_d :
                                       ((m2ae4_1_argbuf_select_d[1] && (! m2ae4_1_argbuf_emit_q[0])) ? m2aeH_1_argbuf_d :
                                        ((m2ae4_1_argbuf_select_d[2] && (! m2ae4_1_argbuf_emit_q[0])) ? m3ae5_1_argbuf_d :
                                         ((m2ae4_1_argbuf_select_d[3] && (! m2ae4_1_argbuf_emit_q[0])) ? m3aeI_1_argbuf_d :
                                          ((m2ae4_1_argbuf_select_d[4] && (! m2ae4_1_argbuf_emit_q[0])) ? \q4'aex_1_argbuf_d  :
                                           ((m2ae4_1_argbuf_select_d[5] && (! m2ae4_1_argbuf_emit_q[0])) ? wsjQ_1_1_argbuf_d :
                                            {16'd0, 1'd0}))))));
  assign readMerge_choice_QTree_Int_d = ((m2ae4_1_argbuf_select_d[0] && (! m2ae4_1_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                         ((m2ae4_1_argbuf_select_d[1] && (! m2ae4_1_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                          ((m2ae4_1_argbuf_select_d[2] && (! m2ae4_1_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                           ((m2ae4_1_argbuf_select_d[3] && (! m2ae4_1_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                            ((m2ae4_1_argbuf_select_d[4] && (! m2ae4_1_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                             ((m2ae4_1_argbuf_select_d[5] && (! m2ae4_1_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                              {3'd0, 1'd0}))))));
  
  /* demux (Ty C6,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C6) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm2ae4_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm2aeH_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm3ae5_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm3aeI_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intq4'aex_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntwsjQ_1_1_argbuf,QTree_Int)] */
  logic [5:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[3:1])
        3'd0: destructReadOut_QTree_Int_onehotd = 6'd1;
        3'd1: destructReadOut_QTree_Int_onehotd = 6'd2;
        3'd2: destructReadOut_QTree_Int_onehotd = 6'd4;
        3'd3: destructReadOut_QTree_Int_onehotd = 6'd8;
        3'd4: destructReadOut_QTree_Int_onehotd = 6'd16;
        3'd5: destructReadOut_QTree_Int_onehotd = 6'd32;
        default: destructReadOut_QTree_Int_onehotd = 6'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 6'd0;
  assign readPointer_QTree_Intm2ae4_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intm2aeH_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intm3ae5_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[2]};
  assign readPointer_QTree_Intm3aeI_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[3]};
  assign \readPointer_QTree_Intq4'aex_1_argbuf_d  = {destructReadOut_QTree_Int_d[66:1],
                                                     destructReadOut_QTree_Int_onehotd[4]};
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[5]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_IntwsjQ_1_1_argbuf_r,
                                                                                \readPointer_QTree_Intq4'aex_1_argbuf_r ,
                                                                                readPointer_QTree_Intm3aeI_1_argbuf_r,
                                                                                readPointer_QTree_Intm3ae5_1_argbuf_r,
                                                                                readPointer_QTree_Intm2aeH_1_argbuf_r,
                                                                                readPointer_QTree_Intm2ae4_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C29,
           Ty QTree_Int) : [(lizzieLet10_1_argbuf,QTree_Int),
                            (lizzieLet12_1_argbuf,QTree_Int),
                            (lizzieLet15_1_argbuf,QTree_Int),
                            (lizzieLet16_1_argbuf,QTree_Int),
                            (lizzieLet17_1_argbuf,QTree_Int),
                            (lizzieLet18_1_argbuf,QTree_Int),
                            (lizzieLet20_1_argbuf,QTree_Int),
                            (lizzieLet22_1_argbuf,QTree_Int),
                            (lizzieLet23_1_argbuf,QTree_Int),
                            (lizzieLet25_1_argbuf,QTree_Int),
                            (lizzieLet28_2_1_argbuf,QTree_Int),
                            (lizzieLet29_1_1_argbuf,QTree_Int),
                            (lizzieLet30_1_1_argbuf,QTree_Int),
                            (lizzieLet31_1_argbuf,QTree_Int),
                            (lizzieLet33_1_1_argbuf,QTree_Int),
                            (lizzieLet33_1_argbuf,QTree_Int),
                            (lizzieLet34_1_argbuf,QTree_Int),
                            (lizzieLet35_1_argbuf,QTree_Int),
                            (lizzieLet36_1_argbuf,QTree_Int),
                            (lizzieLet38_1_argbuf,QTree_Int),
                            (lizzieLet39_1_argbuf,QTree_Int),
                            (lizzieLet41_1_argbuf,QTree_Int),
                            (lizzieLet42_1_argbuf,QTree_Int),
                            (lizzieLet54_1_argbuf,QTree_Int),
                            (lizzieLet59_1_argbuf,QTree_Int),
                            (lizzieLet64_1_argbuf,QTree_Int),
                            (lizzieLet7_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C29) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [28:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 29'd1 :
                                           (lizzieLet12_1_argbuf_d[0] ? 29'd2 :
                                            (lizzieLet15_1_argbuf_d[0] ? 29'd4 :
                                             (lizzieLet16_1_argbuf_d[0] ? 29'd8 :
                                              (lizzieLet17_1_argbuf_d[0] ? 29'd16 :
                                               (lizzieLet18_1_argbuf_d[0] ? 29'd32 :
                                                (lizzieLet20_1_argbuf_d[0] ? 29'd64 :
                                                 (lizzieLet22_1_argbuf_d[0] ? 29'd128 :
                                                  (lizzieLet23_1_argbuf_d[0] ? 29'd256 :
                                                   (lizzieLet25_1_argbuf_d[0] ? 29'd512 :
                                                    (lizzieLet28_2_1_argbuf_d[0] ? 29'd1024 :
                                                     (lizzieLet29_1_1_argbuf_d[0] ? 29'd2048 :
                                                      (lizzieLet30_1_1_argbuf_d[0] ? 29'd4096 :
                                                       (lizzieLet31_1_argbuf_d[0] ? 29'd8192 :
                                                        (lizzieLet33_1_1_argbuf_d[0] ? 29'd16384 :
                                                         (lizzieLet33_1_argbuf_d[0] ? 29'd32768 :
                                                          (lizzieLet34_1_argbuf_d[0] ? 29'd65536 :
                                                           (lizzieLet35_1_argbuf_d[0] ? 29'd131072 :
                                                            (lizzieLet36_1_argbuf_d[0] ? 29'd262144 :
                                                             (lizzieLet38_1_argbuf_d[0] ? 29'd524288 :
                                                              (lizzieLet39_1_argbuf_d[0] ? 29'd1048576 :
                                                               (lizzieLet41_1_argbuf_d[0] ? 29'd2097152 :
                                                                (lizzieLet42_1_argbuf_d[0] ? 29'd4194304 :
                                                                 (lizzieLet54_1_argbuf_d[0] ? 29'd8388608 :
                                                                  (lizzieLet59_1_argbuf_d[0] ? 29'd16777216 :
                                                                   (lizzieLet64_1_argbuf_d[0] ? 29'd33554432 :
                                                                    (lizzieLet7_1_argbuf_d[0] ? 29'd67108864 :
                                                                     (lizzieLet9_1_argbuf_d[0] ? 29'd134217728 :
                                                                      (dummy_write_QTree_Int_d[0] ? 29'd268435456 :
                                                                       29'd0))))))))))))))))))))))))))))));
  logic [28:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 29'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 29'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                        writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                           writeMerge_data_QTree_Int_r}));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet64_1_argbuf_r,
          lizzieLet59_1_argbuf_r,
          lizzieLet54_1_argbuf_r,
          lizzieLet42_1_argbuf_r,
          lizzieLet41_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet33_1_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_1_argbuf_r,
          lizzieLet29_1_1_argbuf_r,
          lizzieLet28_2_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     29'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                        ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet12_1_argbuf_d :
                                         ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                          ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                           ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                            ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                             ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                              ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                               ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                 ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet28_2_1_argbuf_d :
                                                  ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet29_1_1_argbuf_d :
                                                   ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet30_1_1_argbuf_d :
                                                    ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                     ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet33_1_1_argbuf_d :
                                                      ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                                       ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                        ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                         ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                          ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                                           ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                                            ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet41_1_argbuf_d :
                                                             ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet42_1_argbuf_d :
                                                              ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet54_1_argbuf_d :
                                                               ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet59_1_argbuf_d :
                                                                ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet64_1_argbuf_d :
                                                                 ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                                                  ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                                   ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                                    {66'd0,
                                                                     1'd0})))))))))))))))))))))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_29_dc(1'd1) :
                                          ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_29_dc(1'd1) :
                                           ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_29_dc(1'd1) :
                                            ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_29_dc(1'd1) :
                                             ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_29_dc(1'd1) :
                                              ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C6_29_dc(1'd1) :
                                               ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C7_29_dc(1'd1) :
                                                ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C8_29_dc(1'd1) :
                                                 ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C9_29_dc(1'd1) :
                                                  ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C10_29_dc(1'd1) :
                                                   ((lizzieLet10_1_argbuf_select_d[10] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C11_29_dc(1'd1) :
                                                    ((lizzieLet10_1_argbuf_select_d[11] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C12_29_dc(1'd1) :
                                                     ((lizzieLet10_1_argbuf_select_d[12] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C13_29_dc(1'd1) :
                                                      ((lizzieLet10_1_argbuf_select_d[13] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C14_29_dc(1'd1) :
                                                       ((lizzieLet10_1_argbuf_select_d[14] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C15_29_dc(1'd1) :
                                                        ((lizzieLet10_1_argbuf_select_d[15] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C16_29_dc(1'd1) :
                                                         ((lizzieLet10_1_argbuf_select_d[16] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C17_29_dc(1'd1) :
                                                          ((lizzieLet10_1_argbuf_select_d[17] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C18_29_dc(1'd1) :
                                                           ((lizzieLet10_1_argbuf_select_d[18] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C19_29_dc(1'd1) :
                                                            ((lizzieLet10_1_argbuf_select_d[19] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C20_29_dc(1'd1) :
                                                             ((lizzieLet10_1_argbuf_select_d[20] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C21_29_dc(1'd1) :
                                                              ((lizzieLet10_1_argbuf_select_d[21] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C22_29_dc(1'd1) :
                                                               ((lizzieLet10_1_argbuf_select_d[22] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C23_29_dc(1'd1) :
                                                                ((lizzieLet10_1_argbuf_select_d[23] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C24_29_dc(1'd1) :
                                                                 ((lizzieLet10_1_argbuf_select_d[24] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C25_29_dc(1'd1) :
                                                                  ((lizzieLet10_1_argbuf_select_d[25] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C26_29_dc(1'd1) :
                                                                   ((lizzieLet10_1_argbuf_select_d[26] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C27_29_dc(1'd1) :
                                                                    ((lizzieLet10_1_argbuf_select_d[27] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C28_29_dc(1'd1) :
                                                                     ((lizzieLet10_1_argbuf_select_d[28] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C29_29_dc(1'd1) :
                                                                      {5'd0,
                                                                       1'd0})))))))))))))))))))))))))))));
  
  /* demux (Ty C29,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C29) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet12_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet23_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet25_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet28_2_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet29_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet30_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet33_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet35_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet36_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet38_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet39_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet41_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet42_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet54_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet59_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet64_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [28:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[5:1])
        5'd0: demuxWriteResult_QTree_Int_onehotd = 29'd1;
        5'd1: demuxWriteResult_QTree_Int_onehotd = 29'd2;
        5'd2: demuxWriteResult_QTree_Int_onehotd = 29'd4;
        5'd3: demuxWriteResult_QTree_Int_onehotd = 29'd8;
        5'd4: demuxWriteResult_QTree_Int_onehotd = 29'd16;
        5'd5: demuxWriteResult_QTree_Int_onehotd = 29'd32;
        5'd6: demuxWriteResult_QTree_Int_onehotd = 29'd64;
        5'd7: demuxWriteResult_QTree_Int_onehotd = 29'd128;
        5'd8: demuxWriteResult_QTree_Int_onehotd = 29'd256;
        5'd9: demuxWriteResult_QTree_Int_onehotd = 29'd512;
        5'd10: demuxWriteResult_QTree_Int_onehotd = 29'd1024;
        5'd11: demuxWriteResult_QTree_Int_onehotd = 29'd2048;
        5'd12: demuxWriteResult_QTree_Int_onehotd = 29'd4096;
        5'd13: demuxWriteResult_QTree_Int_onehotd = 29'd8192;
        5'd14: demuxWriteResult_QTree_Int_onehotd = 29'd16384;
        5'd15: demuxWriteResult_QTree_Int_onehotd = 29'd32768;
        5'd16: demuxWriteResult_QTree_Int_onehotd = 29'd65536;
        5'd17: demuxWriteResult_QTree_Int_onehotd = 29'd131072;
        5'd18: demuxWriteResult_QTree_Int_onehotd = 29'd262144;
        5'd19: demuxWriteResult_QTree_Int_onehotd = 29'd524288;
        5'd20: demuxWriteResult_QTree_Int_onehotd = 29'd1048576;
        5'd21: demuxWriteResult_QTree_Int_onehotd = 29'd2097152;
        5'd22: demuxWriteResult_QTree_Int_onehotd = 29'd4194304;
        5'd23: demuxWriteResult_QTree_Int_onehotd = 29'd8388608;
        5'd24: demuxWriteResult_QTree_Int_onehotd = 29'd16777216;
        5'd25: demuxWriteResult_QTree_Int_onehotd = 29'd33554432;
        5'd26: demuxWriteResult_QTree_Int_onehotd = 29'd67108864;
        5'd27: demuxWriteResult_QTree_Int_onehotd = 29'd134217728;
        5'd28: demuxWriteResult_QTree_Int_onehotd = 29'd268435456;
        default: demuxWriteResult_QTree_Int_onehotd = 29'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 29'd0;
  assign writeQTree_IntlizzieLet10_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet12_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet16_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet17_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet23_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[8]};
  assign writeQTree_IntlizzieLet25_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[9]};
  assign writeQTree_IntlizzieLet28_2_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[10]};
  assign writeQTree_IntlizzieLet29_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[11]};
  assign writeQTree_IntlizzieLet30_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[12]};
  assign writeQTree_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[13]};
  assign writeQTree_IntlizzieLet33_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[14]};
  assign writeQTree_IntlizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[15]};
  assign writeQTree_IntlizzieLet34_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[16]};
  assign writeQTree_IntlizzieLet35_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[17]};
  assign writeQTree_IntlizzieLet36_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[18]};
  assign writeQTree_IntlizzieLet38_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[19]};
  assign writeQTree_IntlizzieLet39_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[20]};
  assign writeQTree_IntlizzieLet41_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[21]};
  assign writeQTree_IntlizzieLet42_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[22]};
  assign writeQTree_IntlizzieLet54_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[23]};
  assign writeQTree_IntlizzieLet59_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[24]};
  assign writeQTree_IntlizzieLet64_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[25]};
  assign writeQTree_IntlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[26]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[27]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[28]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet64_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet59_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet54_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet42_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet41_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet39_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet38_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet36_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet35_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet34_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet33_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet33_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet31_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet30_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet29_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet28_2_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet25_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet23_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet22_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet20_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet18_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet17_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet16_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet15_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet12_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet10_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_170,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _170_d = {dconPtr_QTree_Int_d[16:1],
                   dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _170_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__7,Go) > (initHP_CTf'''''''''_f'''''''''_Int,Word16#) */
  assign \initHP_CTf'''''''''_f'''''''''_Int_d  = {16'd0,
                                                   go__7_d[0]};
  assign go__7_r = \initHP_CTf'''''''''_f'''''''''_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf'''''''''_f'''''''''_Int1,Go) > (incrHP_CTf'''''''''_f'''''''''_Int,Word16#) */
  assign \incrHP_CTf'''''''''_f'''''''''_Int_d  = {16'd1,
                                                   \incrHP_CTf'''''''''_f'''''''''_Int1_d [0]};
  assign \incrHP_CTf'''''''''_f'''''''''_Int1_r  = \incrHP_CTf'''''''''_f'''''''''_Int_r ;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CTf'''''''''_f'''''''''_Int2,Go)] > (incrHP_mergeCTf'''''''''_f'''''''''_Int,Go) */
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected ;
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTf'''''''''_f'''''''''_Int_select ))
        \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected  = \incrHP_mergeCTf'''''''''_f'''''''''_Int_select ;
      else
        if (go__8_d[0])
          \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected [0] = 1'd1;
        else if (\incrHP_CTf'''''''''_f'''''''''_Int2_d [0])
          \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_select  <= (\incrHP_mergeCTf'''''''''_f'''''''''_Int_r  ? 2'd0 :
                                                           \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected );
  always_comb
    if (\incrHP_mergeCTf'''''''''_f'''''''''_Int_selected [0])
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_d  = go__8_d;
    else if (\incrHP_mergeCTf'''''''''_f'''''''''_Int_selected [1])
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_d  = \incrHP_CTf'''''''''_f'''''''''_Int2_d ;
    else \incrHP_mergeCTf'''''''''_f'''''''''_Int_d  = 1'd0;
  assign {\incrHP_CTf'''''''''_f'''''''''_Int2_r ,
          go__8_r} = (\incrHP_mergeCTf'''''''''_f'''''''''_Int_r  ? \incrHP_mergeCTf'''''''''_f'''''''''_Int_selected  :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf'''''''''_f'''''''''_Int_buf,Go) > [(incrHP_CTf'''''''''_f'''''''''_Int1,Go),
                                                                   (incrHP_CTf'''''''''_f'''''''''_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_done ;
  assign \incrHP_CTf'''''''''_f'''''''''_Int1_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_d [0] && (! \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted [0]));
  assign \incrHP_CTf'''''''''_f'''''''''_Int2_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_d [0] && (! \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted [1]));
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_done  = (\incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted  | ({\incrHP_CTf'''''''''_f'''''''''_Int2_d [0],
                                                                                                                         \incrHP_CTf'''''''''_f'''''''''_Int1_d [0]} & {\incrHP_CTf'''''''''_f'''''''''_Int2_r ,
                                                                                                                                                                        \incrHP_CTf'''''''''_f'''''''''_Int1_r }));
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_r  = (& \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_emitted  <= (\incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_r  ? 2'd0 :
                                                                \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf'''''''''_f'''''''''_Int,Word16#) (forkHP1_CTf'''''''''_f'''''''''_Int,Word16#) > (addHP_CTf'''''''''_f'''''''''_Int,Word16#) */
  assign \addHP_CTf'''''''''_f'''''''''_Int_d  = {(\incrHP_CTf'''''''''_f'''''''''_Int_d [16:1] + \forkHP1_CTf'''''''''_f'''''''''_Int_d [16:1]),
                                                  (\incrHP_CTf'''''''''_f'''''''''_Int_d [0] && \forkHP1_CTf'''''''''_f'''''''''_Int_d [0])};
  assign {\incrHP_CTf'''''''''_f'''''''''_Int_r ,
          \forkHP1_CTf'''''''''_f'''''''''_Int_r } = {2 {(\addHP_CTf'''''''''_f'''''''''_Int_r  && \addHP_CTf'''''''''_f'''''''''_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf'''''''''_f'''''''''_Int,Word16#),
                      (addHP_CTf'''''''''_f'''''''''_Int,Word16#)] > (mergeHP_CTf'''''''''_f'''''''''_Int,Word16#) */
  logic [1:0] \mergeHP_CTf'''''''''_f'''''''''_Int_selected ;
  logic [1:0] \mergeHP_CTf'''''''''_f'''''''''_Int_select ;
  always_comb
    begin
      \mergeHP_CTf'''''''''_f'''''''''_Int_selected  = 2'd0;
      if ((| \mergeHP_CTf'''''''''_f'''''''''_Int_select ))
        \mergeHP_CTf'''''''''_f'''''''''_Int_selected  = \mergeHP_CTf'''''''''_f'''''''''_Int_select ;
      else
        if (\initHP_CTf'''''''''_f'''''''''_Int_d [0])
          \mergeHP_CTf'''''''''_f'''''''''_Int_selected [0] = 1'd1;
        else if (\addHP_CTf'''''''''_f'''''''''_Int_d [0])
          \mergeHP_CTf'''''''''_f'''''''''_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Int_select  <= 2'd0;
    else
      \mergeHP_CTf'''''''''_f'''''''''_Int_select  <= (\mergeHP_CTf'''''''''_f'''''''''_Int_r  ? 2'd0 :
                                                       \mergeHP_CTf'''''''''_f'''''''''_Int_selected );
  always_comb
    if (\mergeHP_CTf'''''''''_f'''''''''_Int_selected [0])
      \mergeHP_CTf'''''''''_f'''''''''_Int_d  = \initHP_CTf'''''''''_f'''''''''_Int_d ;
    else if (\mergeHP_CTf'''''''''_f'''''''''_Int_selected [1])
      \mergeHP_CTf'''''''''_f'''''''''_Int_d  = \addHP_CTf'''''''''_f'''''''''_Int_d ;
    else \mergeHP_CTf'''''''''_f'''''''''_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTf'''''''''_f'''''''''_Int_r ,
          \initHP_CTf'''''''''_f'''''''''_Int_r } = (\mergeHP_CTf'''''''''_f'''''''''_Int_r  ? \mergeHP_CTf'''''''''_f'''''''''_Int_selected  :
                                                     2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf'''''''''_f'''''''''_Int,Go) > (incrHP_mergeCTf'''''''''_f'''''''''_Int_buf,Go) */
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d ;
  logic \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_r ;
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Int_r  = ((! \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d [0]) || \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf'''''''''_f'''''''''_Int_r )
        \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d  <= \incrHP_mergeCTf'''''''''_f'''''''''_Int_d ;
  Go_t \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf ;
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_r  = (! \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_d  = (\incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf [0] ? \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf  :
                                                            \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_r  && \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf [0]))
        \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf'''''''''_f'''''''''_Int_buf_r ) && (! \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf [0])))
        \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_buf  <= \incrHP_mergeCTf'''''''''_f'''''''''_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf'''''''''_f'''''''''_Int,Word16#) > (mergeHP_CTf'''''''''_f'''''''''_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d ;
  logic \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_r ;
  assign \mergeHP_CTf'''''''''_f'''''''''_Int_r  = ((! \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d [0]) || \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf'''''''''_f'''''''''_Int_r )
        \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d  <= \mergeHP_CTf'''''''''_f'''''''''_Int_d ;
  \Word16#_t  \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf ;
  assign \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_r  = (! \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf [0]);
  assign \mergeHP_CTf'''''''''_f'''''''''_Int_buf_d  = (\mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf [0] ? \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf  :
                                                        \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf'''''''''_f'''''''''_Int_buf_r  && \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf [0]))
        \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf'''''''''_f'''''''''_Int_buf_r ) && (! \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf [0])))
        \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_buf  <= \mergeHP_CTf'''''''''_f'''''''''_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf'''''''''_f'''''''''_Int_buf,Word16#) > [(forkHP1_CTf'''''''''_f'''''''''_Int,Word16#),
                                                                         (forkHP1_CTf'''''''''_f'''''''''_In2,Word16#),
                                                                         (forkHP1_CTf'''''''''_f'''''''''_In3,Word16#)] */
  logic [2:0] \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTf'''''''''_f'''''''''_Int_buf_done ;
  assign \forkHP1_CTf'''''''''_f'''''''''_Int_d  = {\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [16:1],
                                                    (\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted [0]))};
  assign \forkHP1_CTf'''''''''_f'''''''''_In2_d  = {\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [16:1],
                                                    (\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted [1]))};
  assign \forkHP1_CTf'''''''''_f'''''''''_In3_d  = {\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [16:1],
                                                    (\mergeHP_CTf'''''''''_f'''''''''_Int_buf_d [0] && (! \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted [2]))};
  assign \mergeHP_CTf'''''''''_f'''''''''_Int_buf_done  = (\mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted  | ({\forkHP1_CTf'''''''''_f'''''''''_In3_d [0],
                                                                                                                 \forkHP1_CTf'''''''''_f'''''''''_In2_d [0],
                                                                                                                 \forkHP1_CTf'''''''''_f'''''''''_Int_d [0]} & {\forkHP1_CTf'''''''''_f'''''''''_In3_r ,
                                                                                                                                                                \forkHP1_CTf'''''''''_f'''''''''_In2_r ,
                                                                                                                                                                \forkHP1_CTf'''''''''_f'''''''''_Int_r }));
  assign \mergeHP_CTf'''''''''_f'''''''''_Int_buf_r  = (& \mergeHP_CTf'''''''''_f'''''''''_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf'''''''''_f'''''''''_Int_buf_emitted  <= (\mergeHP_CTf'''''''''_f'''''''''_Int_buf_r  ? 3'd0 :
                                                            \mergeHP_CTf'''''''''_f'''''''''_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf'''''''''_f'''''''''_Int) : [(dconReadIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int),
                                                    (dconWriteIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int)] > (memMergeChoice_CTf'''''''''_f'''''''''_Int,C2) (memMergeIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int) */
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Int_select_d ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Int_select_d  = ((| \dconReadIn_CTf'''''''''_f'''''''''_Int_select_q ) ? \dconReadIn_CTf'''''''''_f'''''''''_Int_select_q  :
                                                              (\dconReadIn_CTf'''''''''_f'''''''''_Int_d [0] ? 2'd1 :
                                                               (\dconWriteIn_CTf'''''''''_f'''''''''_Int_d [0] ? 2'd2 :
                                                                2'd0)));
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'''''''''_f'''''''''_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTf'''''''''_f'''''''''_Int_select_q  <= (\dconReadIn_CTf'''''''''_f'''''''''_Int_done  ? 2'd0 :
                                                            \dconReadIn_CTf'''''''''_f'''''''''_Int_select_d );
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q  <= (\dconReadIn_CTf'''''''''_f'''''''''_Int_done  ? 2'd0 :
                                                          \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_d );
  logic [1:0] \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_d ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_d  = (\dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q  | ({\memMergeChoice_CTf'''''''''_f'''''''''_Int_d [0],
                                                                                                                \memMergeIn_CTf'''''''''_f'''''''''_Int_d [0]} & {\memMergeChoice_CTf'''''''''_f'''''''''_Int_r ,
                                                                                                                                                                  \memMergeIn_CTf'''''''''_f'''''''''_Int_r }));
  logic \dconReadIn_CTf'''''''''_f'''''''''_Int_done ;
  assign \dconReadIn_CTf'''''''''_f'''''''''_Int_done  = (& \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_d );
  assign {\dconWriteIn_CTf'''''''''_f'''''''''_Int_r ,
          \dconReadIn_CTf'''''''''_f'''''''''_Int_r } = (\dconReadIn_CTf'''''''''_f'''''''''_Int_done  ? \dconReadIn_CTf'''''''''_f'''''''''_Int_select_d  :
                                                         2'd0);
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_d  = ((\dconReadIn_CTf'''''''''_f'''''''''_Int_select_d [0] && (! \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q [0])) ? \dconReadIn_CTf'''''''''_f'''''''''_Int_d  :
                                                       ((\dconReadIn_CTf'''''''''_f'''''''''_Int_select_d [1] && (! \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q [0])) ? \dconWriteIn_CTf'''''''''_f'''''''''_Int_d  :
                                                        {132'd0, 1'd0}));
  assign \memMergeChoice_CTf'''''''''_f'''''''''_Int_d  = ((\dconReadIn_CTf'''''''''_f'''''''''_Int_select_d [0] && (! \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                           ((\dconReadIn_CTf'''''''''_f'''''''''_Int_select_d [1] && (! \dconReadIn_CTf'''''''''_f'''''''''_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                            {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf'''''''''_f'''''''''_Int,
      Ty MemOut_CTf'''''''''_f'''''''''_Int) : (memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf,MemIn_CTf'''''''''_f'''''''''_Int) > (memOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int) */
  logic [114:0] \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_address ;
  logic [114:0] \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_din ;
  logic [114:0] \memOut_CTf'''''''''_f'''''''''_Int_q ;
  logic \memOut_CTf'''''''''_f'''''''''_Int_valid ;
  logic \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_we ;
  logic \memOut_CTf'''''''''_f'''''''''_Int_we ;
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_din  = \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [132:18];
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_address  = \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [17:2];
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_we  = (\memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [1:1] && \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf'''''''''_f'''''''''_Int_we  <= 1'd0;
        \memOut_CTf'''''''''_f'''''''''_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf'''''''''_f'''''''''_Int_we  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_we ;
        \memOut_CTf'''''''''_f'''''''''_Int_valid  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [0];
        if (\memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_we )
          begin
            \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_mem [\memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_address ] <= \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_din ;
            \memOut_CTf'''''''''_f'''''''''_Int_q  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_din ;
          end
        else
          \memOut_CTf'''''''''_f'''''''''_Int_q  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_mem [\memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_address ];
      end
  assign \memOut_CTf'''''''''_f'''''''''_Int_d  = {\memOut_CTf'''''''''_f'''''''''_Int_q ,
                                                   \memOut_CTf'''''''''_f'''''''''_Int_we ,
                                                   \memOut_CTf'''''''''_f'''''''''_Int_valid };
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_r  = ((! \memOut_CTf'''''''''_f'''''''''_Int_valid ) || \memOut_CTf'''''''''_f'''''''''_Int_r );
  
  /* demux (Ty C2,
       Ty MemOut_CTf'''''''''_f'''''''''_Int) : (memMergeChoice_CTf'''''''''_f'''''''''_Int,C2) (memOut_CTf'''''''''_f'''''''''_Int_dbuf,MemOut_CTf'''''''''_f'''''''''_Int) > [(memReadOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                (memWriteOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int)] */
  logic [1:0] \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf'''''''''_f'''''''''_Int_d [0] && \memOut_CTf'''''''''_f'''''''''_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTf'''''''''_f'''''''''_Int_d [1:1])
        1'd0: \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf'''''''''_f'''''''''_Int_d  = {\memOut_CTf'''''''''_f'''''''''_Int_dbuf_d [116:1],
                                                       \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTf'''''''''_f'''''''''_Int_d  = {\memOut_CTf'''''''''_f'''''''''_Int_dbuf_d [116:1],
                                                        \memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd [1]};
  assign \memOut_CTf'''''''''_f'''''''''_Int_dbuf_r  = (| (\memOut_CTf'''''''''_f'''''''''_Int_dbuf_onehotd  & {\memWriteOut_CTf'''''''''_f'''''''''_Int_r ,
                                                                                                                \memReadOut_CTf'''''''''_f'''''''''_Int_r }));
  assign \memMergeChoice_CTf'''''''''_f'''''''''_Int_r  = \memOut_CTf'''''''''_f'''''''''_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf'''''''''_f'''''''''_Int) : (memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf,MemIn_CTf'''''''''_f'''''''''_Int) > (memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf,MemIn_CTf'''''''''_f'''''''''_Int) */
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_r  = ((! \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d [0]) || \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d  <= {132'd0, 1'd0};
    else
      if (\memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_r )
        \memMergeIn_CTf'''''''''_f'''''''''_Int_dbuf_d  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf'''''''''_f'''''''''_Int) : (memMergeIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int) > (memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf,MemIn_CTf'''''''''_f'''''''''_Int) */
  \MemIn_CTf'''''''''_f'''''''''_Int_t  \memMergeIn_CTf'''''''''_f'''''''''_Int_buf ;
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_r  = (! \memMergeIn_CTf'''''''''_f'''''''''_Int_buf [0]);
  assign \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_d  = (\memMergeIn_CTf'''''''''_f'''''''''_Int_buf [0] ? \memMergeIn_CTf'''''''''_f'''''''''_Int_buf  :
                                                            \memMergeIn_CTf'''''''''_f'''''''''_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'''''''''_f'''''''''_Int_buf  <= {132'd0, 1'd0};
    else
      if ((\memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_r  && \memMergeIn_CTf'''''''''_f'''''''''_Int_buf [0]))
        \memMergeIn_CTf'''''''''_f'''''''''_Int_buf  <= {132'd0, 1'd0};
      else if (((! \memMergeIn_CTf'''''''''_f'''''''''_Int_rbuf_r ) && (! \memMergeIn_CTf'''''''''_f'''''''''_Int_buf [0])))
        \memMergeIn_CTf'''''''''_f'''''''''_Int_buf  <= \memMergeIn_CTf'''''''''_f'''''''''_Int_d ;
  
  /* dbuf (Ty MemOut_CTf'''''''''_f'''''''''_Int) : (memOut_CTf'''''''''_f'''''''''_Int_rbuf,MemOut_CTf'''''''''_f'''''''''_Int) > (memOut_CTf'''''''''_f'''''''''_Int_dbuf,MemOut_CTf'''''''''_f'''''''''_Int) */
  assign \memOut_CTf'''''''''_f'''''''''_Int_rbuf_r  = ((! \memOut_CTf'''''''''_f'''''''''_Int_dbuf_d [0]) || \memOut_CTf'''''''''_f'''''''''_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'''''''''_f'''''''''_Int_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memOut_CTf'''''''''_f'''''''''_Int_rbuf_r )
        \memOut_CTf'''''''''_f'''''''''_Int_dbuf_d  <= \memOut_CTf'''''''''_f'''''''''_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf'''''''''_f'''''''''_Int) : (memOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int) > (memOut_CTf'''''''''_f'''''''''_Int_rbuf,MemOut_CTf'''''''''_f'''''''''_Int) */
  \MemOut_CTf'''''''''_f'''''''''_Int_t  \memOut_CTf'''''''''_f'''''''''_Int_buf ;
  assign \memOut_CTf'''''''''_f'''''''''_Int_r  = (! \memOut_CTf'''''''''_f'''''''''_Int_buf [0]);
  assign \memOut_CTf'''''''''_f'''''''''_Int_rbuf_d  = (\memOut_CTf'''''''''_f'''''''''_Int_buf [0] ? \memOut_CTf'''''''''_f'''''''''_Int_buf  :
                                                        \memOut_CTf'''''''''_f'''''''''_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'''''''''_f'''''''''_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf'''''''''_f'''''''''_Int_rbuf_r  && \memOut_CTf'''''''''_f'''''''''_Int_buf [0]))
        \memOut_CTf'''''''''_f'''''''''_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf'''''''''_f'''''''''_Int_rbuf_r ) && (! \memOut_CTf'''''''''_f'''''''''_Int_buf [0])))
        \memOut_CTf'''''''''_f'''''''''_Int_buf  <= \memOut_CTf'''''''''_f'''''''''_Int_d ;
  
  /* destruct (Ty Pointer_CTf'''''''''_f'''''''''_Int,
          Dcon Pointer_CTf'''''''''_f'''''''''_Int) : (scfarg_0_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > [(destructReadIn_CTf'''''''''_f'''''''''_Int,Word16#)] */
  assign \destructReadIn_CTf'''''''''_f'''''''''_Int_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                           scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf'''''''''_f'''''''''_Int_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''_f'''''''''_Int,
      Dcon ReadIn_CTf'''''''''_f'''''''''_Int) : [(destructReadIn_CTf'''''''''_f'''''''''_Int,Word16#)] > (dconReadIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int) */
  assign \dconReadIn_CTf'''''''''_f'''''''''_Int_d  = \ReadIn_CTf'''''''''_f'''''''''_Int_dc ((& {\destructReadIn_CTf'''''''''_f'''''''''_Int_d [0]}), \destructReadIn_CTf'''''''''_f'''''''''_Int_d );
  assign {\destructReadIn_CTf'''''''''_f'''''''''_Int_r } = {1 {(\dconReadIn_CTf'''''''''_f'''''''''_Int_r  && \dconReadIn_CTf'''''''''_f'''''''''_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTf'''''''''_f'''''''''_Int,
          Dcon ReadOut_CTf'''''''''_f'''''''''_Int) : (memReadOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int) > [(readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf,CTf'''''''''_f'''''''''_Int)] */
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_d  = {\memReadOut_CTf'''''''''_f'''''''''_Int_d [116:2],
                                                                           \memReadOut_CTf'''''''''_f'''''''''_Int_d [0]};
  assign \memReadOut_CTf'''''''''_f'''''''''_Int_r  = \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf'''''''''_f'''''''''_Int) : [(lizzieLet11_1_argbuf,CTf'''''''''_f'''''''''_Int),
                                              (lizzieLet43_1_argbuf,CTf'''''''''_f'''''''''_Int),
                                              (lizzieLet51_1_argbuf,CTf'''''''''_f'''''''''_Int),
                                              (lizzieLet52_1_argbuf,CTf'''''''''_f'''''''''_Int),
                                              (lizzieLet53_1_argbuf,CTf'''''''''_f'''''''''_Int)] > (writeMerge_choice_CTf'''''''''_f'''''''''_Int,C5) (writeMerge_data_CTf'''''''''_f'''''''''_Int,CTf'''''''''_f'''''''''_Int) */
  logic [4:0] lizzieLet11_1_argbuf_select_d;
  assign lizzieLet11_1_argbuf_select_d = ((| lizzieLet11_1_argbuf_select_q) ? lizzieLet11_1_argbuf_select_q :
                                          (lizzieLet11_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet43_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet51_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet52_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet53_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet11_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet11_1_argbuf_select_q <= (lizzieLet11_1_argbuf_done ? 5'd0 :
                                        lizzieLet11_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_argbuf_emit_q <= (lizzieLet11_1_argbuf_done ? 2'd0 :
                                      lizzieLet11_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_argbuf_emit_d;
  assign lizzieLet11_1_argbuf_emit_d = (lizzieLet11_1_argbuf_emit_q | ({\writeMerge_choice_CTf'''''''''_f'''''''''_Int_d [0],
                                                                        \writeMerge_data_CTf'''''''''_f'''''''''_Int_d [0]} & {\writeMerge_choice_CTf'''''''''_f'''''''''_Int_r ,
                                                                                                                               \writeMerge_data_CTf'''''''''_f'''''''''_Int_r }));
  logic lizzieLet11_1_argbuf_done;
  assign lizzieLet11_1_argbuf_done = (& lizzieLet11_1_argbuf_emit_d);
  assign {lizzieLet53_1_argbuf_r,
          lizzieLet52_1_argbuf_r,
          lizzieLet51_1_argbuf_r,
          lizzieLet43_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (lizzieLet11_1_argbuf_done ? lizzieLet11_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf'''''''''_f'''''''''_Int_d  = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet11_1_argbuf_d :
                                                            ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet43_1_argbuf_d :
                                                             ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet51_1_argbuf_d :
                                                              ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet52_1_argbuf_d :
                                                               ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[0])) ? lizzieLet53_1_argbuf_d :
                                                                {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf'''''''''_f'''''''''_Int_d  = ((lizzieLet11_1_argbuf_select_d[0] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                              ((lizzieLet11_1_argbuf_select_d[1] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                               ((lizzieLet11_1_argbuf_select_d[2] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                ((lizzieLet11_1_argbuf_select_d[3] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                 ((lizzieLet11_1_argbuf_select_d[4] && (! lizzieLet11_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                  {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeMerge_choice_CTf'''''''''_f'''''''''_Int,C5) (demuxWriteResult_CTf'''''''''_f'''''''''_Int,Pointer_CTf'''''''''_f'''''''''_Int) > [(writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                          (writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                          (writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                          (writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                          (writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [4:0] \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf'''''''''_f'''''''''_Int_d [0] && \demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [0]))
      unique case (\writeMerge_choice_CTf'''''''''_f'''''''''_Int_d [3:1])
        3'd0:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  = 5'd0;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                                     \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd [0]};
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                                     \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd [1]};
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                                     \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd [2]};
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                                     \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd [3]};
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_d  = {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                                     \demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd [4]};
  assign \demuxWriteResult_CTf'''''''''_f'''''''''_Int_r  = (| (\demuxWriteResult_CTf'''''''''_f'''''''''_Int_onehotd  & {\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_r ,
                                                                                                                          \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_r ,
                                                                                                                          \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_r ,
                                                                                                                          \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_r ,
                                                                                                                          \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_r }));
  assign \writeMerge_choice_CTf'''''''''_f'''''''''_Int_r  = \demuxWriteResult_CTf'''''''''_f'''''''''_Int_r ;
  
  /* dcon (Ty MemIn_CTf'''''''''_f'''''''''_Int,
      Dcon WriteIn_CTf'''''''''_f'''''''''_Int) : [(forkHP1_CTf'''''''''_f'''''''''_In2,Word16#),
                                                   (writeMerge_data_CTf'''''''''_f'''''''''_Int,CTf'''''''''_f'''''''''_Int)] > (dconWriteIn_CTf'''''''''_f'''''''''_Int,MemIn_CTf'''''''''_f'''''''''_Int) */
  assign \dconWriteIn_CTf'''''''''_f'''''''''_Int_d  = \WriteIn_CTf'''''''''_f'''''''''_Int_dc ((& {\forkHP1_CTf'''''''''_f'''''''''_In2_d [0],
                                                                                                    \writeMerge_data_CTf'''''''''_f'''''''''_Int_d [0]}), \forkHP1_CTf'''''''''_f'''''''''_In2_d , \writeMerge_data_CTf'''''''''_f'''''''''_Int_d );
  assign {\forkHP1_CTf'''''''''_f'''''''''_In2_r ,
          \writeMerge_data_CTf'''''''''_f'''''''''_Int_r } = {2 {(\dconWriteIn_CTf'''''''''_f'''''''''_Int_r  && \dconWriteIn_CTf'''''''''_f'''''''''_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTf'''''''''_f'''''''''_Int,
      Dcon Pointer_CTf'''''''''_f'''''''''_Int) : [(forkHP1_CTf'''''''''_f'''''''''_In3,Word16#)] > (dconPtr_CTf'''''''''_f'''''''''_Int,Pointer_CTf'''''''''_f'''''''''_Int) */
  assign \dconPtr_CTf'''''''''_f'''''''''_Int_d  = \Pointer_CTf'''''''''_f'''''''''_Int_dc ((& {\forkHP1_CTf'''''''''_f'''''''''_In3_d [0]}), \forkHP1_CTf'''''''''_f'''''''''_In3_d );
  assign {\forkHP1_CTf'''''''''_f'''''''''_In3_r } = {1 {(\dconPtr_CTf'''''''''_f'''''''''_Int_r  && \dconPtr_CTf'''''''''_f'''''''''_Int_d [0])}};
  
  /* demux (Ty MemOut_CTf'''''''''_f'''''''''_Int,
       Ty Pointer_CTf'''''''''_f'''''''''_Int) : (memWriteOut_CTf'''''''''_f'''''''''_Int,MemOut_CTf'''''''''_f'''''''''_Int) (dconPtr_CTf'''''''''_f'''''''''_Int,Pointer_CTf'''''''''_f'''''''''_Int) > [(_169,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                                                                                           (demuxWriteResult_CTf'''''''''_f'''''''''_Int,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [1:0] \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTf'''''''''_f'''''''''_Int_d [0] && \dconPtr_CTf'''''''''_f'''''''''_Int_d [0]))
      unique case (\memWriteOut_CTf'''''''''_f'''''''''_Int_d [1:1])
        1'd0: \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd  = 2'd2;
        default: \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd  = 2'd0;
  assign _169_d = {\dconPtr_CTf'''''''''_f'''''''''_Int_d [16:1],
                   \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd [0]};
  assign \demuxWriteResult_CTf'''''''''_f'''''''''_Int_d  = {\dconPtr_CTf'''''''''_f'''''''''_Int_d [16:1],
                                                             \dconPtr_CTf'''''''''_f'''''''''_Int_onehotd [1]};
  assign \dconPtr_CTf'''''''''_f'''''''''_Int_r  = (| (\dconPtr_CTf'''''''''_f'''''''''_Int_onehotd  & {\demuxWriteResult_CTf'''''''''_f'''''''''_Int_r ,
                                                                                                        _169_r}));
  assign \memWriteOut_CTf'''''''''_f'''''''''_Int_r  = \dconPtr_CTf'''''''''_f'''''''''_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTf'_f'_Int,Word16#) */
  assign \initHP_CTf'_f'_Int_d  = {16'd0, go__9_d[0]};
  assign go__9_r = \initHP_CTf'_f'_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf'_f'_Int1,Go) > (incrHP_CTf'_f'_Int,Word16#) */
  assign \incrHP_CTf'_f'_Int_d  = {16'd1,
                                   \incrHP_CTf'_f'_Int1_d [0]};
  assign \incrHP_CTf'_f'_Int1_r  = \incrHP_CTf'_f'_Int_r ;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTf'_f'_Int2,Go)] > (incrHP_mergeCTf'_f'_Int,Go) */
  logic [1:0] \incrHP_mergeCTf'_f'_Int_selected ;
  logic [1:0] \incrHP_mergeCTf'_f'_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTf'_f'_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTf'_f'_Int_select ))
        \incrHP_mergeCTf'_f'_Int_selected  = \incrHP_mergeCTf'_f'_Int_select ;
      else
        if (go__10_d[0]) \incrHP_mergeCTf'_f'_Int_selected [0] = 1'd1;
        else if (\incrHP_CTf'_f'_Int2_d [0])
          \incrHP_mergeCTf'_f'_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_f'_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTf'_f'_Int_select  <= (\incrHP_mergeCTf'_f'_Int_r  ? 2'd0 :
                                           \incrHP_mergeCTf'_f'_Int_selected );
  always_comb
    if (\incrHP_mergeCTf'_f'_Int_selected [0])
      \incrHP_mergeCTf'_f'_Int_d  = go__10_d;
    else if (\incrHP_mergeCTf'_f'_Int_selected [1])
      \incrHP_mergeCTf'_f'_Int_d  = \incrHP_CTf'_f'_Int2_d ;
    else \incrHP_mergeCTf'_f'_Int_d  = 1'd0;
  assign {\incrHP_CTf'_f'_Int2_r ,
          go__10_r} = (\incrHP_mergeCTf'_f'_Int_r  ? \incrHP_mergeCTf'_f'_Int_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf'_f'_Int_buf,Go) > [(incrHP_CTf'_f'_Int1,Go),
                                                   (incrHP_CTf'_f'_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTf'_f'_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf'_f'_Int_buf_done ;
  assign \incrHP_CTf'_f'_Int1_d  = (\incrHP_mergeCTf'_f'_Int_buf_d [0] && (! \incrHP_mergeCTf'_f'_Int_buf_emitted [0]));
  assign \incrHP_CTf'_f'_Int2_d  = (\incrHP_mergeCTf'_f'_Int_buf_d [0] && (! \incrHP_mergeCTf'_f'_Int_buf_emitted [1]));
  assign \incrHP_mergeCTf'_f'_Int_buf_done  = (\incrHP_mergeCTf'_f'_Int_buf_emitted  | ({\incrHP_CTf'_f'_Int2_d [0],
                                                                                         \incrHP_CTf'_f'_Int1_d [0]} & {\incrHP_CTf'_f'_Int2_r ,
                                                                                                                        \incrHP_CTf'_f'_Int1_r }));
  assign \incrHP_mergeCTf'_f'_Int_buf_r  = (& \incrHP_mergeCTf'_f'_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_f'_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf'_f'_Int_buf_emitted  <= (\incrHP_mergeCTf'_f'_Int_buf_r  ? 2'd0 :
                                                \incrHP_mergeCTf'_f'_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf'_f'_Int,Word16#) (forkHP1_CTf'_f'_Int,Word16#) > (addHP_CTf'_f'_Int,Word16#) */
  assign \addHP_CTf'_f'_Int_d  = {(\incrHP_CTf'_f'_Int_d [16:1] + \forkHP1_CTf'_f'_Int_d [16:1]),
                                  (\incrHP_CTf'_f'_Int_d [0] && \forkHP1_CTf'_f'_Int_d [0])};
  assign {\incrHP_CTf'_f'_Int_r ,
          \forkHP1_CTf'_f'_Int_r } = {2 {(\addHP_CTf'_f'_Int_r  && \addHP_CTf'_f'_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf'_f'_Int,Word16#),
                      (addHP_CTf'_f'_Int,Word16#)] > (mergeHP_CTf'_f'_Int,Word16#) */
  logic [1:0] \mergeHP_CTf'_f'_Int_selected ;
  logic [1:0] \mergeHP_CTf'_f'_Int_select ;
  always_comb
    begin
      \mergeHP_CTf'_f'_Int_selected  = 2'd0;
      if ((| \mergeHP_CTf'_f'_Int_select ))
        \mergeHP_CTf'_f'_Int_selected  = \mergeHP_CTf'_f'_Int_select ;
      else
        if (\initHP_CTf'_f'_Int_d [0])
          \mergeHP_CTf'_f'_Int_selected [0] = 1'd1;
        else if (\addHP_CTf'_f'_Int_d [0])
          \mergeHP_CTf'_f'_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_f'_Int_select  <= 2'd0;
    else
      \mergeHP_CTf'_f'_Int_select  <= (\mergeHP_CTf'_f'_Int_r  ? 2'd0 :
                                       \mergeHP_CTf'_f'_Int_selected );
  always_comb
    if (\mergeHP_CTf'_f'_Int_selected [0])
      \mergeHP_CTf'_f'_Int_d  = \initHP_CTf'_f'_Int_d ;
    else if (\mergeHP_CTf'_f'_Int_selected [1])
      \mergeHP_CTf'_f'_Int_d  = \addHP_CTf'_f'_Int_d ;
    else \mergeHP_CTf'_f'_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTf'_f'_Int_r ,
          \initHP_CTf'_f'_Int_r } = (\mergeHP_CTf'_f'_Int_r  ? \mergeHP_CTf'_f'_Int_selected  :
                                     2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf'_f'_Int,Go) > (incrHP_mergeCTf'_f'_Int_buf,Go) */
  Go_t \incrHP_mergeCTf'_f'_Int_bufchan_d ;
  logic \incrHP_mergeCTf'_f'_Int_bufchan_r ;
  assign \incrHP_mergeCTf'_f'_Int_r  = ((! \incrHP_mergeCTf'_f'_Int_bufchan_d [0]) || \incrHP_mergeCTf'_f'_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_f'_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf'_f'_Int_r )
        \incrHP_mergeCTf'_f'_Int_bufchan_d  <= \incrHP_mergeCTf'_f'_Int_d ;
  Go_t \incrHP_mergeCTf'_f'_Int_bufchan_buf ;
  assign \incrHP_mergeCTf'_f'_Int_bufchan_r  = (! \incrHP_mergeCTf'_f'_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTf'_f'_Int_buf_d  = (\incrHP_mergeCTf'_f'_Int_bufchan_buf [0] ? \incrHP_mergeCTf'_f'_Int_bufchan_buf  :
                                            \incrHP_mergeCTf'_f'_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \incrHP_mergeCTf'_f'_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf'_f'_Int_buf_r  && \incrHP_mergeCTf'_f'_Int_bufchan_buf [0]))
        \incrHP_mergeCTf'_f'_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf'_f'_Int_buf_r ) && (! \incrHP_mergeCTf'_f'_Int_bufchan_buf [0])))
        \incrHP_mergeCTf'_f'_Int_bufchan_buf  <= \incrHP_mergeCTf'_f'_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf'_f'_Int,Word16#) > (mergeHP_CTf'_f'_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf'_f'_Int_bufchan_d ;
  logic \mergeHP_CTf'_f'_Int_bufchan_r ;
  assign \mergeHP_CTf'_f'_Int_r  = ((! \mergeHP_CTf'_f'_Int_bufchan_d [0]) || \mergeHP_CTf'_f'_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf'_f'_Int_r )
        \mergeHP_CTf'_f'_Int_bufchan_d  <= \mergeHP_CTf'_f'_Int_d ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_bufchan_buf ;
  assign \mergeHP_CTf'_f'_Int_bufchan_r  = (! \mergeHP_CTf'_f'_Int_bufchan_buf [0]);
  assign \mergeHP_CTf'_f'_Int_buf_d  = (\mergeHP_CTf'_f'_Int_bufchan_buf [0] ? \mergeHP_CTf'_f'_Int_bufchan_buf  :
                                        \mergeHP_CTf'_f'_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf'_f'_Int_buf_r  && \mergeHP_CTf'_f'_Int_bufchan_buf [0]))
        \mergeHP_CTf'_f'_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf'_f'_Int_buf_r ) && (! \mergeHP_CTf'_f'_Int_bufchan_buf [0])))
        \mergeHP_CTf'_f'_Int_bufchan_buf  <= \mergeHP_CTf'_f'_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf'_f'_Int_buf,Word16#) > [(forkHP1_CTf'_f'_Int,Word16#),
                                                         (forkHP1_CTf'_f'_In2,Word16#),
                                                         (forkHP1_CTf'_f'_In3,Word16#)] */
  logic [2:0] \mergeHP_CTf'_f'_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTf'_f'_Int_buf_done ;
  assign \forkHP1_CTf'_f'_Int_d  = {\mergeHP_CTf'_f'_Int_buf_d [16:1],
                                    (\mergeHP_CTf'_f'_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_buf_emitted [0]))};
  assign \forkHP1_CTf'_f'_In2_d  = {\mergeHP_CTf'_f'_Int_buf_d [16:1],
                                    (\mergeHP_CTf'_f'_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_buf_emitted [1]))};
  assign \forkHP1_CTf'_f'_In3_d  = {\mergeHP_CTf'_f'_Int_buf_d [16:1],
                                    (\mergeHP_CTf'_f'_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_buf_emitted [2]))};
  assign \mergeHP_CTf'_f'_Int_buf_done  = (\mergeHP_CTf'_f'_Int_buf_emitted  | ({\forkHP1_CTf'_f'_In3_d [0],
                                                                                 \forkHP1_CTf'_f'_In2_d [0],
                                                                                 \forkHP1_CTf'_f'_Int_d [0]} & {\forkHP1_CTf'_f'_In3_r ,
                                                                                                                \forkHP1_CTf'_f'_In2_r ,
                                                                                                                \forkHP1_CTf'_f'_Int_r }));
  assign \mergeHP_CTf'_f'_Int_buf_r  = (& \mergeHP_CTf'_f'_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTf'_f'_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf'_f'_Int_buf_emitted  <= (\mergeHP_CTf'_f'_Int_buf_r  ? 3'd0 :
                                            \mergeHP_CTf'_f'_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf'_f'_Int) : [(dconReadIn_CTf'_f'_Int,MemIn_CTf'_f'_Int),
                                    (dconWriteIn_CTf'_f'_Int,MemIn_CTf'_f'_Int)] > (memMergeChoice_CTf'_f'_Int,C2) (memMergeIn_CTf'_f'_Int,MemIn_CTf'_f'_Int) */
  logic [1:0] \dconReadIn_CTf'_f'_Int_select_d ;
  assign \dconReadIn_CTf'_f'_Int_select_d  = ((| \dconReadIn_CTf'_f'_Int_select_q ) ? \dconReadIn_CTf'_f'_Int_select_q  :
                                              (\dconReadIn_CTf'_f'_Int_d [0] ? 2'd1 :
                                               (\dconWriteIn_CTf'_f'_Int_d [0] ? 2'd2 :
                                                2'd0)));
  logic [1:0] \dconReadIn_CTf'_f'_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf'_f'_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTf'_f'_Int_select_q  <= (\dconReadIn_CTf'_f'_Int_done  ? 2'd0 :
                                            \dconReadIn_CTf'_f'_Int_select_d );
  logic [1:0] \dconReadIn_CTf'_f'_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \dconReadIn_CTf'_f'_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf'_f'_Int_emit_q  <= (\dconReadIn_CTf'_f'_Int_done  ? 2'd0 :
                                          \dconReadIn_CTf'_f'_Int_emit_d );
  logic [1:0] \dconReadIn_CTf'_f'_Int_emit_d ;
  assign \dconReadIn_CTf'_f'_Int_emit_d  = (\dconReadIn_CTf'_f'_Int_emit_q  | ({\memMergeChoice_CTf'_f'_Int_d [0],
                                                                                \memMergeIn_CTf'_f'_Int_d [0]} & {\memMergeChoice_CTf'_f'_Int_r ,
                                                                                                                  \memMergeIn_CTf'_f'_Int_r }));
  logic \dconReadIn_CTf'_f'_Int_done ;
  assign \dconReadIn_CTf'_f'_Int_done  = (& \dconReadIn_CTf'_f'_Int_emit_d );
  assign {\dconWriteIn_CTf'_f'_Int_r ,
          \dconReadIn_CTf'_f'_Int_r } = (\dconReadIn_CTf'_f'_Int_done  ? \dconReadIn_CTf'_f'_Int_select_d  :
                                         2'd0);
  assign \memMergeIn_CTf'_f'_Int_d  = ((\dconReadIn_CTf'_f'_Int_select_d [0] && (! \dconReadIn_CTf'_f'_Int_emit_q [0])) ? \dconReadIn_CTf'_f'_Int_d  :
                                       ((\dconReadIn_CTf'_f'_Int_select_d [1] && (! \dconReadIn_CTf'_f'_Int_emit_q [0])) ? \dconWriteIn_CTf'_f'_Int_d  :
                                        {132'd0, 1'd0}));
  assign \memMergeChoice_CTf'_f'_Int_d  = ((\dconReadIn_CTf'_f'_Int_select_d [0] && (! \dconReadIn_CTf'_f'_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                           ((\dconReadIn_CTf'_f'_Int_select_d [1] && (! \dconReadIn_CTf'_f'_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                            {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf'_f'_Int,
      Ty MemOut_CTf'_f'_Int) : (memMergeIn_CTf'_f'_Int_dbuf,MemIn_CTf'_f'_Int) > (memOut_CTf'_f'_Int,MemOut_CTf'_f'_Int) */
  logic [114:0] \memMergeIn_CTf'_f'_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf'_f'_Int_dbuf_address ;
  logic [114:0] \memMergeIn_CTf'_f'_Int_dbuf_din ;
  logic [114:0] \memOut_CTf'_f'_Int_q ;
  logic \memOut_CTf'_f'_Int_valid ;
  logic \memMergeIn_CTf'_f'_Int_dbuf_we ;
  logic \memOut_CTf'_f'_Int_we ;
  assign \memMergeIn_CTf'_f'_Int_dbuf_din  = \memMergeIn_CTf'_f'_Int_dbuf_d [132:18];
  assign \memMergeIn_CTf'_f'_Int_dbuf_address  = \memMergeIn_CTf'_f'_Int_dbuf_d [17:2];
  assign \memMergeIn_CTf'_f'_Int_dbuf_we  = (\memMergeIn_CTf'_f'_Int_dbuf_d [1:1] && \memMergeIn_CTf'_f'_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf'_f'_Int_we  <= 1'd0;
        \memOut_CTf'_f'_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf'_f'_Int_we  <= \memMergeIn_CTf'_f'_Int_dbuf_we ;
        \memOut_CTf'_f'_Int_valid  <= \memMergeIn_CTf'_f'_Int_dbuf_d [0];
        if (\memMergeIn_CTf'_f'_Int_dbuf_we )
          begin
            \memMergeIn_CTf'_f'_Int_dbuf_mem [\memMergeIn_CTf'_f'_Int_dbuf_address ] <= \memMergeIn_CTf'_f'_Int_dbuf_din ;
            \memOut_CTf'_f'_Int_q  <= \memMergeIn_CTf'_f'_Int_dbuf_din ;
          end
        else
          \memOut_CTf'_f'_Int_q  <= \memMergeIn_CTf'_f'_Int_dbuf_mem [\memMergeIn_CTf'_f'_Int_dbuf_address ];
      end
  assign \memOut_CTf'_f'_Int_d  = {\memOut_CTf'_f'_Int_q ,
                                   \memOut_CTf'_f'_Int_we ,
                                   \memOut_CTf'_f'_Int_valid };
  assign \memMergeIn_CTf'_f'_Int_dbuf_r  = ((! \memOut_CTf'_f'_Int_valid ) || \memOut_CTf'_f'_Int_r );
  
  /* demux (Ty C2,
       Ty MemOut_CTf'_f'_Int) : (memMergeChoice_CTf'_f'_Int,C2) (memOut_CTf'_f'_Int_dbuf,MemOut_CTf'_f'_Int) > [(memReadOut_CTf'_f'_Int,MemOut_CTf'_f'_Int),
                                                                                                                (memWriteOut_CTf'_f'_Int,MemOut_CTf'_f'_Int)] */
  logic [1:0] \memOut_CTf'_f'_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf'_f'_Int_d [0] && \memOut_CTf'_f'_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTf'_f'_Int_d [1:1])
        1'd0: \memOut_CTf'_f'_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf'_f'_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf'_f'_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf'_f'_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf'_f'_Int_d  = {\memOut_CTf'_f'_Int_dbuf_d [116:1],
                                       \memOut_CTf'_f'_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTf'_f'_Int_d  = {\memOut_CTf'_f'_Int_dbuf_d [116:1],
                                        \memOut_CTf'_f'_Int_dbuf_onehotd [1]};
  assign \memOut_CTf'_f'_Int_dbuf_r  = (| (\memOut_CTf'_f'_Int_dbuf_onehotd  & {\memWriteOut_CTf'_f'_Int_r ,
                                                                                \memReadOut_CTf'_f'_Int_r }));
  assign \memMergeChoice_CTf'_f'_Int_r  = \memOut_CTf'_f'_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf'_f'_Int) : (memMergeIn_CTf'_f'_Int_rbuf,MemIn_CTf'_f'_Int) > (memMergeIn_CTf'_f'_Int_dbuf,MemIn_CTf'_f'_Int) */
  assign \memMergeIn_CTf'_f'_Int_rbuf_r  = ((! \memMergeIn_CTf'_f'_Int_dbuf_d [0]) || \memMergeIn_CTf'_f'_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'_f'_Int_dbuf_d  <= {132'd0, 1'd0};
    else
      if (\memMergeIn_CTf'_f'_Int_rbuf_r )
        \memMergeIn_CTf'_f'_Int_dbuf_d  <= \memMergeIn_CTf'_f'_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf'_f'_Int) : (memMergeIn_CTf'_f'_Int,MemIn_CTf'_f'_Int) > (memMergeIn_CTf'_f'_Int_rbuf,MemIn_CTf'_f'_Int) */
  \MemIn_CTf'_f'_Int_t  \memMergeIn_CTf'_f'_Int_buf ;
  assign \memMergeIn_CTf'_f'_Int_r  = (! \memMergeIn_CTf'_f'_Int_buf [0]);
  assign \memMergeIn_CTf'_f'_Int_rbuf_d  = (\memMergeIn_CTf'_f'_Int_buf [0] ? \memMergeIn_CTf'_f'_Int_buf  :
                                            \memMergeIn_CTf'_f'_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'_f'_Int_buf  <= {132'd0, 1'd0};
    else
      if ((\memMergeIn_CTf'_f'_Int_rbuf_r  && \memMergeIn_CTf'_f'_Int_buf [0]))
        \memMergeIn_CTf'_f'_Int_buf  <= {132'd0, 1'd0};
      else if (((! \memMergeIn_CTf'_f'_Int_rbuf_r ) && (! \memMergeIn_CTf'_f'_Int_buf [0])))
        \memMergeIn_CTf'_f'_Int_buf  <= \memMergeIn_CTf'_f'_Int_d ;
  
  /* dbuf (Ty MemOut_CTf'_f'_Int) : (memOut_CTf'_f'_Int_rbuf,MemOut_CTf'_f'_Int) > (memOut_CTf'_f'_Int_dbuf,MemOut_CTf'_f'_Int) */
  assign \memOut_CTf'_f'_Int_rbuf_r  = ((! \memOut_CTf'_f'_Int_dbuf_d [0]) || \memOut_CTf'_f'_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memOut_CTf'_f'_Int_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memOut_CTf'_f'_Int_rbuf_r )
        \memOut_CTf'_f'_Int_dbuf_d  <= \memOut_CTf'_f'_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf'_f'_Int) : (memOut_CTf'_f'_Int,MemOut_CTf'_f'_Int) > (memOut_CTf'_f'_Int_rbuf,MemOut_CTf'_f'_Int) */
  \MemOut_CTf'_f'_Int_t  \memOut_CTf'_f'_Int_buf ;
  assign \memOut_CTf'_f'_Int_r  = (! \memOut_CTf'_f'_Int_buf [0]);
  assign \memOut_CTf'_f'_Int_rbuf_d  = (\memOut_CTf'_f'_Int_buf [0] ? \memOut_CTf'_f'_Int_buf  :
                                        \memOut_CTf'_f'_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \memOut_CTf'_f'_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memOut_CTf'_f'_Int_rbuf_r  && \memOut_CTf'_f'_Int_buf [0]))
        \memOut_CTf'_f'_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memOut_CTf'_f'_Int_rbuf_r ) && (! \memOut_CTf'_f'_Int_buf [0])))
        \memOut_CTf'_f'_Int_buf  <= \memOut_CTf'_f'_Int_d ;
  
  /* destruct (Ty Pointer_CTf'_f'_Int,
          Dcon Pointer_CTf'_f'_Int) : (scfarg_0_2_1_argbuf,Pointer_CTf'_f'_Int) > [(destructReadIn_CTf'_f'_Int,Word16#)] */
  assign \destructReadIn_CTf'_f'_Int_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                           scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTf'_f'_Int_r ;
  
  /* dcon (Ty MemIn_CTf'_f'_Int,
      Dcon ReadIn_CTf'_f'_Int) : [(destructReadIn_CTf'_f'_Int,Word16#)] > (dconReadIn_CTf'_f'_Int,MemIn_CTf'_f'_Int) */
  assign \dconReadIn_CTf'_f'_Int_d  = \ReadIn_CTf'_f'_Int_dc ((& {\destructReadIn_CTf'_f'_Int_d [0]}), \destructReadIn_CTf'_f'_Int_d );
  assign {\destructReadIn_CTf'_f'_Int_r } = {1 {(\dconReadIn_CTf'_f'_Int_r  && \dconReadIn_CTf'_f'_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTf'_f'_Int,
          Dcon ReadOut_CTf'_f'_Int) : (memReadOut_CTf'_f'_Int,MemOut_CTf'_f'_Int) > [(readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf,CTf'_f'_Int)] */
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_d  = {\memReadOut_CTf'_f'_Int_d [116:2],
                                                           \memReadOut_CTf'_f'_Int_d [0]};
  assign \memReadOut_CTf'_f'_Int_r  = \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf'_f'_Int) : [(lizzieLet21_1_argbuf,CTf'_f'_Int),
                              (lizzieLet44_1_argbuf,CTf'_f'_Int),
                              (lizzieLet56_1_argbuf,CTf'_f'_Int),
                              (lizzieLet57_1_argbuf,CTf'_f'_Int),
                              (lizzieLet58_1_argbuf,CTf'_f'_Int)] > (writeMerge_choice_CTf'_f'_Int,C5) (writeMerge_data_CTf'_f'_Int,CTf'_f'_Int) */
  logic [4:0] lizzieLet21_1_argbuf_select_d;
  assign lizzieLet21_1_argbuf_select_d = ((| lizzieLet21_1_argbuf_select_q) ? lizzieLet21_1_argbuf_select_q :
                                          (lizzieLet21_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet44_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet56_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet57_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet58_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet21_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet21_1_argbuf_select_q <= (lizzieLet21_1_argbuf_done ? 5'd0 :
                                        lizzieLet21_1_argbuf_select_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet21_1_argbuf_emit_q <= (lizzieLet21_1_argbuf_done ? 2'd0 :
                                      lizzieLet21_1_argbuf_emit_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_d;
  assign lizzieLet21_1_argbuf_emit_d = (lizzieLet21_1_argbuf_emit_q | ({\writeMerge_choice_CTf'_f'_Int_d [0],
                                                                        \writeMerge_data_CTf'_f'_Int_d [0]} & {\writeMerge_choice_CTf'_f'_Int_r ,
                                                                                                               \writeMerge_data_CTf'_f'_Int_r }));
  logic lizzieLet21_1_argbuf_done;
  assign lizzieLet21_1_argbuf_done = (& lizzieLet21_1_argbuf_emit_d);
  assign {lizzieLet58_1_argbuf_r,
          lizzieLet57_1_argbuf_r,
          lizzieLet56_1_argbuf_r,
          lizzieLet44_1_argbuf_r,
          lizzieLet21_1_argbuf_r} = (lizzieLet21_1_argbuf_done ? lizzieLet21_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTf'_f'_Int_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                            ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet44_1_argbuf_d :
                                             ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet56_1_argbuf_d :
                                              ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet57_1_argbuf_d :
                                               ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet58_1_argbuf_d :
                                                {115'd0, 1'd0})))));
  assign \writeMerge_choice_CTf'_f'_Int_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                              ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                               ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                 ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                  {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf'_f'_Int) : (writeMerge_choice_CTf'_f'_Int,C5) (demuxWriteResult_CTf'_f'_Int,Pointer_CTf'_f'_Int) > [(writeCTf'_f'_IntlizzieLet21_1_argbuf,Pointer_CTf'_f'_Int),
                                                                                                                          (writeCTf'_f'_IntlizzieLet44_1_argbuf,Pointer_CTf'_f'_Int),
                                                                                                                          (writeCTf'_f'_IntlizzieLet56_1_argbuf,Pointer_CTf'_f'_Int),
                                                                                                                          (writeCTf'_f'_IntlizzieLet57_1_argbuf,Pointer_CTf'_f'_Int),
                                                                                                                          (writeCTf'_f'_IntlizzieLet58_1_argbuf,Pointer_CTf'_f'_Int)] */
  logic [4:0] \demuxWriteResult_CTf'_f'_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf'_f'_Int_d [0] && \demuxWriteResult_CTf'_f'_Int_d [0]))
      unique case (\writeMerge_choice_CTf'_f'_Int_d [3:1])
        3'd0: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd16;
        default: \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf'_f'_Int_onehotd  = 5'd0;
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_d [16:1],
                                                     \demuxWriteResult_CTf'_f'_Int_onehotd [0]};
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_d [16:1],
                                                     \demuxWriteResult_CTf'_f'_Int_onehotd [1]};
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_d [16:1],
                                                     \demuxWriteResult_CTf'_f'_Int_onehotd [2]};
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_d [16:1],
                                                     \demuxWriteResult_CTf'_f'_Int_onehotd [3]};
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_d [16:1],
                                                     \demuxWriteResult_CTf'_f'_Int_onehotd [4]};
  assign \demuxWriteResult_CTf'_f'_Int_r  = (| (\demuxWriteResult_CTf'_f'_Int_onehotd  & {\writeCTf'_f'_IntlizzieLet58_1_argbuf_r ,
                                                                                          \writeCTf'_f'_IntlizzieLet57_1_argbuf_r ,
                                                                                          \writeCTf'_f'_IntlizzieLet56_1_argbuf_r ,
                                                                                          \writeCTf'_f'_IntlizzieLet44_1_argbuf_r ,
                                                                                          \writeCTf'_f'_IntlizzieLet21_1_argbuf_r }));
  assign \writeMerge_choice_CTf'_f'_Int_r  = \demuxWriteResult_CTf'_f'_Int_r ;
  
  /* dcon (Ty MemIn_CTf'_f'_Int,
      Dcon WriteIn_CTf'_f'_Int) : [(forkHP1_CTf'_f'_In2,Word16#),
                                   (writeMerge_data_CTf'_f'_Int,CTf'_f'_Int)] > (dconWriteIn_CTf'_f'_Int,MemIn_CTf'_f'_Int) */
  assign \dconWriteIn_CTf'_f'_Int_d  = \WriteIn_CTf'_f'_Int_dc ((& {\forkHP1_CTf'_f'_In2_d [0],
                                                                    \writeMerge_data_CTf'_f'_Int_d [0]}), \forkHP1_CTf'_f'_In2_d , \writeMerge_data_CTf'_f'_Int_d );
  assign {\forkHP1_CTf'_f'_In2_r ,
          \writeMerge_data_CTf'_f'_Int_r } = {2 {(\dconWriteIn_CTf'_f'_Int_r  && \dconWriteIn_CTf'_f'_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTf'_f'_Int,
      Dcon Pointer_CTf'_f'_Int) : [(forkHP1_CTf'_f'_In3,Word16#)] > (dconPtr_CTf'_f'_Int,Pointer_CTf'_f'_Int) */
  assign \dconPtr_CTf'_f'_Int_d  = \Pointer_CTf'_f'_Int_dc ((& {\forkHP1_CTf'_f'_In3_d [0]}), \forkHP1_CTf'_f'_In3_d );
  assign {\forkHP1_CTf'_f'_In3_r } = {1 {(\dconPtr_CTf'_f'_Int_r  && \dconPtr_CTf'_f'_Int_d [0])}};
  
  /* demux (Ty MemOut_CTf'_f'_Int,
       Ty Pointer_CTf'_f'_Int) : (memWriteOut_CTf'_f'_Int,MemOut_CTf'_f'_Int) (dconPtr_CTf'_f'_Int,Pointer_CTf'_f'_Int) > [(_168,Pointer_CTf'_f'_Int),
                                                                                                                           (demuxWriteResult_CTf'_f'_Int,Pointer_CTf'_f'_Int)] */
  logic [1:0] \dconPtr_CTf'_f'_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTf'_f'_Int_d [0] && \dconPtr_CTf'_f'_Int_d [0]))
      unique case (\memWriteOut_CTf'_f'_Int_d [1:1])
        1'd0: \dconPtr_CTf'_f'_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf'_f'_Int_onehotd  = 2'd2;
        default: \dconPtr_CTf'_f'_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf'_f'_Int_onehotd  = 2'd0;
  assign _168_d = {\dconPtr_CTf'_f'_Int_d [16:1],
                   \dconPtr_CTf'_f'_Int_onehotd [0]};
  assign \demuxWriteResult_CTf'_f'_Int_d  = {\dconPtr_CTf'_f'_Int_d [16:1],
                                             \dconPtr_CTf'_f'_Int_onehotd [1]};
  assign \dconPtr_CTf'_f'_Int_r  = (| (\dconPtr_CTf'_f'_Int_onehotd  & {\demuxWriteResult_CTf'_f'_Int_r ,
                                                                        _168_r}));
  assign \memWriteOut_CTf'_f'_Int_r  = \dconPtr_CTf'_f'_Int_r ;
  
  /* const (Ty Word16#,Lit 0) : (go__11,Go) > (initHP_CTf_f_Int,Word16#) */
  assign initHP_CTf_f_Int_d = {16'd0, go__11_d[0]};
  assign go__11_r = initHP_CTf_f_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf_f_Int1,Go) > (incrHP_CTf_f_Int,Word16#) */
  assign incrHP_CTf_f_Int_d = {16'd1, incrHP_CTf_f_Int1_d[0]};
  assign incrHP_CTf_f_Int1_r = incrHP_CTf_f_Int_r;
  
  /* merge (Ty Go) : [(go__12,Go),
                 (incrHP_CTf_f_Int2,Go)] > (incrHP_mergeCTf_f_Int,Go) */
  logic [1:0] incrHP_mergeCTf_f_Int_selected;
  logic [1:0] incrHP_mergeCTf_f_Int_select;
  always_comb
    begin
      incrHP_mergeCTf_f_Int_selected = 2'd0;
      if ((| incrHP_mergeCTf_f_Int_select))
        incrHP_mergeCTf_f_Int_selected = incrHP_mergeCTf_f_Int_select;
      else
        if (go__12_d[0]) incrHP_mergeCTf_f_Int_selected[0] = 1'd1;
        else if (incrHP_CTf_f_Int2_d[0])
          incrHP_mergeCTf_f_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_select <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_select <= (incrHP_mergeCTf_f_Int_r ? 2'd0 :
                                       incrHP_mergeCTf_f_Int_selected);
  always_comb
    if (incrHP_mergeCTf_f_Int_selected[0])
      incrHP_mergeCTf_f_Int_d = go__12_d;
    else if (incrHP_mergeCTf_f_Int_selected[1])
      incrHP_mergeCTf_f_Int_d = incrHP_CTf_f_Int2_d;
    else incrHP_mergeCTf_f_Int_d = 1'd0;
  assign {incrHP_CTf_f_Int2_r,
          go__12_r} = (incrHP_mergeCTf_f_Int_r ? incrHP_mergeCTf_f_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_f_Int_buf,Go) > [(incrHP_CTf_f_Int1,Go),
                                                 (incrHP_CTf_f_Int2,Go)] */
  logic [1:0] incrHP_mergeCTf_f_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTf_f_Int_buf_done;
  assign incrHP_CTf_f_Int1_d = (incrHP_mergeCTf_f_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_buf_emitted[0]));
  assign incrHP_CTf_f_Int2_d = (incrHP_mergeCTf_f_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_buf_emitted[1]));
  assign incrHP_mergeCTf_f_Int_buf_done = (incrHP_mergeCTf_f_Int_buf_emitted | ({incrHP_CTf_f_Int2_d[0],
                                                                                 incrHP_CTf_f_Int1_d[0]} & {incrHP_CTf_f_Int2_r,
                                                                                                            incrHP_CTf_f_Int1_r}));
  assign incrHP_mergeCTf_f_Int_buf_r = (& incrHP_mergeCTf_f_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_buf_emitted <= (incrHP_mergeCTf_f_Int_buf_r ? 2'd0 :
                                            incrHP_mergeCTf_f_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf_f_Int,Word16#) (forkHP1_CTf_f_Int,Word16#) > (addHP_CTf_f_Int,Word16#) */
  assign addHP_CTf_f_Int_d = {(incrHP_CTf_f_Int_d[16:1] + forkHP1_CTf_f_Int_d[16:1]),
                              (incrHP_CTf_f_Int_d[0] && forkHP1_CTf_f_Int_d[0])};
  assign {incrHP_CTf_f_Int_r,
          forkHP1_CTf_f_Int_r} = {2 {(addHP_CTf_f_Int_r && addHP_CTf_f_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf_f_Int,Word16#),
                      (addHP_CTf_f_Int,Word16#)] > (mergeHP_CTf_f_Int,Word16#) */
  logic [1:0] mergeHP_CTf_f_Int_selected;
  logic [1:0] mergeHP_CTf_f_Int_select;
  always_comb
    begin
      mergeHP_CTf_f_Int_selected = 2'd0;
      if ((| mergeHP_CTf_f_Int_select))
        mergeHP_CTf_f_Int_selected = mergeHP_CTf_f_Int_select;
      else
        if (initHP_CTf_f_Int_d[0]) mergeHP_CTf_f_Int_selected[0] = 1'd1;
        else if (addHP_CTf_f_Int_d[0])
          mergeHP_CTf_f_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_select <= 2'd0;
    else
      mergeHP_CTf_f_Int_select <= (mergeHP_CTf_f_Int_r ? 2'd0 :
                                   mergeHP_CTf_f_Int_selected);
  always_comb
    if (mergeHP_CTf_f_Int_selected[0])
      mergeHP_CTf_f_Int_d = initHP_CTf_f_Int_d;
    else if (mergeHP_CTf_f_Int_selected[1])
      mergeHP_CTf_f_Int_d = addHP_CTf_f_Int_d;
    else mergeHP_CTf_f_Int_d = {16'd0, 1'd0};
  assign {addHP_CTf_f_Int_r,
          initHP_CTf_f_Int_r} = (mergeHP_CTf_f_Int_r ? mergeHP_CTf_f_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf_f_Int,Go) > (incrHP_mergeCTf_f_Int_buf,Go) */
  Go_t incrHP_mergeCTf_f_Int_bufchan_d;
  logic incrHP_mergeCTf_f_Int_bufchan_r;
  assign incrHP_mergeCTf_f_Int_r = ((! incrHP_mergeCTf_f_Int_bufchan_d[0]) || incrHP_mergeCTf_f_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_f_Int_r)
        incrHP_mergeCTf_f_Int_bufchan_d <= incrHP_mergeCTf_f_Int_d;
  Go_t incrHP_mergeCTf_f_Int_bufchan_buf;
  assign incrHP_mergeCTf_f_Int_bufchan_r = (! incrHP_mergeCTf_f_Int_bufchan_buf[0]);
  assign incrHP_mergeCTf_f_Int_buf_d = (incrHP_mergeCTf_f_Int_bufchan_buf[0] ? incrHP_mergeCTf_f_Int_bufchan_buf :
                                        incrHP_mergeCTf_f_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTf_f_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_f_Int_buf_r && incrHP_mergeCTf_f_Int_bufchan_buf[0]))
        incrHP_mergeCTf_f_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_f_Int_buf_r) && (! incrHP_mergeCTf_f_Int_bufchan_buf[0])))
        incrHP_mergeCTf_f_Int_bufchan_buf <= incrHP_mergeCTf_f_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf_f_Int,Word16#) > (mergeHP_CTf_f_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_f_Int_bufchan_d;
  logic mergeHP_CTf_f_Int_bufchan_r;
  assign mergeHP_CTf_f_Int_r = ((! mergeHP_CTf_f_Int_bufchan_d[0]) || mergeHP_CTf_f_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTf_f_Int_r)
        mergeHP_CTf_f_Int_bufchan_d <= mergeHP_CTf_f_Int_d;
  \Word16#_t  mergeHP_CTf_f_Int_bufchan_buf;
  assign mergeHP_CTf_f_Int_bufchan_r = (! mergeHP_CTf_f_Int_bufchan_buf[0]);
  assign mergeHP_CTf_f_Int_buf_d = (mergeHP_CTf_f_Int_bufchan_buf[0] ? mergeHP_CTf_f_Int_bufchan_buf :
                                    mergeHP_CTf_f_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_f_Int_buf_r && mergeHP_CTf_f_Int_bufchan_buf[0]))
        mergeHP_CTf_f_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_f_Int_buf_r) && (! mergeHP_CTf_f_Int_bufchan_buf[0])))
        mergeHP_CTf_f_Int_bufchan_buf <= mergeHP_CTf_f_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_f_Int_buf,Word16#) > [(forkHP1_CTf_f_Int,Word16#),
                                                       (forkHP1_CTf_f_In2,Word16#),
                                                       (forkHP1_CTf_f_In3,Word16#)] */
  logic [2:0] mergeHP_CTf_f_Int_buf_emitted;
  logic [2:0] mergeHP_CTf_f_Int_buf_done;
  assign forkHP1_CTf_f_Int_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[0]))};
  assign forkHP1_CTf_f_In2_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[1]))};
  assign forkHP1_CTf_f_In3_d = {mergeHP_CTf_f_Int_buf_d[16:1],
                                (mergeHP_CTf_f_Int_buf_d[0] && (! mergeHP_CTf_f_Int_buf_emitted[2]))};
  assign mergeHP_CTf_f_Int_buf_done = (mergeHP_CTf_f_Int_buf_emitted | ({forkHP1_CTf_f_In3_d[0],
                                                                         forkHP1_CTf_f_In2_d[0],
                                                                         forkHP1_CTf_f_Int_d[0]} & {forkHP1_CTf_f_In3_r,
                                                                                                    forkHP1_CTf_f_In2_r,
                                                                                                    forkHP1_CTf_f_Int_r}));
  assign mergeHP_CTf_f_Int_buf_r = (& mergeHP_CTf_f_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_f_Int_buf_emitted <= (mergeHP_CTf_f_Int_buf_r ? 3'd0 :
                                        mergeHP_CTf_f_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf_f_Int) : [(dconReadIn_CTf_f_Int,MemIn_CTf_f_Int),
                                  (dconWriteIn_CTf_f_Int,MemIn_CTf_f_Int)] > (memMergeChoice_CTf_f_Int,C2) (memMergeIn_CTf_f_Int,MemIn_CTf_f_Int) */
  logic [1:0] dconReadIn_CTf_f_Int_select_d;
  assign dconReadIn_CTf_f_Int_select_d = ((| dconReadIn_CTf_f_Int_select_q) ? dconReadIn_CTf_f_Int_select_q :
                                          (dconReadIn_CTf_f_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_CTf_f_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_CTf_f_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_select_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_select_q <= (dconReadIn_CTf_f_Int_done ? 2'd0 :
                                        dconReadIn_CTf_f_Int_select_d);
  logic [1:0] dconReadIn_CTf_f_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTf_f_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_emit_q <= (dconReadIn_CTf_f_Int_done ? 2'd0 :
                                      dconReadIn_CTf_f_Int_emit_d);
  logic [1:0] dconReadIn_CTf_f_Int_emit_d;
  assign dconReadIn_CTf_f_Int_emit_d = (dconReadIn_CTf_f_Int_emit_q | ({memMergeChoice_CTf_f_Int_d[0],
                                                                        memMergeIn_CTf_f_Int_d[0]} & {memMergeChoice_CTf_f_Int_r,
                                                                                                      memMergeIn_CTf_f_Int_r}));
  logic dconReadIn_CTf_f_Int_done;
  assign dconReadIn_CTf_f_Int_done = (& dconReadIn_CTf_f_Int_emit_d);
  assign {dconWriteIn_CTf_f_Int_r,
          dconReadIn_CTf_f_Int_r} = (dconReadIn_CTf_f_Int_done ? dconReadIn_CTf_f_Int_select_d :
                                     2'd0);
  assign memMergeIn_CTf_f_Int_d = ((dconReadIn_CTf_f_Int_select_d[0] && (! dconReadIn_CTf_f_Int_emit_q[0])) ? dconReadIn_CTf_f_Int_d :
                                   ((dconReadIn_CTf_f_Int_select_d[1] && (! dconReadIn_CTf_f_Int_emit_q[0])) ? dconWriteIn_CTf_f_Int_d :
                                    {180'd0, 1'd0}));
  assign memMergeChoice_CTf_f_Int_d = ((dconReadIn_CTf_f_Int_select_d[0] && (! dconReadIn_CTf_f_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_CTf_f_Int_select_d[1] && (! dconReadIn_CTf_f_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf_f_Int,
      Ty MemOut_CTf_f_Int) : (memMergeIn_CTf_f_Int_dbuf,MemIn_CTf_f_Int) > (memOut_CTf_f_Int,MemOut_CTf_f_Int) */
  logic [162:0] memMergeIn_CTf_f_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_f_Int_dbuf_address;
  logic [162:0] memMergeIn_CTf_f_Int_dbuf_din;
  logic [162:0] memOut_CTf_f_Int_q;
  logic memOut_CTf_f_Int_valid;
  logic memMergeIn_CTf_f_Int_dbuf_we;
  logic memOut_CTf_f_Int_we;
  assign memMergeIn_CTf_f_Int_dbuf_din = memMergeIn_CTf_f_Int_dbuf_d[180:18];
  assign memMergeIn_CTf_f_Int_dbuf_address = memMergeIn_CTf_f_Int_dbuf_d[17:2];
  assign memMergeIn_CTf_f_Int_dbuf_we = (memMergeIn_CTf_f_Int_dbuf_d[1:1] && memMergeIn_CTf_f_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_f_Int_we <= 1'd0;
        memOut_CTf_f_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_f_Int_we <= memMergeIn_CTf_f_Int_dbuf_we;
        memOut_CTf_f_Int_valid <= memMergeIn_CTf_f_Int_dbuf_d[0];
        if (memMergeIn_CTf_f_Int_dbuf_we)
          begin
            memMergeIn_CTf_f_Int_dbuf_mem[memMergeIn_CTf_f_Int_dbuf_address] <= memMergeIn_CTf_f_Int_dbuf_din;
            memOut_CTf_f_Int_q <= memMergeIn_CTf_f_Int_dbuf_din;
          end
        else
          memOut_CTf_f_Int_q <= memMergeIn_CTf_f_Int_dbuf_mem[memMergeIn_CTf_f_Int_dbuf_address];
      end
  assign memOut_CTf_f_Int_d = {memOut_CTf_f_Int_q,
                               memOut_CTf_f_Int_we,
                               memOut_CTf_f_Int_valid};
  assign memMergeIn_CTf_f_Int_dbuf_r = ((! memOut_CTf_f_Int_valid) || memOut_CTf_f_Int_r);
  
  /* demux (Ty C2,
       Ty MemOut_CTf_f_Int) : (memMergeChoice_CTf_f_Int,C2) (memOut_CTf_f_Int_dbuf,MemOut_CTf_f_Int) > [(memReadOut_CTf_f_Int,MemOut_CTf_f_Int),
                                                                                                        (memWriteOut_CTf_f_Int,MemOut_CTf_f_Int)] */
  logic [1:0] memOut_CTf_f_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_f_Int_d[0] && memOut_CTf_f_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTf_f_Int_d[1:1])
        1'd0: memOut_CTf_f_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_f_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTf_f_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_f_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_f_Int_d = {memOut_CTf_f_Int_dbuf_d[164:1],
                                   memOut_CTf_f_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTf_f_Int_d = {memOut_CTf_f_Int_dbuf_d[164:1],
                                    memOut_CTf_f_Int_dbuf_onehotd[1]};
  assign memOut_CTf_f_Int_dbuf_r = (| (memOut_CTf_f_Int_dbuf_onehotd & {memWriteOut_CTf_f_Int_r,
                                                                        memReadOut_CTf_f_Int_r}));
  assign memMergeChoice_CTf_f_Int_r = memOut_CTf_f_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf_f_Int) : (memMergeIn_CTf_f_Int_rbuf,MemIn_CTf_f_Int) > (memMergeIn_CTf_f_Int_dbuf,MemIn_CTf_f_Int) */
  assign memMergeIn_CTf_f_Int_rbuf_r = ((! memMergeIn_CTf_f_Int_dbuf_d[0]) || memMergeIn_CTf_f_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_Int_dbuf_d <= {180'd0, 1'd0};
    else
      if (memMergeIn_CTf_f_Int_rbuf_r)
        memMergeIn_CTf_f_Int_dbuf_d <= memMergeIn_CTf_f_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf_f_Int) : (memMergeIn_CTf_f_Int,MemIn_CTf_f_Int) > (memMergeIn_CTf_f_Int_rbuf,MemIn_CTf_f_Int) */
  MemIn_CTf_f_Int_t memMergeIn_CTf_f_Int_buf;
  assign memMergeIn_CTf_f_Int_r = (! memMergeIn_CTf_f_Int_buf[0]);
  assign memMergeIn_CTf_f_Int_rbuf_d = (memMergeIn_CTf_f_Int_buf[0] ? memMergeIn_CTf_f_Int_buf :
                                        memMergeIn_CTf_f_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CTf_f_Int_buf <= {180'd0, 1'd0};
    else
      if ((memMergeIn_CTf_f_Int_rbuf_r && memMergeIn_CTf_f_Int_buf[0]))
        memMergeIn_CTf_f_Int_buf <= {180'd0, 1'd0};
      else if (((! memMergeIn_CTf_f_Int_rbuf_r) && (! memMergeIn_CTf_f_Int_buf[0])))
        memMergeIn_CTf_f_Int_buf <= memMergeIn_CTf_f_Int_d;
  
  /* dbuf (Ty MemOut_CTf_f_Int) : (memOut_CTf_f_Int_rbuf,MemOut_CTf_f_Int) > (memOut_CTf_f_Int_dbuf,MemOut_CTf_f_Int) */
  assign memOut_CTf_f_Int_rbuf_r = ((! memOut_CTf_f_Int_dbuf_d[0]) || memOut_CTf_f_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_dbuf_d <= {164'd0, 1'd0};
    else
      if (memOut_CTf_f_Int_rbuf_r)
        memOut_CTf_f_Int_dbuf_d <= memOut_CTf_f_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf_f_Int) : (memOut_CTf_f_Int,MemOut_CTf_f_Int) > (memOut_CTf_f_Int_rbuf,MemOut_CTf_f_Int) */
  MemOut_CTf_f_Int_t memOut_CTf_f_Int_buf;
  assign memOut_CTf_f_Int_r = (! memOut_CTf_f_Int_buf[0]);
  assign memOut_CTf_f_Int_rbuf_d = (memOut_CTf_f_Int_buf[0] ? memOut_CTf_f_Int_buf :
                                    memOut_CTf_f_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTf_f_Int_buf <= {164'd0, 1'd0};
    else
      if ((memOut_CTf_f_Int_rbuf_r && memOut_CTf_f_Int_buf[0]))
        memOut_CTf_f_Int_buf <= {164'd0, 1'd0};
      else if (((! memOut_CTf_f_Int_rbuf_r) && (! memOut_CTf_f_Int_buf[0])))
        memOut_CTf_f_Int_buf <= memOut_CTf_f_Int_d;
  
  /* destruct (Ty Pointer_CTf_f_Int,
          Dcon Pointer_CTf_f_Int) : (scfarg_0_3_1_argbuf,Pointer_CTf_f_Int) > [(destructReadIn_CTf_f_Int,Word16#)] */
  assign destructReadIn_CTf_f_Int_d = {scfarg_0_3_1_argbuf_d[16:1],
                                       scfarg_0_3_1_argbuf_d[0]};
  assign scfarg_0_3_1_argbuf_r = destructReadIn_CTf_f_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int,
      Dcon ReadIn_CTf_f_Int) : [(destructReadIn_CTf_f_Int,Word16#)] > (dconReadIn_CTf_f_Int,MemIn_CTf_f_Int) */
  assign dconReadIn_CTf_f_Int_d = ReadIn_CTf_f_Int_dc((& {destructReadIn_CTf_f_Int_d[0]}), destructReadIn_CTf_f_Int_d);
  assign {destructReadIn_CTf_f_Int_r} = {1 {(dconReadIn_CTf_f_Int_r && dconReadIn_CTf_f_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTf_f_Int,
          Dcon ReadOut_CTf_f_Int) : (memReadOut_CTf_f_Int,MemOut_CTf_f_Int) > [(readPointer_CTf_f_Intscfarg_0_3_1_argbuf,CTf_f_Int)] */
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_d = {memReadOut_CTf_f_Int_d[164:2],
                                                       memReadOut_CTf_f_Int_d[0]};
  assign memReadOut_CTf_f_Int_r = readPointer_CTf_f_Intscfarg_0_3_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CTf_f_Int) : [(lizzieLet40_1_argbuf,CTf_f_Int),
                                  (lizzieLet45_1_argbuf,CTf_f_Int),
                                  (lizzieLet61_1_argbuf,CTf_f_Int),
                                  (lizzieLet62_1_argbuf,CTf_f_Int),
                                  (lizzieLet63_1_argbuf,CTf_f_Int)] > (writeMerge_choice_CTf_f_Int,C5) (writeMerge_data_CTf_f_Int,CTf_f_Int) */
  logic [4:0] lizzieLet40_1_argbuf_select_d;
  assign lizzieLet40_1_argbuf_select_d = ((| lizzieLet40_1_argbuf_select_q) ? lizzieLet40_1_argbuf_select_q :
                                          (lizzieLet40_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet45_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet61_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet62_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet63_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet40_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet40_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet40_1_argbuf_select_q <= (lizzieLet40_1_argbuf_done ? 5'd0 :
                                        lizzieLet40_1_argbuf_select_d);
  logic [1:0] lizzieLet40_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet40_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet40_1_argbuf_emit_q <= (lizzieLet40_1_argbuf_done ? 2'd0 :
                                      lizzieLet40_1_argbuf_emit_d);
  logic [1:0] lizzieLet40_1_argbuf_emit_d;
  assign lizzieLet40_1_argbuf_emit_d = (lizzieLet40_1_argbuf_emit_q | ({writeMerge_choice_CTf_f_Int_d[0],
                                                                        writeMerge_data_CTf_f_Int_d[0]} & {writeMerge_choice_CTf_f_Int_r,
                                                                                                           writeMerge_data_CTf_f_Int_r}));
  logic lizzieLet40_1_argbuf_done;
  assign lizzieLet40_1_argbuf_done = (& lizzieLet40_1_argbuf_emit_d);
  assign {lizzieLet63_1_argbuf_r,
          lizzieLet62_1_argbuf_r,
          lizzieLet61_1_argbuf_r,
          lizzieLet45_1_argbuf_r,
          lizzieLet40_1_argbuf_r} = (lizzieLet40_1_argbuf_done ? lizzieLet40_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_f_Int_d = ((lizzieLet40_1_argbuf_select_d[0] && (! lizzieLet40_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                        ((lizzieLet40_1_argbuf_select_d[1] && (! lizzieLet40_1_argbuf_emit_q[0])) ? lizzieLet45_1_argbuf_d :
                                         ((lizzieLet40_1_argbuf_select_d[2] && (! lizzieLet40_1_argbuf_emit_q[0])) ? lizzieLet61_1_argbuf_d :
                                          ((lizzieLet40_1_argbuf_select_d[3] && (! lizzieLet40_1_argbuf_emit_q[0])) ? lizzieLet62_1_argbuf_d :
                                           ((lizzieLet40_1_argbuf_select_d[4] && (! lizzieLet40_1_argbuf_emit_q[0])) ? lizzieLet63_1_argbuf_d :
                                            {163'd0, 1'd0})))));
  assign writeMerge_choice_CTf_f_Int_d = ((lizzieLet40_1_argbuf_select_d[0] && (! lizzieLet40_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                          ((lizzieLet40_1_argbuf_select_d[1] && (! lizzieLet40_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                           ((lizzieLet40_1_argbuf_select_d[2] && (! lizzieLet40_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                            ((lizzieLet40_1_argbuf_select_d[3] && (! lizzieLet40_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                             ((lizzieLet40_1_argbuf_select_d[4] && (! lizzieLet40_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf_f_Int) : (writeMerge_choice_CTf_f_Int,C5) (demuxWriteResult_CTf_f_Int,Pointer_CTf_f_Int) > [(writeCTf_f_IntlizzieLet40_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet45_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet61_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet62_1_argbuf,Pointer_CTf_f_Int),
                                                                                                                  (writeCTf_f_IntlizzieLet63_1_argbuf,Pointer_CTf_f_Int)] */
  logic [4:0] demuxWriteResult_CTf_f_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_f_Int_d[0] && demuxWriteResult_CTf_f_Int_d[0]))
      unique case (writeMerge_choice_CTf_f_Int_d[3:1])
        3'd0: demuxWriteResult_CTf_f_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_f_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_f_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_f_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_f_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTf_f_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_f_Int_onehotd = 5'd0;
  assign writeCTf_f_IntlizzieLet40_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[0]};
  assign writeCTf_f_IntlizzieLet45_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[1]};
  assign writeCTf_f_IntlizzieLet61_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[2]};
  assign writeCTf_f_IntlizzieLet62_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[3]};
  assign writeCTf_f_IntlizzieLet63_1_argbuf_d = {demuxWriteResult_CTf_f_Int_d[16:1],
                                                 demuxWriteResult_CTf_f_Int_onehotd[4]};
  assign demuxWriteResult_CTf_f_Int_r = (| (demuxWriteResult_CTf_f_Int_onehotd & {writeCTf_f_IntlizzieLet63_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet62_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet61_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet45_1_argbuf_r,
                                                                                  writeCTf_f_IntlizzieLet40_1_argbuf_r}));
  assign writeMerge_choice_CTf_f_Int_r = demuxWriteResult_CTf_f_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int,
      Dcon WriteIn_CTf_f_Int) : [(forkHP1_CTf_f_In2,Word16#),
                                 (writeMerge_data_CTf_f_Int,CTf_f_Int)] > (dconWriteIn_CTf_f_Int,MemIn_CTf_f_Int) */
  assign dconWriteIn_CTf_f_Int_d = WriteIn_CTf_f_Int_dc((& {forkHP1_CTf_f_In2_d[0],
                                                            writeMerge_data_CTf_f_Int_d[0]}), forkHP1_CTf_f_In2_d, writeMerge_data_CTf_f_Int_d);
  assign {forkHP1_CTf_f_In2_r,
          writeMerge_data_CTf_f_Int_r} = {2 {(dconWriteIn_CTf_f_Int_r && dconWriteIn_CTf_f_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTf_f_Int,
      Dcon Pointer_CTf_f_Int) : [(forkHP1_CTf_f_In3,Word16#)] > (dconPtr_CTf_f_Int,Pointer_CTf_f_Int) */
  assign dconPtr_CTf_f_Int_d = Pointer_CTf_f_Int_dc((& {forkHP1_CTf_f_In3_d[0]}), forkHP1_CTf_f_In3_d);
  assign {forkHP1_CTf_f_In3_r} = {1 {(dconPtr_CTf_f_Int_r && dconPtr_CTf_f_Int_d[0])}};
  
  /* demux (Ty MemOut_CTf_f_Int,
       Ty Pointer_CTf_f_Int) : (memWriteOut_CTf_f_Int,MemOut_CTf_f_Int) (dconPtr_CTf_f_Int,Pointer_CTf_f_Int) > [(_167,Pointer_CTf_f_Int),
                                                                                                                 (demuxWriteResult_CTf_f_Int,Pointer_CTf_f_Int)] */
  logic [1:0] dconPtr_CTf_f_Int_onehotd;
  always_comb
    if ((memWriteOut_CTf_f_Int_d[0] && dconPtr_CTf_f_Int_d[0]))
      unique case (memWriteOut_CTf_f_Int_d[1:1])
        1'd0: dconPtr_CTf_f_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTf_f_Int_onehotd = 2'd2;
        default: dconPtr_CTf_f_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_f_Int_onehotd = 2'd0;
  assign _167_d = {dconPtr_CTf_f_Int_d[16:1],
                   dconPtr_CTf_f_Int_onehotd[0]};
  assign demuxWriteResult_CTf_f_Int_d = {dconPtr_CTf_f_Int_d[16:1],
                                         dconPtr_CTf_f_Int_onehotd[1]};
  assign dconPtr_CTf_f_Int_r = (| (dconPtr_CTf_f_Int_onehotd & {demuxWriteResult_CTf_f_Int_r,
                                                                _167_r}));
  assign memWriteOut_CTf_f_Int_r = dconPtr_CTf_f_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* mergectrl (Ty C2,
           Ty Pointer_MaskQTree) : [(m1ae3_1_argbuf,Pointer_MaskQTree),
                                    (q4aew_1_argbuf,Pointer_MaskQTree)] > (readMerge_choice_MaskQTree,C2) (readMerge_data_MaskQTree,Pointer_MaskQTree) */
  logic [1:0] m1ae3_1_argbuf_select_d;
  assign m1ae3_1_argbuf_select_d = ((| m1ae3_1_argbuf_select_q) ? m1ae3_1_argbuf_select_q :
                                    (m1ae3_1_argbuf_d[0] ? 2'd1 :
                                     (q4aew_1_argbuf_d[0] ? 2'd2 :
                                      2'd0)));
  logic [1:0] m1ae3_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae3_1_argbuf_select_q <= 2'd0;
    else
      m1ae3_1_argbuf_select_q <= (m1ae3_1_argbuf_done ? 2'd0 :
                                  m1ae3_1_argbuf_select_d);
  logic [1:0] m1ae3_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae3_1_argbuf_emit_q <= 2'd0;
    else
      m1ae3_1_argbuf_emit_q <= (m1ae3_1_argbuf_done ? 2'd0 :
                                m1ae3_1_argbuf_emit_d);
  logic [1:0] m1ae3_1_argbuf_emit_d;
  assign m1ae3_1_argbuf_emit_d = (m1ae3_1_argbuf_emit_q | ({readMerge_choice_MaskQTree_d[0],
                                                            readMerge_data_MaskQTree_d[0]} & {readMerge_choice_MaskQTree_r,
                                                                                              readMerge_data_MaskQTree_r}));
  logic m1ae3_1_argbuf_done;
  assign m1ae3_1_argbuf_done = (& m1ae3_1_argbuf_emit_d);
  assign {q4aew_1_argbuf_r,
          m1ae3_1_argbuf_r} = (m1ae3_1_argbuf_done ? m1ae3_1_argbuf_select_d :
                               2'd0);
  assign readMerge_data_MaskQTree_d = ((m1ae3_1_argbuf_select_d[0] && (! m1ae3_1_argbuf_emit_q[0])) ? m1ae3_1_argbuf_d :
                                       ((m1ae3_1_argbuf_select_d[1] && (! m1ae3_1_argbuf_emit_q[0])) ? q4aew_1_argbuf_d :
                                        {16'd0, 1'd0}));
  assign readMerge_choice_MaskQTree_d = ((m1ae3_1_argbuf_select_d[0] && (! m1ae3_1_argbuf_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((m1ae3_1_argbuf_select_d[1] && (! m1ae3_1_argbuf_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* demux (Ty C2,
       Ty MaskQTree) : (readMerge_choice_MaskQTree,C2) (destructReadOut_MaskQTree,MaskQTree) > [(readPointer_MaskQTreem1ae3_1_argbuf,MaskQTree),
                                                                                                (readPointer_MaskQTreeq4aew_1_argbuf,MaskQTree)] */
  logic [1:0] destructReadOut_MaskQTree_onehotd;
  always_comb
    if ((readMerge_choice_MaskQTree_d[0] && destructReadOut_MaskQTree_d[0]))
      unique case (readMerge_choice_MaskQTree_d[1:1])
        1'd0: destructReadOut_MaskQTree_onehotd = 2'd1;
        1'd1: destructReadOut_MaskQTree_onehotd = 2'd2;
        default: destructReadOut_MaskQTree_onehotd = 2'd0;
      endcase
    else destructReadOut_MaskQTree_onehotd = 2'd0;
  assign readPointer_MaskQTreem1ae3_1_argbuf_d = {destructReadOut_MaskQTree_d[66:1],
                                                  destructReadOut_MaskQTree_onehotd[0]};
  assign readPointer_MaskQTreeq4aew_1_argbuf_d = {destructReadOut_MaskQTree_d[66:1],
                                                  destructReadOut_MaskQTree_onehotd[1]};
  assign destructReadOut_MaskQTree_r = (| (destructReadOut_MaskQTree_onehotd & {readPointer_MaskQTreeq4aew_1_argbuf_r,
                                                                                readPointer_MaskQTreem1ae3_1_argbuf_r}));
  assign readMerge_choice_MaskQTree_r = destructReadOut_MaskQTree_r;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (readMerge_data_MaskQTree,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {readMerge_data_MaskQTree_d[16:1],
                                       readMerge_data_MaskQTree_d[0]};
  assign readMerge_data_MaskQTree_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(destructReadOut_MaskQTree,MaskQTree)] */
  assign destructReadOut_MaskQTree_d = {memReadOut_MaskQTree_d[67:2],
                                        memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = destructReadOut_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_166,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _166_d = {dconPtr_MaskQTree_d[16:1],
                   dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _166_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1a8v_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2a8w_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m3a8x_2,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnz_IntTupGo___Pointer_QTree_Intgo_6,Go),
                                                                                                                ($wnnz_IntTupGo___Pointer_QTree_IntwsjQ,Pointer_QTree_Int)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_d  = {\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [16:1],
                                                       (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_done  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_d [0],
                                                                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0]} & {\$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_r ,
                                                                                                                                                             \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r }));
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                         \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnz_IntTupGo___Pointer_QTree_Intgo_6,Go) > [(go_6_1,Go),
                                                              (go_6_2,Go)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done ;
  assign go_6_1_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted [0]));
  assign go_6_2_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted [1]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done  = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  | ({go_6_2_d[0],
                                                                                                               go_6_1_d[0]} & {go_6_2_r,
                                                                                                                               go_6_1_r}));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Intgo_6_r  ? 2'd0 :
                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_6_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_IntwsjQ,Pointer_QTree_Int) > (wsjQ_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_r ;
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_r  = ((! \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d [0]) || \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d  <= {16'd0,
                                                             1'd0};
    else
      if (\$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_r )
        \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d  <= \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_d ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf ;
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_r  = (! \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf [0]);
  assign wsjQ_1_argbuf_d = (\$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf [0] ? \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf  :
                            \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf  <= {16'd0,
                                                               1'd0};
    else
      if ((wsjQ_1_argbuf_r && \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf [0]))
        \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf  <= {16'd0,
                                                                 1'd0};
      else if (((! wsjQ_1_argbuf_r) && (! \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf [0])))
        \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_buf  <= \$wnnz_IntTupGo___Pointer_QTree_IntwsjQ_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_Int_resbuf,Int#)] > (es_6_1I#,Int) */
  assign \es_6_1I#_d  = \I#_dc ((& {\$wnnz_Int_resbuf_d [0]}), \$wnnz_Int_resbuf_d );
  assign {\$wnnz_Int_resbuf_r } = {1 {(\es_6_1I#_r  && \es_6_1I#_d [0])}};
  
  /* mergectrl (Ty C2,
           Ty TupGo___MyDTInt_Bool___Int) : [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int)] > (applyfnInt_Bool_5_choice,C2) (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) */
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d = ((| applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q :
                                                                   (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] ? 2'd1 :
                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0] ? 2'd2 :
                                                                     2'd0)));
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                                 applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                               applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q | ({applyfnInt_Bool_5_choice_d[0],
                                                                                                                          applyfnInt_Bool_5_data_d[0]} & {applyfnInt_Bool_5_choice_r,
                                                                                                                                                          applyfnInt_Bool_5_data_r}));
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  assign {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r} = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d :
                                                              2'd0);
  assign applyfnInt_Bool_5_data_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d :
                                     ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d :
                                      {32'd0, 1'd0}));
  assign applyfnInt_Bool_5_choice_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_1,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_1_bufchan_d;
  logic applyfnInt_Bool_5_1_bufchan_r;
  assign applyfnInt_Bool_5_1_r = ((! applyfnInt_Bool_5_1_bufchan_d[0]) || applyfnInt_Bool_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_1_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_1_r)
        applyfnInt_Bool_5_1_bufchan_d <= applyfnInt_Bool_5_1_d;
  MyBool_t applyfnInt_Bool_5_1_bufchan_buf;
  assign applyfnInt_Bool_5_1_bufchan_r = (! applyfnInt_Bool_5_1_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (applyfnInt_Bool_5_1_bufchan_buf[0] ? applyfnInt_Bool_5_1_bufchan_buf :
                                       applyfnInt_Bool_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && applyfnInt_Bool_5_1_bufchan_buf[0]))
        applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! applyfnInt_Bool_5_1_bufchan_buf[0])))
        applyfnInt_Bool_5_1_bufchan_buf <= applyfnInt_Bool_5_1_bufchan_d;
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_2,MyBool) > (applyfnInt_Bool_5_2_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_2_bufchan_d;
  logic applyfnInt_Bool_5_2_bufchan_r;
  assign applyfnInt_Bool_5_2_r = ((! applyfnInt_Bool_5_2_bufchan_d[0]) || applyfnInt_Bool_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_2_r)
        applyfnInt_Bool_5_2_bufchan_d <= applyfnInt_Bool_5_2_d;
  MyBool_t applyfnInt_Bool_5_2_bufchan_buf;
  assign applyfnInt_Bool_5_2_bufchan_r = (! applyfnInt_Bool_5_2_bufchan_buf[0]);
  assign applyfnInt_Bool_5_2_argbuf_d = (applyfnInt_Bool_5_2_bufchan_buf[0] ? applyfnInt_Bool_5_2_bufchan_buf :
                                         applyfnInt_Bool_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_2_argbuf_r && applyfnInt_Bool_5_2_bufchan_buf[0]))
        applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_2_argbuf_r) && (! applyfnInt_Bool_5_2_bufchan_buf[0])))
        applyfnInt_Bool_5_2_bufchan_buf <= applyfnInt_Bool_5_2_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_2_argbuf,MyBool) > [(es_6_1_1,MyBool),
                                                          (es_6_1_2,MyBool)] */
  logic [1:0] applyfnInt_Bool_5_2_argbuf_emitted;
  logic [1:0] applyfnInt_Bool_5_2_argbuf_done;
  assign es_6_1_1_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[0]))};
  assign es_6_1_2_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[1]))};
  assign applyfnInt_Bool_5_2_argbuf_done = (applyfnInt_Bool_5_2_argbuf_emitted | ({es_6_1_2_d[0],
                                                                                   es_6_1_1_d[0]} & {es_6_1_2_r,
                                                                                                     es_6_1_1_r}));
  assign applyfnInt_Bool_5_2_argbuf_r = (& applyfnInt_Bool_5_2_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_argbuf_emitted <= 2'd0;
    else
      applyfnInt_Bool_5_2_argbuf_emitted <= (applyfnInt_Bool_5_2_argbuf_r ? 2'd0 :
                                             applyfnInt_Bool_5_2_argbuf_done);
  
  /* demux (Ty C2,
       Ty MyBool) : (applyfnInt_Bool_5_choice,C2) (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > [(applyfnInt_Bool_5_1,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_2,MyBool)] */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd;
  always_comb
    if ((applyfnInt_Bool_5_choice_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[0]))
      unique case (applyfnInt_Bool_5_choice_d[1:1])
        1'd0:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd1;
        1'd1:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd2;
        default:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
      endcase
    else
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
  assign applyfnInt_Bool_5_1_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[0]};
  assign applyfnInt_Bool_5_2_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[1]};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = (| (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd & {applyfnInt_Bool_5_2_r,
                                                                                                                                                                  applyfnInt_Bool_5_1_r}));
  assign applyfnInt_Bool_5_choice_r = lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5_data_emitted;
  logic [2:0] applyfnInt_Bool_5_data_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5_data_d[32:1],
                                                              (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[2]))};
  assign applyfnInt_Bool_5_data_done = (applyfnInt_Bool_5_data_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r}));
  assign applyfnInt_Bool_5_data_r = (& applyfnInt_Bool_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_data_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_data_emitted <= (applyfnInt_Bool_5_data_r ? 3'd0 :
                                         applyfnInt_Bool_5_data_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_2_1,MyBool),
                                                        (es_2_2,MyBool),
                                                        (es_2_3,MyBool),
                                                        (es_2_4,MyBool),
                                                        (es_2_5,MyBool)] */
  logic [4:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [4:0] applyfnInt_Bool_5_resbuf_done;
  assign es_2_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_2_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_2_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign es_2_4_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[3]))};
  assign es_2_5_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[4]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_2_5_d[0],
                                                                               es_2_4_d[0],
                                                                               es_2_3_d[0],
                                                                               es_2_2_d[0],
                                                                               es_2_1_d[0]} & {es_2_5_r,
                                                                                               es_2_4_r,
                                                                                               es_2_3_r,
                                                                                               es_2_2_r,
                                                                                               es_2_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 5'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 5'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* mergectrl (Ty C3,
           Ty TupMyDTInt_Int_Int___Int___Int) : [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int)] > (applyfnInt_Int_Int_5_choice,C3) (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d = ((| applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q :
                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] ? 3'd1 :
                                                                           (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0] ? 3'd2 :
                                                                            (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0] ? 3'd4 :
                                                                             3'd0))));
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 3'd0 :
                                                                        applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 2'd0 :
                                                                      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q | ({applyfnInt_Int_Int_5_choice_d[0],
                                                                                                                                        applyfnInt_Int_Int_5_data_d[0]} & {applyfnInt_Int_Int_5_choice_r,
                                                                                                                                                                           applyfnInt_Int_Int_5_data_r}));
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  assign {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r} = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d :
                                                                     3'd0);
  assign applyfnInt_Int_Int_5_data_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d :
                                        ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d :
                                         ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d :
                                          {64'd0, 1'd0})));
  assign applyfnInt_Int_Int_5_choice_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int) > [(arg0_2_1,MyDTInt_Int_Int),
                                                                                                          (arg0_2_2,MyDTInt_Int_Int),
                                                                                                          (arg0_2_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                                               arg0_2_2_d[0],
                                                                                                                                               arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                                                 arg0_2_2_r,
                                                                                                                                                                 arg0_2_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_1,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_Int_5_1_bufchan_d;
  logic applyfnInt_Int_Int_5_1_bufchan_r;
  assign applyfnInt_Int_Int_5_1_r = ((! applyfnInt_Int_Int_5_1_bufchan_d[0]) || applyfnInt_Int_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_1_r)
        applyfnInt_Int_Int_5_1_bufchan_d <= applyfnInt_Int_Int_5_1_d;
  Int_t applyfnInt_Int_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_Int_5_1_bufchan_r = (! applyfnInt_Int_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (applyfnInt_Int_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_Int_5_1_bufchan_buf :
                                          applyfnInt_Int_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && applyfnInt_Int_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! applyfnInt_Int_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_Int_5_1_bufchan_buf <= applyfnInt_Int_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2,Int) > (applyfnInt_Int_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_bufchan_d;
  logic applyfnInt_Int_Int_5_2_bufchan_r;
  assign applyfnInt_Int_Int_5_2_r = ((! applyfnInt_Int_Int_5_2_bufchan_d[0]) || applyfnInt_Int_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_r)
        applyfnInt_Int_Int_5_2_bufchan_d <= applyfnInt_Int_Int_5_2_d;
  Int_t applyfnInt_Int_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_bufchan_r = (! applyfnInt_Int_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_2_argbuf_d = (applyfnInt_Int_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_bufchan_buf :
                                            applyfnInt_Int_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_2_argbuf_r && applyfnInt_Int_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_2_argbuf_r) && (! applyfnInt_Int_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_bufchan_buf <= applyfnInt_Int_Int_5_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_2_argbuf,Int)] > (es_3_1QVal_Int,QTree_Int) */
  assign es_3_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_2_argbuf_d[0]}), applyfnInt_Int_Int_5_2_argbuf_d);
  assign {applyfnInt_Int_Int_5_2_argbuf_r} = {1 {(es_3_1QVal_Int_r && es_3_1QVal_Int_d[0])}};
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3,Int) > (applyfnInt_Int_Int_5_3_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_bufchan_d;
  logic applyfnInt_Int_Int_5_3_bufchan_r;
  assign applyfnInt_Int_Int_5_3_r = ((! applyfnInt_Int_Int_5_3_bufchan_d[0]) || applyfnInt_Int_Int_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_r)
        applyfnInt_Int_Int_5_3_bufchan_d <= applyfnInt_Int_Int_5_3_d;
  Int_t applyfnInt_Int_Int_5_3_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_bufchan_r = (! applyfnInt_Int_Int_5_3_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_3_argbuf_d = (applyfnInt_Int_Int_5_3_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_bufchan_buf :
                                            applyfnInt_Int_Int_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_3_argbuf_r && applyfnInt_Int_Int_5_3_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_3_argbuf_r) && (! applyfnInt_Int_Int_5_3_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_bufchan_buf <= applyfnInt_Int_Int_5_3_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3_argbuf,Int) > (es_5_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_3_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_3_argbuf_r = ((! applyfnInt_Int_Int_5_3_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_3_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_argbuf_r)
        applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= applyfnInt_Int_Int_5_3_argbuf_d;
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]);
  assign es_5_1_1_argbuf_d = (applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_argbuf_bufchan_buf :
                              applyfnInt_Int_Int_5_3_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_5_1_1_argbuf_r && applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_5_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  
  /* demux (Ty C3,
       Ty Int) : (applyfnInt_Int_Int_5_choice,C3) (es_0_1_1I#_mux_mux_mux,Int) > [(applyfnInt_Int_Int_5_1,Int),
                                                                                  (applyfnInt_Int_Int_5_2,Int),
                                                                                  (applyfnInt_Int_Int_5_3,Int)] */
  logic [2:0] \es_0_1_1I#_mux_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_Int_5_choice_d[0] && \es_0_1_1I#_mux_mux_mux_d [0]))
      unique case (applyfnInt_Int_Int_5_choice_d[2:1])
        2'd0: \es_0_1_1I#_mux_mux_mux_onehotd  = 3'd1;
        2'd1: \es_0_1_1I#_mux_mux_mux_onehotd  = 3'd2;
        2'd2: \es_0_1_1I#_mux_mux_mux_onehotd  = 3'd4;
        default: \es_0_1_1I#_mux_mux_mux_onehotd  = 3'd0;
      endcase
    else \es_0_1_1I#_mux_mux_mux_onehotd  = 3'd0;
  assign applyfnInt_Int_Int_5_1_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [0]};
  assign applyfnInt_Int_Int_5_2_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [1]};
  assign applyfnInt_Int_Int_5_3_d = {\es_0_1_1I#_mux_mux_mux_d [32:1],
                                     \es_0_1_1I#_mux_mux_mux_onehotd [2]};
  assign \es_0_1_1I#_mux_mux_mux_r  = (| (\es_0_1_1I#_mux_mux_mux_onehotd  & {applyfnInt_Int_Int_5_3_r,
                                                                              applyfnInt_Int_Int_5_2_r,
                                                                              applyfnInt_Int_Int_5_1_r}));
  assign applyfnInt_Int_Int_5_choice_r = \es_0_1_1I#_mux_mux_mux_r ;
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2,MyDTInt_Int_Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_Int_5_data_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d = (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5_data_d[32:1],
                                                                     (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d = {applyfnInt_Int_Int_5_data_d[64:33],
                                                                       (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_Int_5_data_done = (applyfnInt_Int_Int_5_data_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_2_r}));
  assign applyfnInt_Int_Int_5_data_r = (& applyfnInt_Int_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5_data_emitted <= (applyfnInt_Int_Int_5_data_r ? 3'd0 :
                                            applyfnInt_Int_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > (es_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_resbuf_r = ((! applyfnInt_Int_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_resbuf_r)
        applyfnInt_Int_Int_5_resbuf_bufchan_d <= applyfnInt_Int_Int_5_resbuf_d;
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (applyfnInt_Int_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_resbuf_bufchan_buf :
                            applyfnInt_Int_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_Int_5_resbuf_bufchan_d;
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_main1,Int)] */
  assign arg0_1Dcon_main1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                               (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_main1,Int) > [(arg0_1Dcon_main1_1,Int),
                                          (arg0_1Dcon_main1_2,Int),
                                          (arg0_1Dcon_main1_3,Int),
                                          (arg0_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_1Dcon_main1_emitted;
  logic [3:0] arg0_1Dcon_main1_done;
  assign arg0_1Dcon_main1_1_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[0]))};
  assign arg0_1Dcon_main1_2_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[1]))};
  assign arg0_1Dcon_main1_3_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[2]))};
  assign arg0_1Dcon_main1_4_d = {arg0_1Dcon_main1_d[32:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[3]))};
  assign arg0_1Dcon_main1_done = (arg0_1Dcon_main1_emitted | ({arg0_1Dcon_main1_4_d[0],
                                                               arg0_1Dcon_main1_3_d[0],
                                                               arg0_1Dcon_main1_2_d[0],
                                                               arg0_1Dcon_main1_1_d[0]} & {arg0_1Dcon_main1_4_r,
                                                                                           arg0_1Dcon_main1_3_r,
                                                                                           arg0_1Dcon_main1_2_r,
                                                                                           arg0_1Dcon_main1_1_r}));
  assign arg0_1Dcon_main1_r = (& arg0_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_1Dcon_main1_emitted <= (arg0_1Dcon_main1_r ? 4'd0 :
                                   arg0_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_main1_1I#,Int) > [(xahT_destruct,Int#)] */
  assign xahT_destruct_d = {\arg0_1Dcon_main1_1I#_d [32:1],
                            \arg0_1Dcon_main1_1I#_d [0]};
  assign \arg0_1Dcon_main1_1I#_r  = xahT_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_main1_2,Int) (arg0_1Dcon_main1_1,Int) > [(arg0_1Dcon_main1_1I#,Int)] */
  assign \arg0_1Dcon_main1_1I#_d  = {arg0_1Dcon_main1_1_d[32:1],
                                     (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0])};
  assign arg0_1Dcon_main1_1_r = (\arg0_1Dcon_main1_1I#_r  && (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0]));
  assign arg0_1Dcon_main1_2_r = (\arg0_1Dcon_main1_1I#_r  && (arg0_1Dcon_main1_2_d[0] && arg0_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_main1_3,Int) (arg0_2Dcon_main1,Go) > [(arg0_1Dcon_main1_3I#,Go)] */
  assign \arg0_1Dcon_main1_3I#_d  = (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]);
  assign arg0_2Dcon_main1_r = (\arg0_1Dcon_main1_3I#_r  && (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]));
  assign arg0_1Dcon_main1_3_r = (\arg0_1Dcon_main1_3I#_r  && (arg0_1Dcon_main1_3_d[0] && arg0_2Dcon_main1_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_main1_3I#,Go) > [(arg0_1Dcon_main1_3I#_1,Go),
                                            (arg0_1Dcon_main1_3I#_2,Go),
                                            (arg0_1Dcon_main1_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_main1_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_main1_3I#_done ;
  assign \arg0_1Dcon_main1_3I#_1_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [0]));
  assign \arg0_1Dcon_main1_3I#_2_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [1]));
  assign \arg0_1Dcon_main1_3I#_3_d  = (\arg0_1Dcon_main1_3I#_d [0] && (! \arg0_1Dcon_main1_3I#_emitted [2]));
  assign \arg0_1Dcon_main1_3I#_done  = (\arg0_1Dcon_main1_3I#_emitted  | ({\arg0_1Dcon_main1_3I#_3_d [0],
                                                                           \arg0_1Dcon_main1_3I#_2_d [0],
                                                                           \arg0_1Dcon_main1_3I#_1_d [0]} & {\arg0_1Dcon_main1_3I#_3_r ,
                                                                                                             \arg0_1Dcon_main1_3I#_2_r ,
                                                                                                             \arg0_1Dcon_main1_3I#_1_r }));
  assign \arg0_1Dcon_main1_3I#_r  = (& \arg0_1Dcon_main1_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_main1_3I#_emitted  <= (\arg0_1Dcon_main1_3I#_r  ? 3'd0 :
                                         \arg0_1Dcon_main1_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_main1_3I#_1,Go) > (arg0_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_main1_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_main1_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_main1_3I#_1_r  = ((! \arg0_1Dcon_main1_3I#_1_bufchan_d [0]) || \arg0_1Dcon_main1_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_main1_3I#_1_r )
        \arg0_1Dcon_main1_3I#_1_bufchan_d  <= \arg0_1Dcon_main1_3I#_1_d ;
  Go_t \arg0_1Dcon_main1_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_main1_3I#_1_bufchan_r  = (! \arg0_1Dcon_main1_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_1Dcon_main1_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_main1_3I#_1_bufchan_buf  :
                                              \arg0_1Dcon_main1_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_main1_3I#_1_argbuf_r  && \arg0_1Dcon_main1_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_1Dcon_main1_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_main1_3I#_1_bufchan_buf  <= \arg0_1Dcon_main1_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_1Dcon_main1_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_main1_3I#_1_argbuf_0_d  = {32'd0,
                                                \arg0_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_main1_3I#_1_argbuf_r  = \arg0_1Dcon_main1_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_main1_3I#_1_argbuf_0,Int#) (xahT_destruct,Int#) > (lizzieLet1_1wild1Xt_1_Eq,Bool) */
  assign lizzieLet1_1wild1Xt_1_Eq_d = {(\arg0_1Dcon_main1_3I#_1_argbuf_0_d [32:1] == xahT_destruct_d[32:1]),
                                       (\arg0_1Dcon_main1_3I#_1_argbuf_0_d [0] && xahT_destruct_d[0])};
  assign {\arg0_1Dcon_main1_3I#_1_argbuf_0_r ,
          xahT_destruct_r} = {2 {(lizzieLet1_1wild1Xt_1_Eq_r && lizzieLet1_1wild1Xt_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_main1_3I#_2,Go) > (arg0_1Dcon_main1_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_main1_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_main1_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_main1_3I#_2_r  = ((! \arg0_1Dcon_main1_3I#_2_bufchan_d [0]) || \arg0_1Dcon_main1_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_main1_3I#_2_r )
        \arg0_1Dcon_main1_3I#_2_bufchan_d  <= \arg0_1Dcon_main1_3I#_2_d ;
  Go_t \arg0_1Dcon_main1_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_main1_3I#_2_bufchan_r  = (! \arg0_1Dcon_main1_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_main1_3I#_2_argbuf_d  = (\arg0_1Dcon_main1_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_main1_3I#_2_bufchan_buf  :
                                              \arg0_1Dcon_main1_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_main1_3I#_2_argbuf_r  && \arg0_1Dcon_main1_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_main1_3I#_2_argbuf_r ) && (! \arg0_1Dcon_main1_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_main1_3I#_2_bufchan_buf  <= \arg0_1Dcon_main1_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_main1_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_main1_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_main1_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_main1_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_main1_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_main1_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_main1_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7,Go) > [(arg0_2Dcon_main1,Go)] */
  assign arg0_2Dcon_main1_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  assign arg0_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_7_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1,Int) > [(arg0_2_1Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_2_1Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[32:1],
                                          (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_r = (\arg0_2_1Dcon_$fNumInt_$c+_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (\arg0_2_1Dcon_$fNumInt_$c+_r  && (arg0_2_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_1_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_2_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_2_2Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                          (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_2_2Dcon_$fNumInt_$c+_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_2_2_r = (\arg0_2_2Dcon_$fNumInt_$c+_r  && (arg0_2_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_1,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_2,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_3,Int),
                                                   (arg0_2_2Dcon_$fNumInt_$c+_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_done ;
  assign \arg0_2_2Dcon_$fNumInt_$c+_1_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_2_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_4_d  = {\arg0_2_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_2_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_done  = (\arg0_2_2Dcon_$fNumInt_$c+_emitted  | ({\arg0_2_2Dcon_$fNumInt_$c+_4_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_3_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_2_d [0],
                                                                                     \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$c+_4_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_3_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_2_r ,
                                                                                                                            \arg0_2_2Dcon_$fNumInt_$c+_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$c+_r  = (& \arg0_2_2Dcon_$fNumInt_$c+_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_2Dcon_$fNumInt_$c+_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$c+_emitted  <= (\arg0_2_2Dcon_$fNumInt_$c+_r  ? 4'd0 :
                                              \arg0_2_2Dcon_$fNumInt_$c+_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c+_1I#,Int) > [(xa1lV_destruct,Int#)] */
  assign xa1lV_destruct_d = {\arg0_2_2Dcon_$fNumInt_$c+_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$c+_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$c+_1I#_r  = xa1lV_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_2,Int) (arg0_2_2Dcon_$fNumInt_$c+_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$c+_1_d [32:1],
                                              (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$c+_1_r  = (\arg0_2_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_2_r  = (\arg0_2_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3,Int) (arg0_2_1Dcon_$fNumInt_$c+,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_d  = {\arg0_2_1Dcon_$fNumInt_$c+_d [32:1],
                                              (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0])};
  assign \arg0_2_1Dcon_$fNumInt_$c+_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_2_1Dcon_$fNumInt_$c+_d [0]));
  
  /* fork (Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_1,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_2,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_3,Int),
                                                       (arg0_2_2Dcon_$fNumInt_$c+_3I#_4,Int)] */
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted ;
  logic [3:0] \arg0_2_2Dcon_$fNumInt_$c+_3I#_done ;
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [0]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [1]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [2]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_2_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted [3]))};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_done  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  | ({\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0],
                                                                                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]} & {\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r ,
                                                                                                                                        \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r }));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_r  = (& \arg0_2_2Dcon_$fNumInt_$c+_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  <= 4'd0;
    else
      \arg0_2_2Dcon_$fNumInt_$c+_3I#_emitted  <= (\arg0_2_2Dcon_$fNumInt_$c+_3I#_r  ? 4'd0 :
                                                  \arg0_2_2Dcon_$fNumInt_$c+_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#,Int) > [(ya1lW_destruct,Int#)] */
  assign ya1lW_destruct_d = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d [32:1],
                             \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d [0]};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  = ya1lW_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_2,Int) (arg0_2_2Dcon_$fNumInt_$c+_3I#_1,Int) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#,Int)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_d  = {\arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0])};
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_2_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_2_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_3,Int) (xa1lV_destruct,Int#) > [(arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#,Int#)] */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d  = {xa1lV_destruct_d[32:1],
                                                  (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0])};
  assign xa1lV_destruct_r = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3_r  = (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  
  /* op_add (Ty Int#) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#,Int#) (ya1lW_destruct,Int#) > (arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#) */
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d  = {(\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d [32:1] + ya1lW_destruct_d[32:1]),
                                                                 (\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_d [0] && ya1lW_destruct_d[0])};
  assign {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_r ,
          ya1lW_destruct_r} = {2 {(\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r  && \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0]}), \arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d );
  assign {\arg0_2_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r } = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_3I#_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_3I#_4_r  = (\es_0_1_1I#_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_1_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_2Dcon_$fNumInt_$c+_4,Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  assign \arg0_2_2Dcon_$fNumInt_$c+_4_r  = (\es_0_1_1I#_mux_mux_r  && (\arg0_2_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int_Int) [(es_0_1_1I#_mux_mux,Int)] > (es_0_1_1I#_mux_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_mux_d  = {\es_0_1_1I#_mux_mux_d [32:1],
                                       (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0])};
  assign \es_0_1_1I#_mux_mux_r  = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  assign arg0_2_3_r = (\es_0_1_1I#_mux_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) > [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8,Go),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1,Pointer_QTree_Int),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] */
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted;
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done;
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[0]));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[16:1],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[1]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[32:17],
                                                                                (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[2]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted | ({call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]} & {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_r,
                                                                                                                                                                                                                                        call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r}));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r = (& call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= 3'd0;
    else
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r ? 3'd0 :
                                                                                  call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_Int_goConst,Go) > (call_$wnnz_Int_initBufi,Go) */
  Go_t call_$wnnz_Int_goConst_buf;
  assign call_$wnnz_Int_goConst_r = (! call_$wnnz_Int_goConst_buf[0]);
  assign call_$wnnz_Int_initBufi_d = (call_$wnnz_Int_goConst_buf[0] ? call_$wnnz_Int_goConst_buf :
                                      call_$wnnz_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_Int_initBufi_r && call_$wnnz_Int_goConst_buf[0]))
        call_$wnnz_Int_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_Int_initBufi_r) && (! call_$wnnz_Int_goConst_buf[0])))
        call_$wnnz_Int_goConst_buf <= call_$wnnz_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_Int_goMux1,Go),
                           (lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf,Go),
                           (lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf,Go),
                           (lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_8_goMux_choice,C5) (go_8_goMux_data,Go) */
  logic [4:0] call_$wnnz_Int_goMux1_select_d;
  assign call_$wnnz_Int_goMux1_select_d = ((| call_$wnnz_Int_goMux1_select_q) ? call_$wnnz_Int_goMux1_select_q :
                                           (call_$wnnz_Int_goMux1_d[0] ? 5'd1 :
                                            (lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_d[0] ? 5'd2 :
                                             (lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_d[0] ? 5'd4 :
                                              (lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_d[0] ? 5'd8 :
                                               (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                5'd0))))));
  logic [4:0] call_$wnnz_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_Int_goMux1_select_q <= (call_$wnnz_Int_goMux1_done ? 5'd0 :
                                         call_$wnnz_Int_goMux1_select_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_Int_goMux1_emit_q <= (call_$wnnz_Int_goMux1_done ? 2'd0 :
                                       call_$wnnz_Int_goMux1_emit_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_d;
  assign call_$wnnz_Int_goMux1_emit_d = (call_$wnnz_Int_goMux1_emit_q | ({go_8_goMux_choice_d[0],
                                                                          go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                   go_8_goMux_data_r}));
  logic call_$wnnz_Int_goMux1_done;
  assign call_$wnnz_Int_goMux1_done = (& call_$wnnz_Int_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_r,
          lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_r,
          lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_r,
          call_$wnnz_Int_goMux1_r} = (call_$wnnz_Int_goMux1_done ? call_$wnnz_Int_goMux1_select_d :
                                      5'd0);
  assign go_8_goMux_data_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? call_$wnnz_Int_goMux1_d :
                              ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_d :
                               ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_d :
                                ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_d :
                                 ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_8_goMux_choice_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_Int_initBuf,Go) > [(call_$wnnz_Int_unlockFork1,Go),
                                              (call_$wnnz_Int_unlockFork2,Go),
                                              (call_$wnnz_Int_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_Int_initBuf_emitted;
  logic [2:0] call_$wnnz_Int_initBuf_done;
  assign call_$wnnz_Int_unlockFork1_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[0]));
  assign call_$wnnz_Int_unlockFork2_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[1]));
  assign call_$wnnz_Int_unlockFork3_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[2]));
  assign call_$wnnz_Int_initBuf_done = (call_$wnnz_Int_initBuf_emitted | ({call_$wnnz_Int_unlockFork3_d[0],
                                                                           call_$wnnz_Int_unlockFork2_d[0],
                                                                           call_$wnnz_Int_unlockFork1_d[0]} & {call_$wnnz_Int_unlockFork3_r,
                                                                                                               call_$wnnz_Int_unlockFork2_r,
                                                                                                               call_$wnnz_Int_unlockFork1_r}));
  assign call_$wnnz_Int_initBuf_r = (& call_$wnnz_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_Int_initBuf_emitted <= (call_$wnnz_Int_initBuf_r ? 3'd0 :
                                         call_$wnnz_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_Int_initBufi,Go) > (call_$wnnz_Int_initBuf,Go) */
  assign call_$wnnz_Int_initBufi_r = ((! call_$wnnz_Int_initBuf_d[0]) || call_$wnnz_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_Int_initBufi_r)
        call_$wnnz_Int_initBuf_d <= call_$wnnz_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_Int_unlockFork1,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8,Go)] > (call_$wnnz_Int_goMux1,Go) */
  assign call_$wnnz_Int_goMux1_d = (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]);
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]));
  assign call_$wnnz_Int_unlockFork1_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_8_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_Int_unlockFork2,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1,Pointer_QTree_Int)] > (call_$wnnz_Int_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_Int_goMux2_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d[0]));
  assign call_$wnnz_Int_unlockFork2_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwsjQ_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz_Int) : (call_$wnnz_Int_unlockFork3,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] > (call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int) */
  assign call_$wnnz_Int_goMux3_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[16:1],
                                    (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  assign call_$wnnz_Int_unlockFork3_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int) : (call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int) > [(call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9,Go),
                                                                                                                                                                                                                                                                                                                   (call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                                                                   (call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                   (call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [3:0] \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted ;
  logic [3:0] \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_done ;
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d  = (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [0] && (! \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted [0]));
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [16:1],
                                                                                                                                       (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [0] && (! \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted [1]))};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [32:17],
                                                                                                                                        (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [0] && (! \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted [2]))};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [48:33],
                                                                                                                                        (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [0] && (! \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted [3]))};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_done  = (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted  | ({\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d [0],
                                                                                                                                                                                                                                                                         \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d [0],
                                                                                                                                                                                                                                                                         \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d [0],
                                                                                                                                                                                                                                                                         \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d [0]} & {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                          \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_r ,
                                                                                                                                                                                                                                                                                                                                                                                                          \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_r ,
                                                                                                                                                                                                                                                                                                                                                                                                          \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_r }));
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_r  = (& \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted  <= 4'd0;
    else
      \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_emitted  <= (\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_r  ? 4'd0 :
                                                                                                                                        \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_done );
  
  /* rbuf (Ty Go) : (call_f'''''''''_f'''''''''_Int_goConst,Go) > (call_f'''''''''_f'''''''''_Int_initBufi,Go) */
  Go_t \call_f'''''''''_f'''''''''_Int_goConst_buf ;
  assign \call_f'''''''''_f'''''''''_Int_goConst_r  = (! \call_f'''''''''_f'''''''''_Int_goConst_buf [0]);
  assign \call_f'''''''''_f'''''''''_Int_initBufi_d  = (\call_f'''''''''_f'''''''''_Int_goConst_buf [0] ? \call_f'''''''''_f'''''''''_Int_goConst_buf  :
                                                        \call_f'''''''''_f'''''''''_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_f'''''''''_f'''''''''_Int_initBufi_r  && \call_f'''''''''_f'''''''''_Int_goConst_buf [0]))
        \call_f'''''''''_f'''''''''_Int_goConst_buf  <= 1'd0;
      else if (((! \call_f'''''''''_f'''''''''_Int_initBufi_r ) && (! \call_f'''''''''_f'''''''''_Int_goConst_buf [0])))
        \call_f'''''''''_f'''''''''_Int_goConst_buf  <= \call_f'''''''''_f'''''''''_Int_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_f'''''''''_f'''''''''_Int_goMux1,Go),
                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf,Go),
                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf,Go),
                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf,Go),
                     (lizzieLet6_4MQNode_3QNode_Int_1_argbuf,Go)] > (go_9_goMux_choice,C5) (go_9_goMux_data,Go) */
  logic [4:0] \call_f'''''''''_f'''''''''_Int_goMux1_select_d ;
  assign \call_f'''''''''_f'''''''''_Int_goMux1_select_d  = ((| \call_f'''''''''_f'''''''''_Int_goMux1_select_q ) ? \call_f'''''''''_f'''''''''_Int_goMux1_select_q  :
                                                             (\call_f'''''''''_f'''''''''_Int_goMux1_d [0] ? 5'd1 :
                                                              (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_d [0] ? 5'd2 :
                                                               (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_d [0] ? 5'd4 :
                                                                (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_d [0] ? 5'd8 :
                                                                 (lizzieLet6_4MQNode_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                                  5'd0))))));
  logic [4:0] \call_f'''''''''_f'''''''''_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Int_goMux1_select_q  <= 5'd0;
    else
      \call_f'''''''''_f'''''''''_Int_goMux1_select_q  <= (\call_f'''''''''_f'''''''''_Int_goMux1_done  ? 5'd0 :
                                                           \call_f'''''''''_f'''''''''_Int_goMux1_select_d );
  logic [1:0] \call_f'''''''''_f'''''''''_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_f'''''''''_f'''''''''_Int_goMux1_emit_q  <= (\call_f'''''''''_f'''''''''_Int_goMux1_done  ? 2'd0 :
                                                         \call_f'''''''''_f'''''''''_Int_goMux1_emit_d );
  logic [1:0] \call_f'''''''''_f'''''''''_Int_goMux1_emit_d ;
  assign \call_f'''''''''_f'''''''''_Int_goMux1_emit_d  = (\call_f'''''''''_f'''''''''_Int_goMux1_emit_q  | ({go_9_goMux_choice_d[0],
                                                                                                              go_9_goMux_data_d[0]} & {go_9_goMux_choice_r,
                                                                                                                                       go_9_goMux_data_r}));
  logic \call_f'''''''''_f'''''''''_Int_goMux1_done ;
  assign \call_f'''''''''_f'''''''''_Int_goMux1_done  = (& \call_f'''''''''_f'''''''''_Int_goMux1_emit_d );
  assign {lizzieLet6_4MQNode_3QNode_Int_1_argbuf_r,
          \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_r ,
          \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_r ,
          \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_r ,
          \call_f'''''''''_f'''''''''_Int_goMux1_r } = (\call_f'''''''''_f'''''''''_Int_goMux1_done  ? \call_f'''''''''_f'''''''''_Int_goMux1_select_d  :
                                                        5'd0);
  assign go_9_goMux_data_d = ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [0] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [0])) ? \call_f'''''''''_f'''''''''_Int_goMux1_d  :
                              ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [1] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_d  :
                               ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [2] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_d  :
                                ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [3] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [0])) ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_d  :
                                 ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [4] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [0])) ? lizzieLet6_4MQNode_3QNode_Int_1_argbuf_d :
                                  1'd0)))));
  assign go_9_goMux_choice_d = ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [0] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [1] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [2] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [3] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_f'''''''''_f'''''''''_Int_goMux1_select_d [4] && (! \call_f'''''''''_f'''''''''_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f'''''''''_f'''''''''_Int_initBuf,Go) > [(call_f'''''''''_f'''''''''_Int_unlockFork1,Go),
                                                              (call_f'''''''''_f'''''''''_Int_unlockFork2,Go),
                                                              (call_f'''''''''_f'''''''''_Int_unlockFork3,Go),
                                                              (call_f'''''''''_f'''''''''_Int_unlockFork4,Go)] */
  logic [3:0] \call_f'''''''''_f'''''''''_Int_initBuf_emitted ;
  logic [3:0] \call_f'''''''''_f'''''''''_Int_initBuf_done ;
  assign \call_f'''''''''_f'''''''''_Int_unlockFork1_d  = (\call_f'''''''''_f'''''''''_Int_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Int_initBuf_emitted [0]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork2_d  = (\call_f'''''''''_f'''''''''_Int_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Int_initBuf_emitted [1]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork3_d  = (\call_f'''''''''_f'''''''''_Int_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Int_initBuf_emitted [2]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork4_d  = (\call_f'''''''''_f'''''''''_Int_initBuf_d [0] && (! \call_f'''''''''_f'''''''''_Int_initBuf_emitted [3]));
  assign \call_f'''''''''_f'''''''''_Int_initBuf_done  = (\call_f'''''''''_f'''''''''_Int_initBuf_emitted  | ({\call_f'''''''''_f'''''''''_Int_unlockFork4_d [0],
                                                                                                               \call_f'''''''''_f'''''''''_Int_unlockFork3_d [0],
                                                                                                               \call_f'''''''''_f'''''''''_Int_unlockFork2_d [0],
                                                                                                               \call_f'''''''''_f'''''''''_Int_unlockFork1_d [0]} & {\call_f'''''''''_f'''''''''_Int_unlockFork4_r ,
                                                                                                                                                                     \call_f'''''''''_f'''''''''_Int_unlockFork3_r ,
                                                                                                                                                                     \call_f'''''''''_f'''''''''_Int_unlockFork2_r ,
                                                                                                                                                                     \call_f'''''''''_f'''''''''_Int_unlockFork1_r }));
  assign \call_f'''''''''_f'''''''''_Int_initBuf_r  = (& \call_f'''''''''_f'''''''''_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Int_initBuf_emitted  <= 4'd0;
    else
      \call_f'''''''''_f'''''''''_Int_initBuf_emitted  <= (\call_f'''''''''_f'''''''''_Int_initBuf_r  ? 4'd0 :
                                                           \call_f'''''''''_f'''''''''_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f'''''''''_f'''''''''_Int_initBufi,Go) > (call_f'''''''''_f'''''''''_Int_initBuf,Go) */
  assign \call_f'''''''''_f'''''''''_Int_initBufi_r  = ((! \call_f'''''''''_f'''''''''_Int_initBuf_d [0]) || \call_f'''''''''_f'''''''''_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'''''''''_f'''''''''_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f'''''''''_f'''''''''_Int_initBufi_r )
        \call_f'''''''''_f'''''''''_Int_initBuf_d  <= \call_f'''''''''_f'''''''''_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f'''''''''_f'''''''''_Int_unlockFork1,Go) [(call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9,Go)] > (call_f'''''''''_f'''''''''_Int_goMux1,Go) */
  assign \call_f'''''''''_f'''''''''_Int_goMux1_d  = (\call_f'''''''''_f'''''''''_Int_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d [0]);
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_r  = (\call_f'''''''''_f'''''''''_Int_goMux1_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d [0]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork1_r  = (\call_f'''''''''_f'''''''''_Int_goMux1_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork1_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intgo_9_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_f'''''''''_f'''''''''_Int_unlockFork2,Go) [(call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew,Pointer_MaskQTree)] > (call_f'''''''''_f'''''''''_Int_goMux2,Pointer_MaskQTree) */
  assign \call_f'''''''''_f'''''''''_Int_goMux2_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d [16:1],
                                                      (\call_f'''''''''_f'''''''''_Int_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d [0])};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_r  = (\call_f'''''''''_f'''''''''_Int_goMux2_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d [0]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork2_r  = (\call_f'''''''''_f'''''''''_Int_goMux2_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork2_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4aew_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f'''''''''_f'''''''''_Int_unlockFork3,Go) [(call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex,Pointer_QTree_Int)] > (call_f'''''''''_f'''''''''_Int_goMux3,Pointer_QTree_Int) */
  assign \call_f'''''''''_f'''''''''_Int_goMux3_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d [16:1],
                                                      (\call_f'''''''''_f'''''''''_Int_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d [0])};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_r  = (\call_f'''''''''_f'''''''''_Int_goMux3_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d [0]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork3_r  = (\call_f'''''''''_f'''''''''_Int_goMux3_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork3_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intq4'aex_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf'''''''''_f'''''''''_Int) : (call_f'''''''''_f'''''''''_Int_unlockFork4,Go) [(call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1,Pointer_CTf'''''''''_f'''''''''_Int)] > (call_f'''''''''_f'''''''''_Int_goMux4,Pointer_CTf'''''''''_f'''''''''_Int) */
  assign \call_f'''''''''_f'''''''''_Int_goMux4_d  = {\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d [16:1],
                                                      (\call_f'''''''''_f'''''''''_Int_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d [0])};
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_r  = (\call_f'''''''''_f'''''''''_Int_goMux4_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d [0]));
  assign \call_f'''''''''_f'''''''''_Int_unlockFork4_r  = (\call_f'''''''''_f'''''''''_Int_goMux4_r  && (\call_f'''''''''_f'''''''''_Int_unlockFork4_d [0] && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Intsc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int) : (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int) > [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10,Go),
                                                                                                                                                                                                                                                                                                                                                      (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                      (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                      (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                      (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                      (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2,Pointer_CTf'_f'_Int)] */
  logic [5:0] \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted ;
  logic [5:0] \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_done ;
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d  = (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [0]));
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [16:1],
                                                                                                                                        (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [1]))};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [32:17],
                                                                                                                                        (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [2]))};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d  = (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [3]));
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d  = (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [4]));
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [48:33],
                                                                                                                                         (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0] && (! \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted [5]))};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_done  = (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted  | ({\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d [0],
                                                                                                                                                                                                                                                                           \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d [0],
                                                                                                                                                                                                                                                                           \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d [0],
                                                                                                                                                                                                                                                                           \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d [0],
                                                                                                                                                                                                                                                                           \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d [0],
                                                                                                                                                                                                                                                                           \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d [0]} & {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_r }));
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_r  = (& \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted  <= 6'd0;
    else
      \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_emitted  <= (\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_r  ? 6'd0 :
                                                                                                                                         \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_done );
  
  /* rbuf (Ty Go) : (call_f'_f'_Int_goConst,Go) > (call_f'_f'_Int_initBufi,Go) */
  Go_t \call_f'_f'_Int_goConst_buf ;
  assign \call_f'_f'_Int_goConst_r  = (! \call_f'_f'_Int_goConst_buf [0]);
  assign \call_f'_f'_Int_initBufi_d  = (\call_f'_f'_Int_goConst_buf [0] ? \call_f'_f'_Int_goConst_buf  :
                                        \call_f'_f'_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_f'_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_f'_f'_Int_initBufi_r  && \call_f'_f'_Int_goConst_buf [0]))
        \call_f'_f'_Int_goConst_buf  <= 1'd0;
      else if (((! \call_f'_f'_Int_initBufi_r ) && (! \call_f'_f'_Int_goConst_buf [0])))
        \call_f'_f'_Int_goConst_buf  <= \call_f'_f'_Int_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f'_f'_Int_goMux1,Go),
                           (lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf,Go),
                           (lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf,Go),
                           (lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf,Go),
                           (lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_10_goMux_choice,C5) (go_10_goMux_data,Go) */
  logic [4:0] \call_f'_f'_Int_goMux1_select_d ;
  assign \call_f'_f'_Int_goMux1_select_d  = ((| \call_f'_f'_Int_goMux1_select_q ) ? \call_f'_f'_Int_goMux1_select_q  :
                                             (\call_f'_f'_Int_goMux1_d [0] ? 5'd1 :
                                              (\lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_d [0] ? 5'd2 :
                                               (\lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_d [0] ? 5'd4 :
                                                (\lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_d [0] ? 5'd8 :
                                                 (lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                  5'd0))))));
  logic [4:0] \call_f'_f'_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_f'_Int_goMux1_select_q  <= 5'd0;
    else
      \call_f'_f'_Int_goMux1_select_q  <= (\call_f'_f'_Int_goMux1_done  ? 5'd0 :
                                           \call_f'_f'_Int_goMux1_select_d );
  logic [1:0] \call_f'_f'_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_f'_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_f'_f'_Int_goMux1_emit_q  <= (\call_f'_f'_Int_goMux1_done  ? 2'd0 :
                                         \call_f'_f'_Int_goMux1_emit_d );
  logic [1:0] \call_f'_f'_Int_goMux1_emit_d ;
  assign \call_f'_f'_Int_goMux1_emit_d  = (\call_f'_f'_Int_goMux1_emit_q  | ({go_10_goMux_choice_d[0],
                                                                              go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                        go_10_goMux_data_r}));
  logic \call_f'_f'_Int_goMux1_done ;
  assign \call_f'_f'_Int_goMux1_done  = (& \call_f'_f'_Int_goMux1_emit_d );
  assign {lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_r,
          \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_r ,
          \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_r ,
          \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_r ,
          \call_f'_f'_Int_goMux1_r } = (\call_f'_f'_Int_goMux1_done  ? \call_f'_f'_Int_goMux1_select_d  :
                                        5'd0);
  assign go_10_goMux_data_d = ((\call_f'_f'_Int_goMux1_select_d [0] && (! \call_f'_f'_Int_goMux1_emit_q [0])) ? \call_f'_f'_Int_goMux1_d  :
                               ((\call_f'_f'_Int_goMux1_select_d [1] && (! \call_f'_f'_Int_goMux1_emit_q [0])) ? \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_d  :
                                ((\call_f'_f'_Int_goMux1_select_d [2] && (! \call_f'_f'_Int_goMux1_emit_q [0])) ? \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_d  :
                                 ((\call_f'_f'_Int_goMux1_select_d [3] && (! \call_f'_f'_Int_goMux1_emit_q [0])) ? \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_d  :
                                  ((\call_f'_f'_Int_goMux1_select_d [4] && (! \call_f'_f'_Int_goMux1_emit_q [0])) ? lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_10_goMux_choice_d = ((\call_f'_f'_Int_goMux1_select_d [0] && (! \call_f'_f'_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_f'_f'_Int_goMux1_select_d [1] && (! \call_f'_f'_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_f'_f'_Int_goMux1_select_d [2] && (! \call_f'_f'_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_f'_f'_Int_goMux1_select_d [3] && (! \call_f'_f'_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_f'_f'_Int_goMux1_select_d [4] && (! \call_f'_f'_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f'_f'_Int_initBuf,Go) > [(call_f'_f'_Int_unlockFork1,Go),
                                              (call_f'_f'_Int_unlockFork2,Go),
                                              (call_f'_f'_Int_unlockFork3,Go),
                                              (call_f'_f'_Int_unlockFork4,Go),
                                              (call_f'_f'_Int_unlockFork5,Go),
                                              (call_f'_f'_Int_unlockFork6,Go)] */
  logic [5:0] \call_f'_f'_Int_initBuf_emitted ;
  logic [5:0] \call_f'_f'_Int_initBuf_done ;
  assign \call_f'_f'_Int_unlockFork1_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [0]));
  assign \call_f'_f'_Int_unlockFork2_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [1]));
  assign \call_f'_f'_Int_unlockFork3_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [2]));
  assign \call_f'_f'_Int_unlockFork4_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [3]));
  assign \call_f'_f'_Int_unlockFork5_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [4]));
  assign \call_f'_f'_Int_unlockFork6_d  = (\call_f'_f'_Int_initBuf_d [0] && (! \call_f'_f'_Int_initBuf_emitted [5]));
  assign \call_f'_f'_Int_initBuf_done  = (\call_f'_f'_Int_initBuf_emitted  | ({\call_f'_f'_Int_unlockFork6_d [0],
                                                                               \call_f'_f'_Int_unlockFork5_d [0],
                                                                               \call_f'_f'_Int_unlockFork4_d [0],
                                                                               \call_f'_f'_Int_unlockFork3_d [0],
                                                                               \call_f'_f'_Int_unlockFork2_d [0],
                                                                               \call_f'_f'_Int_unlockFork1_d [0]} & {\call_f'_f'_Int_unlockFork6_r ,
                                                                                                                     \call_f'_f'_Int_unlockFork5_r ,
                                                                                                                     \call_f'_f'_Int_unlockFork4_r ,
                                                                                                                     \call_f'_f'_Int_unlockFork3_r ,
                                                                                                                     \call_f'_f'_Int_unlockFork2_r ,
                                                                                                                     \call_f'_f'_Int_unlockFork1_r }));
  assign \call_f'_f'_Int_initBuf_r  = (& \call_f'_f'_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_f'_Int_initBuf_emitted  <= 6'd0;
    else
      \call_f'_f'_Int_initBuf_emitted  <= (\call_f'_f'_Int_initBuf_r  ? 6'd0 :
                                           \call_f'_f'_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f'_f'_Int_initBufi,Go) > (call_f'_f'_Int_initBuf,Go) */
  assign \call_f'_f'_Int_initBufi_r  = ((! \call_f'_f'_Int_initBuf_d [0]) || \call_f'_f'_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_f'_f'_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f'_f'_Int_initBufi_r )
        \call_f'_f'_Int_initBuf_d  <= \call_f'_f'_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f'_f'_Int_unlockFork1,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10,Go)] > (call_f'_f'_Int_goMux1,Go) */
  assign \call_f'_f'_Int_goMux1_d  = (\call_f'_f'_Int_unlockFork1_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d [0]);
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_r  = (\call_f'_f'_Int_goMux1_r  && (\call_f'_f'_Int_unlockFork1_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d [0]));
  assign \call_f'_f'_Int_unlockFork1_r  = (\call_f'_f'_Int_goMux1_r  && (\call_f'_f'_Int_unlockFork1_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intgo_10_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f'_f'_Int_unlockFork2,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH,Pointer_QTree_Int)] > (call_f'_f'_Int_goMux2,Pointer_QTree_Int) */
  assign \call_f'_f'_Int_goMux2_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d [16:1],
                                      (\call_f'_f'_Int_unlockFork2_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d [0])};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_r  = (\call_f'_f'_Int_goMux2_r  && (\call_f'_f'_Int_unlockFork2_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d [0]));
  assign \call_f'_f'_Int_unlockFork2_r  = (\call_f'_f'_Int_goMux2_r  && (\call_f'_f'_Int_unlockFork2_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm2aeH_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f'_f'_Int_unlockFork3,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI,Pointer_QTree_Int)] > (call_f'_f'_Int_goMux3,Pointer_QTree_Int) */
  assign \call_f'_f'_Int_goMux3_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d [16:1],
                                      (\call_f'_f'_Int_unlockFork3_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d [0])};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_r  = (\call_f'_f'_Int_goMux3_r  && (\call_f'_f'_Int_unlockFork3_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d [0]));
  assign \call_f'_f'_Int_unlockFork3_r  = (\call_f'_f'_Int_goMux3_r  && (\call_f'_f'_Int_unlockFork3_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intm3aeI_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f'_f'_Int_unlockFork4,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ,MyDTInt_Bool)] > (call_f'_f'_Int_goMux4,MyDTInt_Bool) */
  assign \call_f'_f'_Int_goMux4_d  = (\call_f'_f'_Int_unlockFork4_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d [0]);
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_r  = (\call_f'_f'_Int_goMux4_r  && (\call_f'_f'_Int_unlockFork4_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d [0]));
  assign \call_f'_f'_Int_unlockFork4_r  = (\call_f'_f'_Int_goMux4_r  && (\call_f'_f'_Int_unlockFork4_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intis_zaeJ_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f'_f'_Int_unlockFork5,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK,MyDTInt_Int_Int)] > (call_f'_f'_Int_goMux5,MyDTInt_Int_Int) */
  assign \call_f'_f'_Int_goMux5_d  = (\call_f'_f'_Int_unlockFork5_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d [0]);
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_r  = (\call_f'_f'_Int_goMux5_r  && (\call_f'_f'_Int_unlockFork5_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d [0]));
  assign \call_f'_f'_Int_unlockFork5_r  = (\call_f'_f'_Int_goMux5_r  && (\call_f'_f'_Int_unlockFork5_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intop_addaeK_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf'_f'_Int) : (call_f'_f'_Int_unlockFork6,Go) [(call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2,Pointer_CTf'_f'_Int)] > (call_f'_f'_Int_goMux6,Pointer_CTf'_f'_Int) */
  assign \call_f'_f'_Int_goMux6_d  = {\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d [16:1],
                                      (\call_f'_f'_Int_unlockFork6_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d [0])};
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_r  = (\call_f'_f'_Int_goMux6_r  && (\call_f'_f'_Int_unlockFork6_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d [0]));
  assign \call_f'_f'_Int_unlockFork6_r  = (\call_f'_f'_Int_goMux6_r  && (\call_f'_f'_Int_unlockFork6_d [0] && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Intsc_0_2_d [0]));
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) : (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) > [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11,Go),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                          (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3,Pointer_CTf_f_Int)] */
  logic [6:0] call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted;
  logic [6:0] call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done;
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d = (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[0]));
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[16:1],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[1]))};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[32:17],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[2]))};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[48:33],
                                                                                                                                                      (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[3]))};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d = (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[4]));
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d = (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[5]));
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[64:49],
                                                                                                                                                       (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0] && (! call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted[6]))};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done = (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted | ({call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d[0],
                                                                                                                                                                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d[0]} & {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                        call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_r}));
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r = (& call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted <= 7'd0;
    else
      call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_emitted <= (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r ? 7'd0 :
                                                                                                                                                       call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_done);
  
  /* rbuf (Ty Go) : (call_f_f_Int_goConst,Go) > (call_f_f_Int_initBufi,Go) */
  Go_t call_f_f_Int_goConst_buf;
  assign call_f_f_Int_goConst_r = (! call_f_f_Int_goConst_buf[0]);
  assign call_f_f_Int_initBufi_d = (call_f_f_Int_goConst_buf[0] ? call_f_f_Int_goConst_buf :
                                    call_f_f_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goConst_buf <= 1'd0;
    else
      if ((call_f_f_Int_initBufi_r && call_f_f_Int_goConst_buf[0]))
        call_f_f_Int_goConst_buf <= 1'd0;
      else if (((! call_f_f_Int_initBufi_r) && (! call_f_f_Int_goConst_buf[0])))
        call_f_f_Int_goConst_buf <= call_f_f_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_f_Int_goMux1,Go),
                           (lizzieLet60_3Lcall_f_f_Int3_1_argbuf,Go),
                           (lizzieLet60_3Lcall_f_f_Int2_1_argbuf,Go),
                           (lizzieLet60_3Lcall_f_f_Int1_1_argbuf,Go),
                           (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] call_f_f_Int_goMux1_select_d;
  assign call_f_f_Int_goMux1_select_d = ((| call_f_f_Int_goMux1_select_q) ? call_f_f_Int_goMux1_select_q :
                                         (call_f_f_Int_goMux1_d[0] ? 5'd1 :
                                          (lizzieLet60_3Lcall_f_f_Int3_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet60_3Lcall_f_f_Int2_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet60_3Lcall_f_f_Int1_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] call_f_f_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goMux1_select_q <= 5'd0;
    else
      call_f_f_Int_goMux1_select_q <= (call_f_f_Int_goMux1_done ? 5'd0 :
                                       call_f_f_Int_goMux1_select_d);
  logic [1:0] call_f_f_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_goMux1_emit_q <= 2'd0;
    else
      call_f_f_Int_goMux1_emit_q <= (call_f_f_Int_goMux1_done ? 2'd0 :
                                     call_f_f_Int_goMux1_emit_d);
  logic [1:0] call_f_f_Int_goMux1_emit_d;
  assign call_f_f_Int_goMux1_emit_d = (call_f_f_Int_goMux1_emit_q | ({go_11_goMux_choice_d[0],
                                                                      go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                go_11_goMux_data_r}));
  logic call_f_f_Int_goMux1_done;
  assign call_f_f_Int_goMux1_done = (& call_f_f_Int_goMux1_emit_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_r,
          lizzieLet60_3Lcall_f_f_Int1_1_argbuf_r,
          lizzieLet60_3Lcall_f_f_Int2_1_argbuf_r,
          lizzieLet60_3Lcall_f_f_Int3_1_argbuf_r,
          call_f_f_Int_goMux1_r} = (call_f_f_Int_goMux1_done ? call_f_f_Int_goMux1_select_d :
                                    5'd0);
  assign go_11_goMux_data_d = ((call_f_f_Int_goMux1_select_d[0] && (! call_f_f_Int_goMux1_emit_q[0])) ? call_f_f_Int_goMux1_d :
                               ((call_f_f_Int_goMux1_select_d[1] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f_f_Int3_1_argbuf_d :
                                ((call_f_f_Int_goMux1_select_d[2] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f_f_Int2_1_argbuf_d :
                                 ((call_f_f_Int_goMux1_select_d[3] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet60_3Lcall_f_f_Int1_1_argbuf_d :
                                  ((call_f_f_Int_goMux1_select_d[4] && (! call_f_f_Int_goMux1_emit_q[0])) ? lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((call_f_f_Int_goMux1_select_d[0] && (! call_f_f_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_f_f_Int_goMux1_select_d[1] && (! call_f_f_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_f_f_Int_goMux1_select_d[2] && (! call_f_f_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_f_f_Int_goMux1_select_d[3] && (! call_f_f_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_f_f_Int_goMux1_select_d[4] && (! call_f_f_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_f_Int_initBuf,Go) > [(call_f_f_Int_unlockFork1,Go),
                                            (call_f_f_Int_unlockFork2,Go),
                                            (call_f_f_Int_unlockFork3,Go),
                                            (call_f_f_Int_unlockFork4,Go),
                                            (call_f_f_Int_unlockFork5,Go),
                                            (call_f_f_Int_unlockFork6,Go),
                                            (call_f_f_Int_unlockFork7,Go)] */
  logic [6:0] call_f_f_Int_initBuf_emitted;
  logic [6:0] call_f_f_Int_initBuf_done;
  assign call_f_f_Int_unlockFork1_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[0]));
  assign call_f_f_Int_unlockFork2_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[1]));
  assign call_f_f_Int_unlockFork3_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[2]));
  assign call_f_f_Int_unlockFork4_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[3]));
  assign call_f_f_Int_unlockFork5_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[4]));
  assign call_f_f_Int_unlockFork6_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[5]));
  assign call_f_f_Int_unlockFork7_d = (call_f_f_Int_initBuf_d[0] && (! call_f_f_Int_initBuf_emitted[6]));
  assign call_f_f_Int_initBuf_done = (call_f_f_Int_initBuf_emitted | ({call_f_f_Int_unlockFork7_d[0],
                                                                       call_f_f_Int_unlockFork6_d[0],
                                                                       call_f_f_Int_unlockFork5_d[0],
                                                                       call_f_f_Int_unlockFork4_d[0],
                                                                       call_f_f_Int_unlockFork3_d[0],
                                                                       call_f_f_Int_unlockFork2_d[0],
                                                                       call_f_f_Int_unlockFork1_d[0]} & {call_f_f_Int_unlockFork7_r,
                                                                                                         call_f_f_Int_unlockFork6_r,
                                                                                                         call_f_f_Int_unlockFork5_r,
                                                                                                         call_f_f_Int_unlockFork4_r,
                                                                                                         call_f_f_Int_unlockFork3_r,
                                                                                                         call_f_f_Int_unlockFork2_r,
                                                                                                         call_f_f_Int_unlockFork1_r}));
  assign call_f_f_Int_initBuf_r = (& call_f_f_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_initBuf_emitted <= 7'd0;
    else
      call_f_f_Int_initBuf_emitted <= (call_f_f_Int_initBuf_r ? 7'd0 :
                                       call_f_f_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_f_Int_initBufi,Go) > (call_f_f_Int_initBuf,Go) */
  assign call_f_f_Int_initBufi_r = ((! call_f_f_Int_initBuf_d[0]) || call_f_f_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_f_f_Int_initBufi_r)
        call_f_f_Int_initBuf_d <= call_f_f_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_f_Int_unlockFork1,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11,Go)] > (call_f_f_Int_goMux1,Go) */
  assign call_f_f_Int_goMux1_d = (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d[0]);
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_r = (call_f_f_Int_goMux1_r && (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d[0]));
  assign call_f_f_Int_unlockFork1_r = (call_f_f_Int_goMux1_r && (call_f_f_Int_unlockFork1_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intgo_11_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_f_f_Int_unlockFork2,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3,Pointer_MaskQTree)] > (call_f_f_Int_goMux2,Pointer_MaskQTree) */
  assign call_f_f_Int_goMux2_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d[16:1],
                                  (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d[0])};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_r = (call_f_f_Int_goMux2_r && (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d[0]));
  assign call_f_f_Int_unlockFork2_r = (call_f_f_Int_goMux2_r && (call_f_f_Int_unlockFork2_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm1ae3_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_unlockFork3,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4,Pointer_QTree_Int)] > (call_f_f_Int_goMux3,Pointer_QTree_Int) */
  assign call_f_f_Int_goMux3_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d[16:1],
                                  (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d[0])};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_r = (call_f_f_Int_goMux3_r && (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d[0]));
  assign call_f_f_Int_unlockFork3_r = (call_f_f_Int_goMux3_r && (call_f_f_Int_unlockFork3_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm2ae4_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_unlockFork4,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5,Pointer_QTree_Int)] > (call_f_f_Int_goMux4,Pointer_QTree_Int) */
  assign call_f_f_Int_goMux4_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d[16:1],
                                  (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d[0])};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_r = (call_f_f_Int_goMux4_r && (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d[0]));
  assign call_f_f_Int_unlockFork4_r = (call_f_f_Int_goMux4_r && (call_f_f_Int_unlockFork4_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intm3ae5_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_unlockFork5,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6,MyDTInt_Bool)] > (call_f_f_Int_goMux5,MyDTInt_Bool) */
  assign call_f_f_Int_goMux5_d = (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d[0]);
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_r = (call_f_f_Int_goMux5_r && (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d[0]));
  assign call_f_f_Int_unlockFork5_r = (call_f_f_Int_goMux5_r && (call_f_f_Int_unlockFork5_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intis_zae6_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f_f_Int_unlockFork6,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7,MyDTInt_Int_Int)] > (call_f_f_Int_goMux6,MyDTInt_Int_Int) */
  assign call_f_f_Int_goMux6_d = (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d[0]);
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_r = (call_f_f_Int_goMux6_r && (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d[0]));
  assign call_f_f_Int_unlockFork6_r = (call_f_f_Int_goMux6_r && (call_f_f_Int_unlockFork6_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intop_addae7_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf_f_Int) : (call_f_f_Int_unlockFork7,Go) [(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3,Pointer_CTf_f_Int)] > (call_f_f_Int_goMux7,Pointer_CTf_f_Int) */
  assign call_f_f_Int_goMux7_d = {call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d[16:1],
                                  (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d[0])};
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_r = (call_f_f_Int_goMux7_r && (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d[0]));
  assign call_f_f_Int_unlockFork7_r = (call_f_f_Int_goMux7_r && (call_f_f_Int_unlockFork7_d[0] && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Intsc_0_3_d[0]));
  
  /* buf (Ty QTree_Int) : (es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int,QTree_Int) > (lizzieLet30_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d;
  logic es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_r;
  assign es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_r = ((! es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d[0]) || es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d <= {66'd0,
                                                              1'd0};
    else
      if (es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_r)
        es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d <= es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_d;
  QTree_Int_t es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf;
  assign es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_r = (! es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet30_1_1_argbuf_d = (es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf[0] ? es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf :
                                     es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf <= {66'd0,
                                                                1'd0};
    else
      if ((lizzieLet30_1_1_argbuf_r && es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf[0]))
        es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
      else if (((! lizzieLet30_1_1_argbuf_r) && (! es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf[0])))
        es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_buf <= es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_1,MyBool) (lizzieLet13_5QVal_Int_3QVal_Int_2,Go) > [(es_2_1MyFalse,Go),
                                                                          (es_2_1MyTrue,Go)] */
  logic [1:0] lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd;
  always_comb
    if ((es_2_1_d[0] && lizzieLet13_5QVal_Int_3QVal_Int_2_d[0]))
      unique case (es_2_1_d[1:1])
        1'd0: lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd = 2'd0;
  assign es_2_1MyFalse_d = lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd[0];
  assign es_2_1MyTrue_d = lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd[1];
  assign lizzieLet13_5QVal_Int_3QVal_Int_2_r = (| (lizzieLet13_5QVal_Int_3QVal_Int_2_onehotd & {es_2_1MyTrue_r,
                                                                                                es_2_1MyFalse_r}));
  assign es_2_1_r = lizzieLet13_5QVal_Int_3QVal_Int_2_r;
  
  /* buf (Ty Go) : (es_2_1MyFalse,Go) > (es_2_1MyFalse_1_argbuf,Go) */
  Go_t es_2_1MyFalse_bufchan_d;
  logic es_2_1MyFalse_bufchan_r;
  assign es_2_1MyFalse_r = ((! es_2_1MyFalse_bufchan_d[0]) || es_2_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_1MyFalse_r) es_2_1MyFalse_bufchan_d <= es_2_1MyFalse_d;
  Go_t es_2_1MyFalse_bufchan_buf;
  assign es_2_1MyFalse_bufchan_r = (! es_2_1MyFalse_bufchan_buf[0]);
  assign es_2_1MyFalse_1_argbuf_d = (es_2_1MyFalse_bufchan_buf[0] ? es_2_1MyFalse_bufchan_buf :
                                     es_2_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyFalse_1_argbuf_r && es_2_1MyFalse_bufchan_buf[0]))
        es_2_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyFalse_1_argbuf_r) && (! es_2_1MyFalse_bufchan_buf[0])))
        es_2_1MyFalse_bufchan_buf <= es_2_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_2_1MyTrue,Go) > [(es_2_1MyTrue_1,Go),
                                    (es_2_1MyTrue_2,Go)] */
  logic [1:0] es_2_1MyTrue_emitted;
  logic [1:0] es_2_1MyTrue_done;
  assign es_2_1MyTrue_1_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[0]));
  assign es_2_1MyTrue_2_d = (es_2_1MyTrue_d[0] && (! es_2_1MyTrue_emitted[1]));
  assign es_2_1MyTrue_done = (es_2_1MyTrue_emitted | ({es_2_1MyTrue_2_d[0],
                                                       es_2_1MyTrue_1_d[0]} & {es_2_1MyTrue_2_r,
                                                                               es_2_1MyTrue_1_r}));
  assign es_2_1MyTrue_r = (& es_2_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_emitted <= 2'd0;
    else
      es_2_1MyTrue_emitted <= (es_2_1MyTrue_r ? 2'd0 :
                               es_2_1MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_1MyTrue_1,Go)] > (es_2_1MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_1MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_1MyTrue_1_d[0]}), es_2_1MyTrue_1_d);
  assign {es_2_1MyTrue_1_r} = {1 {(es_2_1MyTrue_1QNone_Int_r && es_2_1MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_1MyTrue_1QNone_Int,QTree_Int) > (lizzieLet16_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_d;
  logic es_2_1MyTrue_1QNone_Int_bufchan_r;
  assign es_2_1MyTrue_1QNone_Int_r = ((! es_2_1MyTrue_1QNone_Int_bufchan_d[0]) || es_2_1MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_1MyTrue_1QNone_Int_r)
        es_2_1MyTrue_1QNone_Int_bufchan_d <= es_2_1MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_1MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_1MyTrue_1QNone_Int_bufchan_r = (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (es_2_1MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_1MyTrue_1QNone_Int_bufchan_buf :
                                   es_2_1MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && es_2_1MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! es_2_1MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_1MyTrue_1QNone_Int_bufchan_buf <= es_2_1MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_1MyTrue_2,Go) > (es_2_1MyTrue_2_argbuf,Go) */
  Go_t es_2_1MyTrue_2_bufchan_d;
  logic es_2_1MyTrue_2_bufchan_r;
  assign es_2_1MyTrue_2_r = ((! es_2_1MyTrue_2_bufchan_d[0]) || es_2_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_1MyTrue_2_r) es_2_1MyTrue_2_bufchan_d <= es_2_1MyTrue_2_d;
  Go_t es_2_1MyTrue_2_bufchan_buf;
  assign es_2_1MyTrue_2_bufchan_r = (! es_2_1MyTrue_2_bufchan_buf[0]);
  assign es_2_1MyTrue_2_argbuf_d = (es_2_1MyTrue_2_bufchan_buf[0] ? es_2_1MyTrue_2_bufchan_buf :
                                    es_2_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyTrue_2_argbuf_r && es_2_1MyTrue_2_bufchan_buf[0]))
        es_2_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyTrue_2_argbuf_r) && (! es_2_1MyTrue_2_bufchan_buf[0])))
        es_2_1MyTrue_2_bufchan_buf <= es_2_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_2_2,MyBool) (lizzieLet13_5QVal_Int_6QVal_Int_2,MyDTInt_Int_Int) > [(es_2_2MyFalse,MyDTInt_Int_Int),
                                                                                                    (_165,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd;
  always_comb
    if ((es_2_2_d[0] && lizzieLet13_5QVal_Int_6QVal_Int_2_d[0]))
      unique case (es_2_2_d[1:1])
        1'd0: lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd = 2'd0;
  assign es_2_2MyFalse_d = lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd[0];
  assign _165_d = lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd[1];
  assign lizzieLet13_5QVal_Int_6QVal_Int_2_r = (| (lizzieLet13_5QVal_Int_6QVal_Int_2_onehotd & {_165_r,
                                                                                                es_2_2MyFalse_r}));
  assign es_2_2_r = lizzieLet13_5QVal_Int_6QVal_Int_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_2_2MyFalse,MyDTInt_Int_Int) > (es_2_2MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_2_2MyFalse_bufchan_d;
  logic es_2_2MyFalse_bufchan_r;
  assign es_2_2MyFalse_r = ((! es_2_2MyFalse_bufchan_d[0]) || es_2_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_2MyFalse_r) es_2_2MyFalse_bufchan_d <= es_2_2MyFalse_d;
  MyDTInt_Int_Int_t es_2_2MyFalse_bufchan_buf;
  assign es_2_2MyFalse_bufchan_r = (! es_2_2MyFalse_bufchan_buf[0]);
  assign es_2_2MyFalse_1_argbuf_d = (es_2_2MyFalse_bufchan_buf[0] ? es_2_2MyFalse_bufchan_buf :
                                     es_2_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyFalse_1_argbuf_r && es_2_2MyFalse_bufchan_buf[0]))
        es_2_2MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyFalse_1_argbuf_r) && (! es_2_2MyFalse_bufchan_buf[0])))
        es_2_2MyFalse_bufchan_buf <= es_2_2MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_2_2MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_2_4MyFalse_1_argbuf,Int),
                                              (es_2_5MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_2_2MyFalse_1_argbuf_d[0],
                                                                                                       es_2_4MyFalse_1_argbuf_d[0],
                                                                                                       es_2_5MyFalse_1_argbuf_d[0]}), es_2_2MyFalse_1_argbuf_d, es_2_4MyFalse_1_argbuf_d, es_2_5MyFalse_1_argbuf_d);
  assign {es_2_2MyFalse_1_argbuf_r,
          es_2_4MyFalse_1_argbuf_r,
          es_2_5MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf'_f'_Int) : (es_2_3,MyBool) (lizzieLet13_5QVal_Int_7QVal_Int,Pointer_CTf'_f'_Int) > [(es_2_3MyFalse,Pointer_CTf'_f'_Int),
                                                                                                          (es_2_3MyTrue,Pointer_CTf'_f'_Int)] */
  logic [1:0] lizzieLet13_5QVal_Int_7QVal_Int_onehotd;
  always_comb
    if ((es_2_3_d[0] && lizzieLet13_5QVal_Int_7QVal_Int_d[0]))
      unique case (es_2_3_d[1:1])
        1'd0: lizzieLet13_5QVal_Int_7QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet13_5QVal_Int_7QVal_Int_onehotd = 2'd2;
        default: lizzieLet13_5QVal_Int_7QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet13_5QVal_Int_7QVal_Int_onehotd = 2'd0;
  assign es_2_3MyFalse_d = {lizzieLet13_5QVal_Int_7QVal_Int_d[16:1],
                            lizzieLet13_5QVal_Int_7QVal_Int_onehotd[0]};
  assign es_2_3MyTrue_d = {lizzieLet13_5QVal_Int_7QVal_Int_d[16:1],
                           lizzieLet13_5QVal_Int_7QVal_Int_onehotd[1]};
  assign lizzieLet13_5QVal_Int_7QVal_Int_r = (| (lizzieLet13_5QVal_Int_7QVal_Int_onehotd & {es_2_3MyTrue_r,
                                                                                            es_2_3MyFalse_r}));
  assign es_2_3_r = lizzieLet13_5QVal_Int_7QVal_Int_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (es_2_3MyFalse,Pointer_CTf'_f'_Int) > (es_2_3MyFalse_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  es_2_3MyFalse_bufchan_d;
  logic es_2_3MyFalse_bufchan_r;
  assign es_2_3MyFalse_r = ((! es_2_3MyFalse_bufchan_d[0]) || es_2_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_2_3MyFalse_r) es_2_3MyFalse_bufchan_d <= es_2_3MyFalse_d;
  \Pointer_CTf'_f'_Int_t  es_2_3MyFalse_bufchan_buf;
  assign es_2_3MyFalse_bufchan_r = (! es_2_3MyFalse_bufchan_buf[0]);
  assign es_2_3MyFalse_1_argbuf_d = (es_2_3MyFalse_bufchan_buf[0] ? es_2_3MyFalse_bufchan_buf :
                                     es_2_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyFalse_1_argbuf_r && es_2_3MyFalse_bufchan_buf[0]))
        es_2_3MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyFalse_1_argbuf_r) && (! es_2_3MyFalse_bufchan_buf[0])))
        es_2_3MyFalse_bufchan_buf <= es_2_3MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (es_2_3MyTrue,Pointer_CTf'_f'_Int) > (es_2_3MyTrue_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  es_2_3MyTrue_bufchan_d;
  logic es_2_3MyTrue_bufchan_r;
  assign es_2_3MyTrue_r = ((! es_2_3MyTrue_bufchan_d[0]) || es_2_3MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_d <= {16'd0, 1'd0};
    else if (es_2_3MyTrue_r) es_2_3MyTrue_bufchan_d <= es_2_3MyTrue_d;
  \Pointer_CTf'_f'_Int_t  es_2_3MyTrue_bufchan_buf;
  assign es_2_3MyTrue_bufchan_r = (! es_2_3MyTrue_bufchan_buf[0]);
  assign es_2_3MyTrue_1_argbuf_d = (es_2_3MyTrue_bufchan_buf[0] ? es_2_3MyTrue_bufchan_buf :
                                    es_2_3MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_3MyTrue_1_argbuf_r && es_2_3MyTrue_bufchan_buf[0]))
        es_2_3MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_3MyTrue_1_argbuf_r) && (! es_2_3MyTrue_bufchan_buf[0])))
        es_2_3MyTrue_bufchan_buf <= es_2_3MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_4,MyBool) (lizzieLet13_5QVal_Int_8QVal_Int_2,Int) > [(es_2_4MyFalse,Int),
                                                                            (_164,Int)] */
  logic [1:0] lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd;
  always_comb
    if ((es_2_4_d[0] && lizzieLet13_5QVal_Int_8QVal_Int_2_d[0]))
      unique case (es_2_4_d[1:1])
        1'd0: lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd = 2'd0;
  assign es_2_4MyFalse_d = {lizzieLet13_5QVal_Int_8QVal_Int_2_d[32:1],
                            lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd[0]};
  assign _164_d = {lizzieLet13_5QVal_Int_8QVal_Int_2_d[32:1],
                   lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd[1]};
  assign lizzieLet13_5QVal_Int_8QVal_Int_2_r = (| (lizzieLet13_5QVal_Int_8QVal_Int_2_onehotd & {_164_r,
                                                                                                es_2_4MyFalse_r}));
  assign es_2_4_r = lizzieLet13_5QVal_Int_8QVal_Int_2_r;
  
  /* buf (Ty Int) : (es_2_4MyFalse,Int) > (es_2_4MyFalse_1_argbuf,Int) */
  Int_t es_2_4MyFalse_bufchan_d;
  logic es_2_4MyFalse_bufchan_r;
  assign es_2_4MyFalse_r = ((! es_2_4MyFalse_bufchan_d[0]) || es_2_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_4MyFalse_r) es_2_4MyFalse_bufchan_d <= es_2_4MyFalse_d;
  Int_t es_2_4MyFalse_bufchan_buf;
  assign es_2_4MyFalse_bufchan_r = (! es_2_4MyFalse_bufchan_buf[0]);
  assign es_2_4MyFalse_1_argbuf_d = (es_2_4MyFalse_bufchan_buf[0] ? es_2_4MyFalse_bufchan_buf :
                                     es_2_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_4MyFalse_1_argbuf_r && es_2_4MyFalse_bufchan_buf[0]))
        es_2_4MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_4MyFalse_1_argbuf_r) && (! es_2_4MyFalse_bufchan_buf[0])))
        es_2_4MyFalse_bufchan_buf <= es_2_4MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_5,MyBool) (vaeM_2,Int) > [(es_2_5MyFalse,Int),
                                                 (_163,Int)] */
  logic [1:0] vaeM_2_onehotd;
  always_comb
    if ((es_2_5_d[0] && vaeM_2_d[0]))
      unique case (es_2_5_d[1:1])
        1'd0: vaeM_2_onehotd = 2'd1;
        1'd1: vaeM_2_onehotd = 2'd2;
        default: vaeM_2_onehotd = 2'd0;
      endcase
    else vaeM_2_onehotd = 2'd0;
  assign es_2_5MyFalse_d = {vaeM_2_d[32:1], vaeM_2_onehotd[0]};
  assign _163_d = {vaeM_2_d[32:1], vaeM_2_onehotd[1]};
  assign vaeM_2_r = (| (vaeM_2_onehotd & {_163_r, es_2_5MyFalse_r}));
  assign es_2_5_r = vaeM_2_r;
  
  /* buf (Ty Int) : (es_2_5MyFalse,Int) > (es_2_5MyFalse_1_argbuf,Int) */
  Int_t es_2_5MyFalse_bufchan_d;
  logic es_2_5MyFalse_bufchan_r;
  assign es_2_5MyFalse_r = ((! es_2_5MyFalse_bufchan_d[0]) || es_2_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_5MyFalse_r) es_2_5MyFalse_bufchan_d <= es_2_5MyFalse_d;
  Int_t es_2_5MyFalse_bufchan_buf;
  assign es_2_5MyFalse_bufchan_r = (! es_2_5MyFalse_bufchan_buf[0]);
  assign es_2_5MyFalse_1_argbuf_d = (es_2_5MyFalse_bufchan_buf[0] ? es_2_5MyFalse_bufchan_buf :
                                     es_2_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_5MyFalse_1_argbuf_r && es_2_5MyFalse_bufchan_buf[0]))
        es_2_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_5MyFalse_1_argbuf_r) && (! es_2_5MyFalse_bufchan_buf[0])))
        es_2_5MyFalse_bufchan_buf <= es_2_5MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_3_1QVal_Int,QTree_Int) > (lizzieLet15_1_argbuf,QTree_Int) */
  QTree_Int_t es_3_1QVal_Int_bufchan_d;
  logic es_3_1QVal_Int_bufchan_r;
  assign es_3_1QVal_Int_r = ((! es_3_1QVal_Int_bufchan_d[0]) || es_3_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_3_1QVal_Int_r) es_3_1QVal_Int_bufchan_d <= es_3_1QVal_Int_d;
  QTree_Int_t es_3_1QVal_Int_bufchan_buf;
  assign es_3_1QVal_Int_bufchan_r = (! es_3_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (es_3_1QVal_Int_bufchan_buf[0] ? es_3_1QVal_Int_bufchan_buf :
                                   es_3_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && es_3_1QVal_Int_bufchan_buf[0]))
        es_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! es_3_1QVal_Int_bufchan_buf[0])))
        es_3_1QVal_Int_bufchan_buf <= es_3_1QVal_Int_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  logic es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_r;
  assign es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_r = ((! es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d[0]) || es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= {32'd0,
                                                                  1'd0};
    else
      if (es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_r)
        es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_d;
  \Int#_t  es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf;
  assign es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_r = (! es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0] ? es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf :
                                 es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                    1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]))
        es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                      1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0])))
        es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  
  /* sink (Ty Int) : (es_6_1I#,Int) > */
  assign {\es_6_1I#_r , \es_6_1I#_dout } = {\es_6_1I#_rout ,
                                            \es_6_1I#_d };
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf_f_Int) : (es_6_1_1,MyBool) (lizzieLet24_5MQNode_6QVal_Int_3QVal_Int,Pointer_CTf_f_Int) > [(es_6_1_1MyFalse,Pointer_CTf_f_Int),
                                                                                                                (es_6_1_1MyTrue,Pointer_CTf_f_Int)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd;
  always_comb
    if ((es_6_1_1_d[0] && lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_d[0]))
      unique case (es_6_1_1_d[1:1])
        1'd0: lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd = 2'd2;
        default: lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd = 2'd0;
  assign es_6_1_1MyFalse_d = {lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_d[16:1],
                              lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd[0]};
  assign es_6_1_1MyTrue_d = {lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_d[16:1],
                             lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_r = (| (lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_onehotd & {es_6_1_1MyTrue_r,
                                                                                                            es_6_1_1MyFalse_r}));
  assign es_6_1_1_r = lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_6_1_1MyFalse,Pointer_CTf_f_Int) > (es_6_1_1MyFalse_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_6_1_1MyFalse_bufchan_d;
  logic es_6_1_1MyFalse_bufchan_r;
  assign es_6_1_1MyFalse_r = ((! es_6_1_1MyFalse_bufchan_d[0]) || es_6_1_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_1MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_6_1_1MyFalse_r)
        es_6_1_1MyFalse_bufchan_d <= es_6_1_1MyFalse_d;
  Pointer_CTf_f_Int_t es_6_1_1MyFalse_bufchan_buf;
  assign es_6_1_1MyFalse_bufchan_r = (! es_6_1_1MyFalse_bufchan_buf[0]);
  assign es_6_1_1MyFalse_1_argbuf_d = (es_6_1_1MyFalse_bufchan_buf[0] ? es_6_1_1MyFalse_bufchan_buf :
                                       es_6_1_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_1MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_6_1_1MyFalse_1_argbuf_r && es_6_1_1MyFalse_bufchan_buf[0]))
        es_6_1_1MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_6_1_1MyFalse_1_argbuf_r) && (! es_6_1_1MyFalse_bufchan_buf[0])))
        es_6_1_1MyFalse_bufchan_buf <= es_6_1_1MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (es_6_1_1MyTrue,Pointer_CTf_f_Int) > (es_6_1_1MyTrue_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t es_6_1_1MyTrue_bufchan_d;
  logic es_6_1_1MyTrue_bufchan_r;
  assign es_6_1_1MyTrue_r = ((! es_6_1_1MyTrue_bufchan_d[0]) || es_6_1_1MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_1MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_6_1_1MyTrue_r) es_6_1_1MyTrue_bufchan_d <= es_6_1_1MyTrue_d;
  Pointer_CTf_f_Int_t es_6_1_1MyTrue_bufchan_buf;
  assign es_6_1_1MyTrue_bufchan_r = (! es_6_1_1MyTrue_bufchan_buf[0]);
  assign es_6_1_1MyTrue_1_argbuf_d = (es_6_1_1MyTrue_bufchan_buf[0] ? es_6_1_1MyTrue_bufchan_buf :
                                      es_6_1_1MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_1MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_6_1_1MyTrue_1_argbuf_r && es_6_1_1MyTrue_bufchan_buf[0]))
        es_6_1_1MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_6_1_1MyTrue_1_argbuf_r) && (! es_6_1_1MyTrue_bufchan_buf[0])))
        es_6_1_1MyTrue_bufchan_buf <= es_6_1_1MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_6_1_2,MyBool) (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2,Go) > [(es_6_1_2MyFalse,Go),
                                                                                    (es_6_1_2MyTrue,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd;
  always_comb
    if ((es_6_1_2_d[0] && lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_d[0]))
      unique case (es_6_1_2_d[1:1])
        1'd0: lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd = 2'd0;
  assign es_6_1_2MyFalse_d = lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd[0];
  assign es_6_1_2MyTrue_d = lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd[1];
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_r = (| (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_onehotd & {es_6_1_2MyTrue_r,
                                                                                                                es_6_1_2MyFalse_r}));
  assign es_6_1_2_r = lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_r;
  
  /* fork (Ty Go) : (es_6_1_2MyFalse,Go) > [(es_6_1_2MyFalse_1,Go),
                                       (es_6_1_2MyFalse_2,Go)] */
  logic [1:0] es_6_1_2MyFalse_emitted;
  logic [1:0] es_6_1_2MyFalse_done;
  assign es_6_1_2MyFalse_1_d = (es_6_1_2MyFalse_d[0] && (! es_6_1_2MyFalse_emitted[0]));
  assign es_6_1_2MyFalse_2_d = (es_6_1_2MyFalse_d[0] && (! es_6_1_2MyFalse_emitted[1]));
  assign es_6_1_2MyFalse_done = (es_6_1_2MyFalse_emitted | ({es_6_1_2MyFalse_2_d[0],
                                                             es_6_1_2MyFalse_1_d[0]} & {es_6_1_2MyFalse_2_r,
                                                                                        es_6_1_2MyFalse_1_r}));
  assign es_6_1_2MyFalse_r = (& es_6_1_2MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyFalse_emitted <= 2'd0;
    else
      es_6_1_2MyFalse_emitted <= (es_6_1_2MyFalse_r ? 2'd0 :
                                  es_6_1_2MyFalse_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(es_6_1_2MyFalse_1,Go)] > (es_6_1_2MyFalse_1QError_Int,QTree_Int) */
  assign es_6_1_2MyFalse_1QError_Int_d = QError_Int_dc((& {es_6_1_2MyFalse_1_d[0]}), es_6_1_2MyFalse_1_d);
  assign {es_6_1_2MyFalse_1_r} = {1 {(es_6_1_2MyFalse_1QError_Int_r && es_6_1_2MyFalse_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_6_1_2MyFalse_1QError_Int,QTree_Int) > (lizzieLet34_1_argbuf,QTree_Int) */
  QTree_Int_t es_6_1_2MyFalse_1QError_Int_bufchan_d;
  logic es_6_1_2MyFalse_1QError_Int_bufchan_r;
  assign es_6_1_2MyFalse_1QError_Int_r = ((! es_6_1_2MyFalse_1QError_Int_bufchan_d[0]) || es_6_1_2MyFalse_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_6_1_2MyFalse_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_6_1_2MyFalse_1QError_Int_r)
        es_6_1_2MyFalse_1QError_Int_bufchan_d <= es_6_1_2MyFalse_1QError_Int_d;
  QTree_Int_t es_6_1_2MyFalse_1QError_Int_bufchan_buf;
  assign es_6_1_2MyFalse_1QError_Int_bufchan_r = (! es_6_1_2MyFalse_1QError_Int_bufchan_buf[0]);
  assign lizzieLet34_1_argbuf_d = (es_6_1_2MyFalse_1QError_Int_bufchan_buf[0] ? es_6_1_2MyFalse_1QError_Int_bufchan_buf :
                                   es_6_1_2MyFalse_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_6_1_2MyFalse_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && es_6_1_2MyFalse_1QError_Int_bufchan_buf[0]))
        es_6_1_2MyFalse_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! es_6_1_2MyFalse_1QError_Int_bufchan_buf[0])))
        es_6_1_2MyFalse_1QError_Int_bufchan_buf <= es_6_1_2MyFalse_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_6_1_2MyFalse_2,Go) > (es_6_1_2MyFalse_2_argbuf,Go) */
  Go_t es_6_1_2MyFalse_2_bufchan_d;
  logic es_6_1_2MyFalse_2_bufchan_r;
  assign es_6_1_2MyFalse_2_r = ((! es_6_1_2MyFalse_2_bufchan_d[0]) || es_6_1_2MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_6_1_2MyFalse_2_r)
        es_6_1_2MyFalse_2_bufchan_d <= es_6_1_2MyFalse_2_d;
  Go_t es_6_1_2MyFalse_2_bufchan_buf;
  assign es_6_1_2MyFalse_2_bufchan_r = (! es_6_1_2MyFalse_2_bufchan_buf[0]);
  assign es_6_1_2MyFalse_2_argbuf_d = (es_6_1_2MyFalse_2_bufchan_buf[0] ? es_6_1_2MyFalse_2_bufchan_buf :
                                       es_6_1_2MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_6_1_2MyFalse_2_argbuf_r && es_6_1_2MyFalse_2_bufchan_buf[0]))
        es_6_1_2MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_6_1_2MyFalse_2_argbuf_r) && (! es_6_1_2MyFalse_2_bufchan_buf[0])))
        es_6_1_2MyFalse_2_bufchan_buf <= es_6_1_2MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_6_1_2MyTrue,Go) > [(es_6_1_2MyTrue_1,Go),
                                      (es_6_1_2MyTrue_2,Go)] */
  logic [1:0] es_6_1_2MyTrue_emitted;
  logic [1:0] es_6_1_2MyTrue_done;
  assign es_6_1_2MyTrue_1_d = (es_6_1_2MyTrue_d[0] && (! es_6_1_2MyTrue_emitted[0]));
  assign es_6_1_2MyTrue_2_d = (es_6_1_2MyTrue_d[0] && (! es_6_1_2MyTrue_emitted[1]));
  assign es_6_1_2MyTrue_done = (es_6_1_2MyTrue_emitted | ({es_6_1_2MyTrue_2_d[0],
                                                           es_6_1_2MyTrue_1_d[0]} & {es_6_1_2MyTrue_2_r,
                                                                                     es_6_1_2MyTrue_1_r}));
  assign es_6_1_2MyTrue_r = (& es_6_1_2MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyTrue_emitted <= 2'd0;
    else
      es_6_1_2MyTrue_emitted <= (es_6_1_2MyTrue_r ? 2'd0 :
                                 es_6_1_2MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_6_1_2MyTrue_1,Go)] > (es_6_1_2MyTrue_1QNone_Int,QTree_Int) */
  assign es_6_1_2MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_6_1_2MyTrue_1_d[0]}), es_6_1_2MyTrue_1_d);
  assign {es_6_1_2MyTrue_1_r} = {1 {(es_6_1_2MyTrue_1QNone_Int_r && es_6_1_2MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_6_1_2MyTrue_1QNone_Int,QTree_Int) > (lizzieLet35_1_argbuf,QTree_Int) */
  QTree_Int_t es_6_1_2MyTrue_1QNone_Int_bufchan_d;
  logic es_6_1_2MyTrue_1QNone_Int_bufchan_r;
  assign es_6_1_2MyTrue_1QNone_Int_r = ((! es_6_1_2MyTrue_1QNone_Int_bufchan_d[0]) || es_6_1_2MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_6_1_2MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_6_1_2MyTrue_1QNone_Int_r)
        es_6_1_2MyTrue_1QNone_Int_bufchan_d <= es_6_1_2MyTrue_1QNone_Int_d;
  QTree_Int_t es_6_1_2MyTrue_1QNone_Int_bufchan_buf;
  assign es_6_1_2MyTrue_1QNone_Int_bufchan_r = (! es_6_1_2MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet35_1_argbuf_d = (es_6_1_2MyTrue_1QNone_Int_bufchan_buf[0] ? es_6_1_2MyTrue_1QNone_Int_bufchan_buf :
                                   es_6_1_2MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_6_1_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && es_6_1_2MyTrue_1QNone_Int_bufchan_buf[0]))
        es_6_1_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! es_6_1_2MyTrue_1QNone_Int_bufchan_buf[0])))
        es_6_1_2MyTrue_1QNone_Int_bufchan_buf <= es_6_1_2MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_6_1_2MyTrue_2,Go) > (es_6_1_2MyTrue_2_argbuf,Go) */
  Go_t es_6_1_2MyTrue_2_bufchan_d;
  logic es_6_1_2MyTrue_2_bufchan_r;
  assign es_6_1_2MyTrue_2_r = ((! es_6_1_2MyTrue_2_bufchan_d[0]) || es_6_1_2MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_6_1_2MyTrue_2_r)
        es_6_1_2MyTrue_2_bufchan_d <= es_6_1_2MyTrue_2_d;
  Go_t es_6_1_2MyTrue_2_bufchan_buf;
  assign es_6_1_2MyTrue_2_bufchan_r = (! es_6_1_2MyTrue_2_bufchan_buf[0]);
  assign es_6_1_2MyTrue_2_argbuf_d = (es_6_1_2MyTrue_2_bufchan_buf[0] ? es_6_1_2MyTrue_2_bufchan_buf :
                                      es_6_1_2MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_6_1_2MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_6_1_2MyTrue_2_argbuf_r && es_6_1_2MyTrue_2_bufchan_buf[0]))
        es_6_1_2MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_6_1_2MyTrue_2_argbuf_r) && (! es_6_1_2MyTrue_2_bufchan_buf[0])))
        es_6_1_2MyTrue_2_bufchan_buf <= es_6_1_2MyTrue_2_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_2_1ww2Xku_1_1_Add32,Int#) (lizzieLet46_4Lcall_$wnnz_Int0,Int#) > (es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32,Int#) */
  assign es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_d = {(es_6_2_1ww2Xku_1_1_Add32_d[32:1] + lizzieLet46_4Lcall_$wnnz_Int0_d[32:1]),
                                                            (es_6_2_1ww2Xku_1_1_Add32_d[0] && lizzieLet46_4Lcall_$wnnz_Int0_d[0])};
  assign {es_6_2_1ww2Xku_1_1_Add32_r,
          lizzieLet46_4Lcall_$wnnz_Int0_r} = {2 {(es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_r && es_4_1_1lizzieLet46_4Lcall_$wnnz_Int0_1_Add32_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_7_1es_8_1es_9_1es_10_1QNode_Int,QTree_Int) > (lizzieLet38_1_argbuf,QTree_Int) */
  QTree_Int_t es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d;
  logic es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_r;
  assign es_7_1es_8_1es_9_1es_10_1QNode_Int_r = ((! es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d[0]) || es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_7_1es_8_1es_9_1es_10_1QNode_Int_r)
        es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d <= es_7_1es_8_1es_9_1es_10_1QNode_Int_d;
  QTree_Int_t es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf;
  assign es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_r = (! es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet38_1_argbuf_d = (es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf[0] ? es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf :
                                   es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf[0]))
        es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf[0])))
        es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_buf <= es_7_1es_8_1es_9_1es_10_1QNode_Int_bufchan_d;
  
  /* mergectrl (Ty C8,
           Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7,TupGo___Pointer_MaskQTree___Pointer_QTree_Int),
                                                                (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8,TupGo___Pointer_MaskQTree___Pointer_QTree_Int)] > (f'''''''''_f'''''''''_Int_choice,C8) (f'''''''''_f'''''''''_Int_data,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  logic [7:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d  = ((| \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_q ) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_q  :
                                                                                                (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_d [0] ? 8'd1 :
                                                                                                 (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_d [0] ? 8'd2 :
                                                                                                  (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_d [0] ? 8'd4 :
                                                                                                   (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_d [0] ? 8'd8 :
                                                                                                    (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_d [0] ? 8'd16 :
                                                                                                     (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_d [0] ? 8'd32 :
                                                                                                      (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_d [0] ? 8'd64 :
                                                                                                       (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_d [0] ? 8'd128 :
                                                                                                        8'd0)))))))));
  logic [7:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_q  <= 8'd0;
    else
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_q  <= (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_done  ? 8'd0 :
                                                                                              \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d );
  logic [1:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q  <= 2'd0;
    else
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q  <= (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_done  ? 2'd0 :
                                                                                            \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_d );
  logic [1:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_d ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_d  = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q  | ({\f'''''''''_f'''''''''_Int_choice_d [0],
                                                                                                                                                                                    \f'''''''''_f'''''''''_Int_data_d [0]} & {\f'''''''''_f'''''''''_Int_choice_r ,
                                                                                                                                                                                                                              \f'''''''''_f'''''''''_Int_data_r }));
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_done ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_done  = (& \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_d );
  assign {\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_r ,
          \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_r } = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_done  ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d  :
                                                                                           8'd0);
  assign \f'''''''''_f'''''''''_Int_data_d  = ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [0] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_d  :
                                               ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [1] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_d  :
                                                ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [2] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_d  :
                                                 ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [3] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_d  :
                                                  ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [4] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_d  :
                                                   ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [5] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_d  :
                                                    ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [6] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_d  :
                                                     ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [7] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [0])) ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_d  :
                                                      {32'd0, 1'd0}))))))));
  assign \f'''''''''_f'''''''''_Int_choice_d  = ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [0] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C1_8_dc(1'd1) :
                                                 ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [1] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C2_8_dc(1'd1) :
                                                  ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [2] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C3_8_dc(1'd1) :
                                                   ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [3] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C4_8_dc(1'd1) :
                                                    ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [4] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C5_8_dc(1'd1) :
                                                     ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [5] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C6_8_dc(1'd1) :
                                                      ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [6] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C7_8_dc(1'd1) :
                                                       ((\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_select_d [7] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_emit_q [1])) ? C8_8_dc(1'd1) :
                                                        {3'd0, 1'd0}))))))));
  
  /* fork (Ty Go) : (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12,Go) > [(go_12_1,Go),
                                                                                                   (go_12_2,Go)] */
  logic [1:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted ;
  logic [1:0] \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_done ;
  assign go_12_1_d = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_d [0] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted [0]));
  assign go_12_2_d = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_d [0] && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted [1]));
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_done  = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted  | ({go_12_2_d[0],
                                                                                                                                                                                         go_12_1_d[0]} & {go_12_2_r,
                                                                                                                                                                                                          go_12_1_r}));
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_r  = (& \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted  <= 2'd0;
    else
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_emitted  <= (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_r  ? 2'd0 :
                                                                                                \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_done );
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1,Pointer_QTree_Int) > (q4'aex_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_r  = ((! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d [0]) || \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d  <= {16'd0,
                                                                                                     1'd0};
    else
      if (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_r )
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d  <= \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_r  = (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf [0]);
  assign \q4'aex_1_1_argbuf_d  = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf  :
                                  \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf  <= {16'd0,
                                                                                                       1'd0};
    else
      if ((\q4'aex_1_1_argbuf_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
      else if (((! \q4'aex_1_1_argbuf_r ) && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_buf  <= \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_bufchan_d ;
  
  /* buf (Ty Pointer_MaskQTree) : (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1,Pointer_MaskQTree) > (q4aew_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_r  = ((! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d [0]) || \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d  <= {16'd0,
                                                                                                    1'd0};
    else
      if (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_r )
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d  <= \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_d ;
  Pointer_MaskQTree_t \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_r  = (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf [0]);
  assign q4aew_1_1_argbuf_d = (\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf  :
                               \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf  <= {16'd0,
                                                                                                      1'd0};
    else
      if ((q4aew_1_1_argbuf_r && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf  <= {16'd0,
                                                                                                        1'd0};
      else if (((! q4aew_1_1_argbuf_r) && (! \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_buf  <= \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_1,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_1_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_1_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_1_r  = ((! \f'''''''''_f'''''''''_Int_1_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_1_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_1_r )
        \f'''''''''_f'''''''''_Int_1_bufchan_d  <= \f'''''''''_f'''''''''_Int_1_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_1_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_1_bufchan_r  = (! \f'''''''''_f'''''''''_Int_1_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_resbuf_d  = (\f'''''''''_f'''''''''_Int_1_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_1_bufchan_buf  :
                                                 \f'''''''''_f'''''''''_Int_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_resbuf_r  && \f'''''''''_f'''''''''_Int_1_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_resbuf_r ) && (! \f'''''''''_f'''''''''_Int_1_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_1_bufchan_buf  <= \f'''''''''_f'''''''''_Int_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_2,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_2_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_2_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_2_r  = ((! \f'''''''''_f'''''''''_Int_2_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_2_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_2_r )
        \f'''''''''_f'''''''''_Int_2_bufchan_d  <= \f'''''''''_f'''''''''_Int_2_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_2_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_2_bufchan_r  = (! \f'''''''''_f'''''''''_Int_2_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_2_argbuf_d  = (\f'''''''''_f'''''''''_Int_2_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_2_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_2_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_2_argbuf_r  && \f'''''''''_f'''''''''_Int_2_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_2_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_2_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_2_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_2_bufchan_buf  <= \f'''''''''_f'''''''''_Int_2_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_3,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_3_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_3_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_3_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_3_r  = ((! \f'''''''''_f'''''''''_Int_3_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_3_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_3_r )
        \f'''''''''_f'''''''''_Int_3_bufchan_d  <= \f'''''''''_f'''''''''_Int_3_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_3_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_3_bufchan_r  = (! \f'''''''''_f'''''''''_Int_3_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_3_argbuf_d  = (\f'''''''''_f'''''''''_Int_3_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_3_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_3_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_3_argbuf_r  && \f'''''''''_f'''''''''_Int_3_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_3_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_3_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_3_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_3_bufchan_buf  <= \f'''''''''_f'''''''''_Int_3_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_4,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_4_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_4_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_4_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_4_r  = ((! \f'''''''''_f'''''''''_Int_4_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_4_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_4_r )
        \f'''''''''_f'''''''''_Int_4_bufchan_d  <= \f'''''''''_f'''''''''_Int_4_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_4_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_4_bufchan_r  = (! \f'''''''''_f'''''''''_Int_4_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_4_argbuf_d  = (\f'''''''''_f'''''''''_Int_4_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_4_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_4_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_4_argbuf_r  && \f'''''''''_f'''''''''_Int_4_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_4_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_4_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_4_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_4_bufchan_buf  <= \f'''''''''_f'''''''''_Int_4_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f'''''''''_f'''''''''_Int_4_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_3_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_2_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_resbuf,Pointer_QTree_Int)] > (es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int,QTree_Int) */
  assign es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_d = QNode_Int_dc((& {\f'''''''''_f'''''''''_Int_4_argbuf_d [0],
                                                                        \f'''''''''_f'''''''''_Int_3_argbuf_d [0],
                                                                        \f'''''''''_f'''''''''_Int_2_argbuf_d [0],
                                                                        \f'''''''''_f'''''''''_Int_resbuf_d [0]}), \f'''''''''_f'''''''''_Int_4_argbuf_d , \f'''''''''_f'''''''''_Int_3_argbuf_d , \f'''''''''_f'''''''''_Int_2_argbuf_d , \f'''''''''_f'''''''''_Int_resbuf_d );
  assign {\f'''''''''_f'''''''''_Int_4_argbuf_r ,
          \f'''''''''_f'''''''''_Int_3_argbuf_r ,
          \f'''''''''_f'''''''''_Int_2_argbuf_r ,
          \f'''''''''_f'''''''''_Int_resbuf_r } = {4 {(es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_r && es_0_2_1es_1_1_1es_2_1_1es_3_1_1QNode_Int_d[0])}};
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_5,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_5_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_5_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_5_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_5_r  = ((! \f'''''''''_f'''''''''_Int_5_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_5_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_5_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_5_r )
        \f'''''''''_f'''''''''_Int_5_bufchan_d  <= \f'''''''''_f'''''''''_Int_5_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_5_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_5_bufchan_r  = (! \f'''''''''_f'''''''''_Int_5_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_5_argbuf_d  = (\f'''''''''_f'''''''''_Int_5_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_5_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_5_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_5_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_5_argbuf_r  && \f'''''''''_f'''''''''_Int_5_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_5_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_5_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_5_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_5_bufchan_buf  <= \f'''''''''_f'''''''''_Int_5_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_6,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_6_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_6_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_6_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_6_r  = ((! \f'''''''''_f'''''''''_Int_6_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_6_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_6_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_6_r )
        \f'''''''''_f'''''''''_Int_6_bufchan_d  <= \f'''''''''_f'''''''''_Int_6_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_6_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_6_bufchan_r  = (! \f'''''''''_f'''''''''_Int_6_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_6_argbuf_d  = (\f'''''''''_f'''''''''_Int_6_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_6_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_6_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_6_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_6_argbuf_r  && \f'''''''''_f'''''''''_Int_6_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_6_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_6_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_6_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_6_bufchan_buf  <= \f'''''''''_f'''''''''_Int_6_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_7,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_7_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_7_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_7_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_7_r  = ((! \f'''''''''_f'''''''''_Int_7_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_7_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_7_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_7_r )
        \f'''''''''_f'''''''''_Int_7_bufchan_d  <= \f'''''''''_f'''''''''_Int_7_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_7_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_7_bufchan_r  = (! \f'''''''''_f'''''''''_Int_7_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_7_argbuf_d  = (\f'''''''''_f'''''''''_Int_7_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_7_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_7_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_7_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_7_argbuf_r  && \f'''''''''_f'''''''''_Int_7_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_7_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_7_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_7_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_7_bufchan_buf  <= \f'''''''''_f'''''''''_Int_7_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_8,Pointer_QTree_Int) > (f'''''''''_f'''''''''_Int_8_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_8_bufchan_d ;
  logic \f'''''''''_f'''''''''_Int_8_bufchan_r ;
  assign \f'''''''''_f'''''''''_Int_8_r  = ((! \f'''''''''_f'''''''''_Int_8_bufchan_d [0]) || \f'''''''''_f'''''''''_Int_8_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_8_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'''''''''_f'''''''''_Int_8_r )
        \f'''''''''_f'''''''''_Int_8_bufchan_d  <= \f'''''''''_f'''''''''_Int_8_d ;
  Pointer_QTree_Int_t \f'''''''''_f'''''''''_Int_8_bufchan_buf ;
  assign \f'''''''''_f'''''''''_Int_8_bufchan_r  = (! \f'''''''''_f'''''''''_Int_8_bufchan_buf [0]);
  assign \f'''''''''_f'''''''''_Int_8_argbuf_d  = (\f'''''''''_f'''''''''_Int_8_bufchan_buf [0] ? \f'''''''''_f'''''''''_Int_8_bufchan_buf  :
                                                   \f'''''''''_f'''''''''_Int_8_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_8_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\f'''''''''_f'''''''''_Int_8_argbuf_r  && \f'''''''''_f'''''''''_Int_8_bufchan_buf [0]))
        \f'''''''''_f'''''''''_Int_8_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \f'''''''''_f'''''''''_Int_8_argbuf_r ) && (! \f'''''''''_f'''''''''_Int_8_bufchan_buf [0])))
        \f'''''''''_f'''''''''_Int_8_bufchan_buf  <= \f'''''''''_f'''''''''_Int_8_bufchan_d ;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(f'''''''''_f'''''''''_Int_8_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_7_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_6_argbuf,Pointer_QTree_Int),
                         (f'''''''''_f'''''''''_Int_5_argbuf,Pointer_QTree_Int)] > (es_7_1es_8_1es_9_1es_10_1QNode_Int,QTree_Int) */
  assign es_7_1es_8_1es_9_1es_10_1QNode_Int_d = QNode_Int_dc((& {\f'''''''''_f'''''''''_Int_8_argbuf_d [0],
                                                                 \f'''''''''_f'''''''''_Int_7_argbuf_d [0],
                                                                 \f'''''''''_f'''''''''_Int_6_argbuf_d [0],
                                                                 \f'''''''''_f'''''''''_Int_5_argbuf_d [0]}), \f'''''''''_f'''''''''_Int_8_argbuf_d , \f'''''''''_f'''''''''_Int_7_argbuf_d , \f'''''''''_f'''''''''_Int_6_argbuf_d , \f'''''''''_f'''''''''_Int_5_argbuf_d );
  assign {\f'''''''''_f'''''''''_Int_8_argbuf_r ,
          \f'''''''''_f'''''''''_Int_7_argbuf_r ,
          \f'''''''''_f'''''''''_Int_6_argbuf_r ,
          \f'''''''''_f'''''''''_Int_5_argbuf_r } = {4 {(es_7_1es_8_1es_9_1es_10_1QNode_Int_r && es_7_1es_8_1es_9_1es_10_1QNode_Int_d[0])}};
  
  /* demux (Ty C8,
       Ty Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_choice,C8) (lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > [(f'''''''''_f'''''''''_Int_1,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_2,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_3,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_4,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_5,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_6,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_7,Pointer_QTree_Int),
                                                                                                                                                             (f'''''''''_f'''''''''_Int_8,Pointer_QTree_Int)] */
  logic [7:0] \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd ;
  always_comb
    if ((\f'''''''''_f'''''''''_Int_choice_d [0] && \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [0]))
      unique case (\f'''''''''_f'''''''''_Int_choice_d [3:1])
        3'd0:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd1;
        3'd1:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd2;
        3'd2:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd4;
        3'd3:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd8;
        3'd4:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd16;
        3'd5:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd32;
        3'd6:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd64;
        3'd7:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd128;
        default:
          \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
      endcase
    else
      \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  = 8'd0;
  assign \f'''''''''_f'''''''''_Int_1_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [0]};
  assign \f'''''''''_f'''''''''_Int_2_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [1]};
  assign \f'''''''''_f'''''''''_Int_3_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [2]};
  assign \f'''''''''_f'''''''''_Int_4_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [3]};
  assign \f'''''''''_f'''''''''_Int_5_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [4]};
  assign \f'''''''''_f'''''''''_Int_6_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [5]};
  assign \f'''''''''_f'''''''''_Int_7_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [6]};
  assign \f'''''''''_f'''''''''_Int_8_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [16:1],
                                            \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd [7]};
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_r  = (| (\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_onehotd  & {\f'''''''''_f'''''''''_Int_8_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_7_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_6_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_5_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_4_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_3_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_2_r ,
                                                                                                                                                                  \f'''''''''_f'''''''''_Int_1_r }));
  assign \f'''''''''_f'''''''''_Int_choice_r  = \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_r ;
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : (f'''''''''_f'''''''''_Int_data,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) > [(f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12,Go),
                                                                                                                                                  (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1,Pointer_MaskQTree),
                                                                                                                                                  (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1,Pointer_QTree_Int)] */
  logic [2:0] \f'''''''''_f'''''''''_Int_data_emitted ;
  logic [2:0] \f'''''''''_f'''''''''_Int_data_done ;
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_d  = (\f'''''''''_f'''''''''_Int_data_d [0] && (! \f'''''''''_f'''''''''_Int_data_emitted [0]));
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_d  = {\f'''''''''_f'''''''''_Int_data_d [16:1],
                                                                                              (\f'''''''''_f'''''''''_Int_data_d [0] && (! \f'''''''''_f'''''''''_Int_data_emitted [1]))};
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_d  = {\f'''''''''_f'''''''''_Int_data_d [32:17],
                                                                                               (\f'''''''''_f'''''''''_Int_data_d [0] && (! \f'''''''''_f'''''''''_Int_data_emitted [2]))};
  assign \f'''''''''_f'''''''''_Int_data_done  = (\f'''''''''_f'''''''''_Int_data_emitted  | ({\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_d [0],
                                                                                               \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_d [0],
                                                                                               \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_d [0]} & {\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4'aex_1_r ,
                                                                                                                                                                                      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intq4aew_1_r ,
                                                                                                                                                                                      \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Intgo_12_r }));
  assign \f'''''''''_f'''''''''_Int_data_r  = (& \f'''''''''_f'''''''''_Int_data_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'''''''''_f'''''''''_Int_data_emitted  <= 3'd0;
    else
      \f'''''''''_f'''''''''_Int_data_emitted  <= (\f'''''''''_f'''''''''_Int_data_r  ? 3'd0 :
                                                   \f'''''''''_f'''''''''_Int_data_done );
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) > [(f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13,Go),
                                                                                                                                                                                                                                                                               (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                               (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                               (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                               (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1,MyDTInt_Int_Int)] */
  logic [4:0] \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted ;
  logic [4:0] \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_d  = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted [0]));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_d  = {\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [16:1],
                                                                                                               (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted [1]))};
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_d  = {\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [32:17],
                                                                                                               (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted [2]))};
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_d  = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted [3]));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_d  = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted [4]));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done  = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted  | ({\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_d [0],
                                                                                                                                                                                                                     \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_d [0],
                                                                                                                                                                                                                     \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_d [0],
                                                                                                                                                                                                                     \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_d [0],
                                                                                                                                                                                                                     \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_d [0]} & {\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_r ,
                                                                                                                                                                                                                                                                                                                             \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_r ,
                                                                                                                                                                                                                                                                                                                             \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_r ,
                                                                                                                                                                                                                                                                                                                             \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_r ,
                                                                                                                                                                                                                                                                                                                             \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_r }));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r  = (& \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted  <= 5'd0;
    else
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted  <= (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r  ? 5'd0 :
                                                                                                              \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done );
  
  /* fork (Ty Go) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13,Go) > [(go_13_1,Go),
                                                                                                                    (go_13_2,Go)] */
  logic [1:0] \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted ;
  logic [1:0] \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_done ;
  assign go_13_1_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted [0]));
  assign go_13_2_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_d [0] && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted [1]));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_done  = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted  | ({go_13_2_d[0],
                                                                                                                                                                                                                           go_13_1_d[0]} & {go_13_2_r,
                                                                                                                                                                                                                                            go_13_1_r}));
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_r  = (& \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted  <= 2'd0;
    else
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_emitted  <= (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_r  ? 2'd0 :
                                                                                                                 \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_13_done );
  
  /* buf (Ty MyDTInt_Bool) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1,MyDTInt_Bool) > (is_zaeJ_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_r ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_r  = ((! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d [0]) || \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_r )
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_d ;
  MyDTInt_Bool_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_r  = (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf [0]);
  assign is_zaeJ_1_1_argbuf_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf [0] ? \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf  :
                                 \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf  <= 1'd0;
    else
      if ((is_zaeJ_1_1_argbuf_r && \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf [0]))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf  <= 1'd0;
      else if (((! is_zaeJ_1_1_argbuf_r) && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf [0])))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_buf  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zaeJ_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1,Pointer_QTree_Int) > (m2aeH_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_r ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_r  = ((! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d [0]) || \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d  <= {16'd0,
                                                                                                                     1'd0};
    else
      if (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_r )
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_d ;
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_r  = (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf [0]);
  assign m2aeH_1_1_argbuf_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf [0] ? \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf  :
                               \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf  <= {16'd0,
                                                                                                                       1'd0};
    else
      if ((m2aeH_1_1_argbuf_r && \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf [0]))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf  <= {16'd0,
                                                                                                                         1'd0};
      else if (((! m2aeH_1_1_argbuf_r) && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf [0])))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_buf  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2aeH_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1,Pointer_QTree_Int) > (m3aeI_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_r ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_r  = ((! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d [0]) || \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d  <= {16'd0,
                                                                                                                     1'd0};
    else
      if (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_r )
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_d ;
  Pointer_QTree_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_r  = (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf [0]);
  assign m3aeI_1_1_argbuf_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf [0] ? \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf  :
                               \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf  <= {16'd0,
                                                                                                                       1'd0};
    else
      if ((m3aeI_1_1_argbuf_r && \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf [0]))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf  <= {16'd0,
                                                                                                                         1'd0};
      else if (((! m3aeI_1_1_argbuf_r) && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf [0])))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_buf  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3aeI_1_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int_Int) : (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1,MyDTInt_Int_Int) > (op_addaeK_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d ;
  logic \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_r ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_r  = ((! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d [0]) || \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_r )
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_d ;
  MyDTInt_Int_Int_t \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf ;
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_r  = (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf [0]);
  assign op_addaeK_1_1_argbuf_d = (\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf [0] ? \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf  :
                                   \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf  <= 1'd0;
    else
      if ((op_addaeK_1_1_argbuf_r && \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf [0]))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf  <= 1'd0;
      else if (((! op_addaeK_1_1_argbuf_r) && (! \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf [0])))
        \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_buf  <= \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addaeK_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'_f'_Int_resbuf,Pointer_QTree_Int) > (lizzieLet14_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'_f'_Int_resbuf_bufchan_d ;
  logic \f'_f'_Int_resbuf_bufchan_r ;
  assign \f'_f'_Int_resbuf_r  = ((! \f'_f'_Int_resbuf_bufchan_d [0]) || \f'_f'_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \f'_f'_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'_f'_Int_resbuf_r )
        \f'_f'_Int_resbuf_bufchan_d  <= \f'_f'_Int_resbuf_d ;
  Pointer_QTree_Int_t \f'_f'_Int_resbuf_bufchan_buf ;
  assign \f'_f'_Int_resbuf_bufchan_r  = (! \f'_f'_Int_resbuf_bufchan_buf [0]);
  assign lizzieLet14_1_1_argbuf_d = (\f'_f'_Int_resbuf_bufchan_buf [0] ? \f'_f'_Int_resbuf_bufchan_buf  :
                                     \f'_f'_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && \f'_f'_Int_resbuf_bufchan_buf [0]))
        \f'_f'_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! \f'_f'_Int_resbuf_bufchan_buf [0])))
        \f'_f'_Int_resbuf_bufchan_buf  <= \f'_f'_Int_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
          Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) > [(f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14,Go),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                         (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1,MyDTInt_Int_Int)] */
  logic [5:0] f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted;
  logic [5:0] f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[0]));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_d = {f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[16:1],
                                                                                                                               (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[1]))};
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_d = {f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[32:17],
                                                                                                                               (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[2]))};
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_d = {f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[48:33],
                                                                                                                               (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[3]))};
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[4]));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted[5]));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted | ({f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_d[0],
                                                                                                                                                                                                                                                     f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0]} & {f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_r,
                                                                                                                                                                                                                                                                                                                                                                             f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r}));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r = (& f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= 6'd0;
    else
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_emitted <= (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r ? 6'd0 :
                                                                                                                              f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_done);
  
  /* fork (Ty Go) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14,Go) > [(go_14_1,Go),
                                                                                                                                      (go_14_2,Go)] */
  logic [1:0] f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted;
  logic [1:0] f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done;
  assign go_14_1_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted[0]));
  assign go_14_2_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_d[0] && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted[1]));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted | ({go_14_2_d[0],
                                                                                                                                                                                                                                                           go_14_1_d[0]} & {go_14_2_r,
                                                                                                                                                                                                                                                                            go_14_1_r}));
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r = (& f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted <= 2'd0;
    else
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_emitted <= (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_r ? 2'd0 :
                                                                                                                                 f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intgo_14_done);
  
  /* buf (Ty MyDTInt_Bool) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1,MyDTInt_Bool) > (is_zae6_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_r = ((! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d <= 1'd0;
    else
      if (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_r)
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_d;
  MyDTInt_Bool_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_r = (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf[0]);
  assign is_zae6_1_1_argbuf_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf :
                                 f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf <= 1'd0;
    else
      if ((is_zae6_1_1_argbuf_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf <= 1'd0;
      else if (((! is_zae6_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_buf <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intis_zae6_1_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1,Pointer_MaskQTree) > (m1ae3_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_r = ((! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_r)
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_d;
  Pointer_MaskQTree_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_r = (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf[0]);
  assign m1ae3_1_1_argbuf_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m1ae3_1_1_argbuf_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m1ae3_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_buf <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm1ae3_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1,Pointer_QTree_Int) > (m2ae4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_r = ((! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_r)
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_d;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_r = (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf[0]);
  assign m2ae4_1_1_argbuf_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m2ae4_1_1_argbuf_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m2ae4_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_buf <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm2ae4_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1,Pointer_QTree_Int) > (m3ae5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_r = ((! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d <= {16'd0,
                                                                                                                                     1'd0};
    else
      if (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_r)
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_d;
  Pointer_QTree_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_r = (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf[0]);
  assign m3ae5_1_1_argbuf_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf :
                               f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf <= {16'd0,
                                                                                                                                       1'd0};
    else
      if ((m3ae5_1_1_argbuf_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf <= {16'd0,
                                                                                                                                         1'd0};
      else if (((! m3ae5_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_buf <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intm3ae5_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1,MyDTInt_Int_Int) > (op_addae7_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d;
  logic f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_r;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_r = ((! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d[0]) || f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d <= 1'd0;
    else
      if (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_r)
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_d;
  MyDTInt_Int_Int_t f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf;
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_r = (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf[0]);
  assign op_addae7_1_1_argbuf_d = (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf[0] ? f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf :
                                   f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf <= 1'd0;
    else
      if ((op_addae7_1_1_argbuf_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf[0]))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf <= 1'd0;
      else if (((! op_addae7_1_1_argbuf_r) && (! f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf[0])))
        f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_buf <= f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Intop_addae7_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_resbuf_bufchan_d;
  logic f_f_Int_resbuf_bufchan_r;
  assign f_f_Int_resbuf_r = ((! f_f_Int_resbuf_bufchan_d[0]) || f_f_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (f_f_Int_resbuf_r) f_f_Int_resbuf_bufchan_d <= f_f_Int_resbuf_d;
  Pointer_QTree_Int_t f_f_Int_resbuf_bufchan_buf;
  assign f_f_Int_resbuf_bufchan_r = (! f_f_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (f_f_Int_resbuf_bufchan_buf[0] ? f_f_Int_resbuf_bufchan_buf :
                            f_f_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_f_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && f_f_Int_resbuf_bufchan_buf[0]))
        f_f_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! f_f_Int_resbuf_bufchan_buf[0])))
        f_f_Int_resbuf_bufchan_buf <= f_f_Int_resbuf_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c+) : [(go_1,Go)] > (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) */
  assign \go_1Dcon_$fNumInt_$c+_d  = \Dcon_$fNumInt_$c+_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_$fNumInt_$c+_r  && \go_1Dcon_$fNumInt_$c+_d [0])}};
  
  /* fork (Ty C5) : (go_10_goMux_choice,C5) > [(go_10_goMux_choice_1,C5),
                                          (go_10_goMux_choice_2,C5),
                                          (go_10_goMux_choice_3,C5),
                                          (go_10_goMux_choice_4,C5),
                                          (go_10_goMux_choice_5,C5)] */
  logic [4:0] go_10_goMux_choice_emitted;
  logic [4:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_3_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[2]))};
  assign go_10_goMux_choice_4_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[3]))};
  assign go_10_goMux_choice_5_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[4]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_5_d[0],
                                                                   go_10_goMux_choice_4_d[0],
                                                                   go_10_goMux_choice_3_d[0],
                                                                   go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_5_r,
                                                                                                 go_10_goMux_choice_4_r,
                                                                                                 go_10_goMux_choice_3_r,
                                                                                                 go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 5'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 5'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C5) [(call_f'_f'_Int_goMux2,Pointer_QTree_Int),
                                                        (q3aeT_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2aeS_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1aeR_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m2aeH_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2aeH_goMux_mux_mux;
  logic [4:0] m2aeH_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[3:1])
      3'd0:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd1,
                                                         \call_f'_f'_Int_goMux2_d };
      3'd1:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd2,
                                                         q3aeT_1_1_argbuf_d};
      3'd2:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd4,
                                                         q2aeS_2_1_argbuf_d};
      3'd3:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd8,
                                                         q1aeR_3_1_argbuf_d};
      3'd4:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd16,
                                                         lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_d};
      default:
        {m2aeH_goMux_mux_onehot, m2aeH_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2aeH_goMux_mux_d = {m2aeH_goMux_mux_mux[16:1],
                              (m2aeH_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (m2aeH_goMux_mux_d[0] && m2aeH_goMux_mux_r);
  assign {lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_r,
          q1aeR_3_1_argbuf_r,
          q2aeS_2_1_argbuf_r,
          q3aeT_1_1_argbuf_r,
          \call_f'_f'_Int_goMux2_r } = (go_10_goMux_choice_1_r ? m2aeH_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_2,C5) [(call_f'_f'_Int_goMux3,Pointer_QTree_Int),
                                                        (t3aeY_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2aeX_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1aeW_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4aeZ_1_argbuf,Pointer_QTree_Int)] > (m3aeI_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m3aeI_goMux_mux_mux;
  logic [4:0] m3aeI_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[3:1])
      3'd0:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd1,
                                                         \call_f'_f'_Int_goMux3_d };
      3'd1:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd2,
                                                         t3aeY_1_1_argbuf_d};
      3'd2:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd4,
                                                         t2aeX_2_1_argbuf_d};
      3'd3:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd8,
                                                         t1aeW_3_1_argbuf_d};
      3'd4:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd16,
                                                         t4aeZ_1_argbuf_d};
      default:
        {m3aeI_goMux_mux_onehot, m3aeI_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3aeI_goMux_mux_d = {m3aeI_goMux_mux_mux[16:1],
                              (m3aeI_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (m3aeI_goMux_mux_d[0] && m3aeI_goMux_mux_r);
  assign {t4aeZ_1_argbuf_r,
          t1aeW_3_1_argbuf_r,
          t2aeX_2_1_argbuf_r,
          t3aeY_1_1_argbuf_r,
          \call_f'_f'_Int_goMux3_r } = (go_10_goMux_choice_2_r ? m3aeI_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_10_goMux_choice_3,C5) [(call_f'_f'_Int_goMux4,MyDTInt_Bool),
                                                   (is_zaeJ_2_2_argbuf,MyDTInt_Bool),
                                                   (is_zaeJ_3_2_argbuf,MyDTInt_Bool),
                                                   (is_zaeJ_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_zaeJ_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_zaeJ_goMux_mux_mux;
  logic [4:0] is_zaeJ_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_3_d[3:1])
      3'd0:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd1,
                                                             \call_f'_f'_Int_goMux4_d };
      3'd1:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd2,
                                                             is_zaeJ_2_2_argbuf_d};
      3'd2:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd4,
                                                             is_zaeJ_3_2_argbuf_d};
      3'd3:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd8,
                                                             is_zaeJ_4_1_argbuf_d};
      3'd4:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd16,
                                                             lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_d};
      default:
        {is_zaeJ_goMux_mux_onehot, is_zaeJ_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_zaeJ_goMux_mux_d = (is_zaeJ_goMux_mux_mux[0] && go_10_goMux_choice_3_d[0]);
  assign go_10_goMux_choice_3_r = (is_zaeJ_goMux_mux_d[0] && is_zaeJ_goMux_mux_r);
  assign {lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_r,
          is_zaeJ_4_1_argbuf_r,
          is_zaeJ_3_2_argbuf_r,
          is_zaeJ_2_2_argbuf_r,
          \call_f'_f'_Int_goMux4_r } = (go_10_goMux_choice_3_r ? is_zaeJ_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_10_goMux_choice_4,C5) [(call_f'_f'_Int_goMux5,MyDTInt_Int_Int),
                                                      (op_addaeK_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addaeK_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addaeK_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_addaeK_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_addaeK_goMux_mux_mux;
  logic [4:0] op_addaeK_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_4_d[3:1])
      3'd0:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd1,
                                                                 \call_f'_f'_Int_goMux5_d };
      3'd1:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd2,
                                                                 op_addaeK_2_2_argbuf_d};
      3'd2:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd4,
                                                                 op_addaeK_3_2_argbuf_d};
      3'd3:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd8,
                                                                 op_addaeK_4_1_argbuf_d};
      3'd4:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_d};
      default:
        {op_addaeK_goMux_mux_onehot, op_addaeK_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_addaeK_goMux_mux_d = (op_addaeK_goMux_mux_mux[0] && go_10_goMux_choice_4_d[0]);
  assign go_10_goMux_choice_4_r = (op_addaeK_goMux_mux_d[0] && op_addaeK_goMux_mux_r);
  assign {lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_r,
          op_addaeK_4_1_argbuf_r,
          op_addaeK_3_2_argbuf_r,
          op_addaeK_2_2_argbuf_r,
          \call_f'_f'_Int_goMux5_r } = (go_10_goMux_choice_4_r ? op_addaeK_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf'_f'_Int) : (go_10_goMux_choice_5,C5) [(call_f'_f'_Int_goMux6,Pointer_CTf'_f'_Int),
                                                          (sca2_2_1_argbuf,Pointer_CTf'_f'_Int),
                                                          (sca1_2_1_argbuf,Pointer_CTf'_f'_Int),
                                                          (sca0_2_1_argbuf,Pointer_CTf'_f'_Int),
                                                          (sca3_2_1_argbuf,Pointer_CTf'_f'_Int)] > (sc_0_2_goMux_mux,Pointer_CTf'_f'_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_f'_f'_Int_goMux6_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_10_goMux_choice_5_d[0])};
  assign go_10_goMux_choice_5_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_f'_f'_Int_goMux6_r } = (go_10_goMux_choice_5_r ? sc_0_2_goMux_mux_onehot :
                                        5'd0);
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5),
                                          (go_11_goMux_choice_3,C5),
                                          (go_11_goMux_choice_4,C5),
                                          (go_11_goMux_choice_5,C5),
                                          (go_11_goMux_choice_6,C5)] */
  logic [5:0] go_11_goMux_choice_emitted;
  logic [5:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_3_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[2]))};
  assign go_11_goMux_choice_4_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[3]))};
  assign go_11_goMux_choice_5_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[4]))};
  assign go_11_goMux_choice_6_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[5]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_6_d[0],
                                                                   go_11_goMux_choice_5_d[0],
                                                                   go_11_goMux_choice_4_d[0],
                                                                   go_11_goMux_choice_3_d[0],
                                                                   go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_6_r,
                                                                                                 go_11_goMux_choice_5_r,
                                                                                                 go_11_goMux_choice_4_r,
                                                                                                 go_11_goMux_choice_3_r,
                                                                                                 go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 6'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 6'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_11_goMux_choice_1,C5) [(call_f_f_Int_goMux2,Pointer_MaskQTree),
                                                        (q3aea_1_1_argbuf,Pointer_MaskQTree),
                                                        (q2ae9_2_1_argbuf,Pointer_MaskQTree),
                                                        (q1ae8_3_1_argbuf,Pointer_MaskQTree),
                                                        (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf,Pointer_MaskQTree)] > (m1ae3_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] m1ae3_goMux_mux_mux;
  logic [4:0] m1ae3_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux2_d};
      3'd1:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd2,
                                                         q3aea_1_1_argbuf_d};
      3'd2:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd4,
                                                         q2ae9_2_1_argbuf_d};
      3'd3:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd8,
                                                         q1ae8_3_1_argbuf_d};
      3'd4:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd16,
                                                         lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_d};
      default:
        {m1ae3_goMux_mux_onehot, m1ae3_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1ae3_goMux_mux_d = {m1ae3_goMux_mux_mux[16:1],
                              (m1ae3_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (m1ae3_goMux_mux_d[0] && m1ae3_goMux_mux_r);
  assign {lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_r,
          q1ae8_3_1_argbuf_r,
          q2ae9_2_1_argbuf_r,
          q3aea_1_1_argbuf_r,
          call_f_f_Int_goMux2_r} = (go_11_goMux_choice_1_r ? m1ae3_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_2,C5) [(call_f_f_Int_goMux3,Pointer_QTree_Int),
                                                        (q3'aep_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2'aeo_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1'aen_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf,Pointer_QTree_Int)] > (m2ae4_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2ae4_goMux_mux_mux;
  logic [4:0] m2ae4_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux3_d};
      3'd1:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd2,
                                                         \q3'aep_1_1_argbuf_d };
      3'd2:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd4,
                                                         \q2'aeo_2_1_argbuf_d };
      3'd3:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd8,
                                                         \q1'aen_3_1_argbuf_d };
      3'd4:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd16,
                                                         lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_d};
      default:
        {m2ae4_goMux_mux_onehot, m2ae4_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ae4_goMux_mux_d = {m2ae4_goMux_mux_mux[16:1],
                              (m2ae4_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (m2ae4_goMux_mux_d[0] && m2ae4_goMux_mux_r);
  assign {lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_r,
          \q1'aen_3_1_argbuf_r ,
          \q2'aeo_2_1_argbuf_r ,
          \q3'aep_1_1_argbuf_r ,
          call_f_f_Int_goMux3_r} = (go_11_goMux_choice_2_r ? m2ae4_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_3,C5) [(call_f_f_Int_goMux4,Pointer_QTree_Int),
                                                        (t3aeu_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2aet_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1aes_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4aev_1_argbuf,Pointer_QTree_Int)] > (m3ae5_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m3ae5_goMux_mux_mux;
  logic [4:0] m3ae5_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_3_d[3:1])
      3'd0:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_goMux4_d};
      3'd1:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd2,
                                                         t3aeu_1_1_argbuf_d};
      3'd2:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd4,
                                                         t2aet_2_1_argbuf_d};
      3'd3:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd8,
                                                         t1aes_3_1_argbuf_d};
      3'd4:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd16,
                                                         t4aev_1_argbuf_d};
      default:
        {m3ae5_goMux_mux_onehot, m3ae5_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m3ae5_goMux_mux_d = {m3ae5_goMux_mux_mux[16:1],
                              (m3ae5_goMux_mux_mux[0] && go_11_goMux_choice_3_d[0])};
  assign go_11_goMux_choice_3_r = (m3ae5_goMux_mux_d[0] && m3ae5_goMux_mux_r);
  assign {t4aev_1_argbuf_r,
          t1aes_3_1_argbuf_r,
          t2aet_2_1_argbuf_r,
          t3aeu_1_1_argbuf_r,
          call_f_f_Int_goMux4_r} = (go_11_goMux_choice_3_r ? m3ae5_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_11_goMux_choice_4,C5) [(call_f_f_Int_goMux5,MyDTInt_Bool),
                                                   (is_zae6_2_2_argbuf,MyDTInt_Bool),
                                                   (is_zae6_3_2_argbuf,MyDTInt_Bool),
                                                   (is_zae6_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_zae6_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_zae6_goMux_mux_mux;
  logic [4:0] is_zae6_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_4_d[3:1])
      3'd0:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd1,
                                                             call_f_f_Int_goMux5_d};
      3'd1:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd2,
                                                             is_zae6_2_2_argbuf_d};
      3'd2:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd4,
                                                             is_zae6_3_2_argbuf_d};
      3'd3:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd8,
                                                             is_zae6_4_1_argbuf_d};
      3'd4:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd16,
                                                             lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_d};
      default:
        {is_zae6_goMux_mux_onehot, is_zae6_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_zae6_goMux_mux_d = (is_zae6_goMux_mux_mux[0] && go_11_goMux_choice_4_d[0]);
  assign go_11_goMux_choice_4_r = (is_zae6_goMux_mux_d[0] && is_zae6_goMux_mux_r);
  assign {lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_r,
          is_zae6_4_1_argbuf_r,
          is_zae6_3_2_argbuf_r,
          is_zae6_2_2_argbuf_r,
          call_f_f_Int_goMux5_r} = (go_11_goMux_choice_4_r ? is_zae6_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_11_goMux_choice_5,C5) [(call_f_f_Int_goMux6,MyDTInt_Int_Int),
                                                      (op_addae7_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addae7_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_addae7_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_addae7_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_addae7_goMux_mux_mux;
  logic [4:0] op_addae7_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_5_d[3:1])
      3'd0:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd1,
                                                                 call_f_f_Int_goMux6_d};
      3'd1:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd2,
                                                                 op_addae7_2_2_argbuf_d};
      3'd2:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd4,
                                                                 op_addae7_3_2_argbuf_d};
      3'd3:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd8,
                                                                 op_addae7_4_1_argbuf_d};
      3'd4:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd16,
                                                                 lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_d};
      default:
        {op_addae7_goMux_mux_onehot, op_addae7_goMux_mux_mux} = {5'd0,
                                                                 1'd0};
    endcase
  assign op_addae7_goMux_mux_d = (op_addae7_goMux_mux_mux[0] && go_11_goMux_choice_5_d[0]);
  assign go_11_goMux_choice_5_r = (op_addae7_goMux_mux_d[0] && op_addae7_goMux_mux_r);
  assign {lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_r,
          op_addae7_4_1_argbuf_r,
          op_addae7_3_2_argbuf_r,
          op_addae7_2_2_argbuf_r,
          call_f_f_Int_goMux6_r} = (go_11_goMux_choice_5_r ? op_addae7_goMux_mux_onehot :
                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf_f_Int) : (go_11_goMux_choice_6,C5) [(call_f_f_Int_goMux7,Pointer_CTf_f_Int),
                                                        (sca2_3_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca1_3_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca0_3_1_argbuf,Pointer_CTf_f_Int),
                                                        (sca3_3_1_argbuf,Pointer_CTf_f_Int)] > (sc_0_3_goMux_mux,Pointer_CTf_f_Int) */
  logic [16:0] sc_0_3_goMux_mux_mux;
  logic [4:0] sc_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_6_d[3:1])
      3'd0:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd1,
                                                           call_f_f_Int_goMux7_d};
      3'd1:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd2,
                                                           sca2_3_1_argbuf_d};
      3'd2:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd4,
                                                           sca1_3_1_argbuf_d};
      3'd3:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd8,
                                                           sca0_3_1_argbuf_d};
      3'd4:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd16,
                                                           sca3_3_1_argbuf_d};
      default:
        {sc_0_3_goMux_mux_onehot, sc_0_3_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_3_goMux_mux_d = {sc_0_3_goMux_mux_mux[16:1],
                               (sc_0_3_goMux_mux_mux[0] && go_11_goMux_choice_6_d[0])};
  assign go_11_goMux_choice_6_r = (sc_0_3_goMux_mux_d[0] && sc_0_3_goMux_mux_r);
  assign {sca3_3_1_argbuf_r,
          sca0_3_1_argbuf_r,
          sca1_3_1_argbuf_r,
          sca2_3_1_argbuf_r,
          call_f_f_Int_goMux7_r} = (go_11_goMux_choice_6_r ? sc_0_3_goMux_mux_onehot :
                                    5'd0);
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Int,
      Dcon Lf'''''''''_f'''''''''_Intsbos) : [(go_12_1,Go)] > (go_12_1Lf'''''''''_f'''''''''_Intsbos,CTf'''''''''_f'''''''''_Int) */
  assign \go_12_1Lf'''''''''_f'''''''''_Intsbos_d  = \Lf'''''''''_f'''''''''_Intsbos_dc ((& {go_12_1_d[0]}), go_12_1_d);
  assign {go_12_1_r} = {1 {(\go_12_1Lf'''''''''_f'''''''''_Intsbos_r  && \go_12_1Lf'''''''''_f'''''''''_Intsbos_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (go_12_1Lf'''''''''_f'''''''''_Intsbos,CTf'''''''''_f'''''''''_Int) > (lizzieLet43_1_argbuf,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d ;
  logic \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_r ;
  assign \go_12_1Lf'''''''''_f'''''''''_Intsbos_r  = ((! \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d [0]) || \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d  <= {115'd0,
                                                            1'd0};
    else
      if (\go_12_1Lf'''''''''_f'''''''''_Intsbos_r )
        \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d  <= \go_12_1Lf'''''''''_f'''''''''_Intsbos_d ;
  \CTf'''''''''_f'''''''''_Int_t  \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf ;
  assign \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_r  = (! \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf [0]);
  assign lizzieLet43_1_argbuf_d = (\go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf [0] ? \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf  :
                                   \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf  <= {115'd0,
                                                              1'd0};
    else
      if ((lizzieLet43_1_argbuf_r && \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf [0]))
        \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf  <= {115'd0,
                                                                1'd0};
      else if (((! lizzieLet43_1_argbuf_r) && (! \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf [0])))
        \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_buf  <= \go_12_1Lf'''''''''_f'''''''''_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_12_2,Go) > (go_12_2_argbuf,Go) */
  Go_t go_12_2_bufchan_d;
  logic go_12_2_bufchan_r;
  assign go_12_2_r = ((! go_12_2_bufchan_d[0]) || go_12_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_d <= 1'd0;
    else if (go_12_2_r) go_12_2_bufchan_d <= go_12_2_d;
  Go_t go_12_2_bufchan_buf;
  assign go_12_2_bufchan_r = (! go_12_2_bufchan_buf[0]);
  assign go_12_2_argbuf_d = (go_12_2_bufchan_buf[0] ? go_12_2_bufchan_buf :
                             go_12_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_buf <= 1'd0;
    else
      if ((go_12_2_argbuf_r && go_12_2_bufchan_buf[0]))
        go_12_2_bufchan_buf <= 1'd0;
      else if (((! go_12_2_argbuf_r) && (! go_12_2_bufchan_buf[0])))
        go_12_2_bufchan_buf <= go_12_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int) : [(go_12_2_argbuf,Go),
                                                                                                   (q4aew_1_1_argbuf,Pointer_MaskQTree),
                                                                                                   (q4'aex_1_1_argbuf,Pointer_QTree_Int),
                                                                                                   (lizzieLet4_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int)] > (call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int) */
  assign \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d  = \TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_dc ((& {go_12_2_argbuf_d[0],
                                                                                                                                                                                                                                q4aew_1_1_argbuf_d[0],
                                                                                                                                                                                                                                \q4'aex_1_1_argbuf_d [0],
                                                                                                                                                                                                                                lizzieLet4_1_1_argbuf_d[0]}), go_12_2_argbuf_d, q4aew_1_1_argbuf_d, \q4'aex_1_1_argbuf_d , lizzieLet4_1_1_argbuf_d);
  assign {go_12_2_argbuf_r,
          q4aew_1_1_argbuf_r,
          \q4'aex_1_1_argbuf_r ,
          lizzieLet4_1_1_argbuf_r} = {4 {(\call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_r  && \call_f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_CTf'''''''''_f'''''''''_Int_1_d [0])}};
  
  /* dcon (Ty CTf'_f'_Int,
      Dcon Lf'_f'_Intsbos) : [(go_13_1,Go)] > (go_13_1Lf'_f'_Intsbos,CTf'_f'_Int) */
  assign \go_13_1Lf'_f'_Intsbos_d  = \Lf'_f'_Intsbos_dc ((& {go_13_1_d[0]}), go_13_1_d);
  assign {go_13_1_r} = {1 {(\go_13_1Lf'_f'_Intsbos_r  && \go_13_1Lf'_f'_Intsbos_d [0])}};
  
  /* buf (Ty CTf'_f'_Int) : (go_13_1Lf'_f'_Intsbos,CTf'_f'_Int) > (lizzieLet44_1_argbuf,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \go_13_1Lf'_f'_Intsbos_bufchan_d ;
  logic \go_13_1Lf'_f'_Intsbos_bufchan_r ;
  assign \go_13_1Lf'_f'_Intsbos_r  = ((! \go_13_1Lf'_f'_Intsbos_bufchan_d [0]) || \go_13_1Lf'_f'_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf'_f'_Intsbos_bufchan_d  <= {115'd0, 1'd0};
    else
      if (\go_13_1Lf'_f'_Intsbos_r )
        \go_13_1Lf'_f'_Intsbos_bufchan_d  <= \go_13_1Lf'_f'_Intsbos_d ;
  \CTf'_f'_Int_t  \go_13_1Lf'_f'_Intsbos_bufchan_buf ;
  assign \go_13_1Lf'_f'_Intsbos_bufchan_r  = (! \go_13_1Lf'_f'_Intsbos_bufchan_buf [0]);
  assign lizzieLet44_1_argbuf_d = (\go_13_1Lf'_f'_Intsbos_bufchan_buf [0] ? \go_13_1Lf'_f'_Intsbos_bufchan_buf  :
                                   \go_13_1Lf'_f'_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf'_f'_Intsbos_bufchan_buf  <= {115'd0, 1'd0};
    else
      if ((lizzieLet44_1_argbuf_r && \go_13_1Lf'_f'_Intsbos_bufchan_buf [0]))
        \go_13_1Lf'_f'_Intsbos_bufchan_buf  <= {115'd0, 1'd0};
      else if (((! lizzieLet44_1_argbuf_r) && (! \go_13_1Lf'_f'_Intsbos_bufchan_buf [0])))
        \go_13_1Lf'_f'_Intsbos_bufchan_buf  <= \go_13_1Lf'_f'_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_13_2,Go) > (go_13_2_argbuf,Go) */
  Go_t go_13_2_bufchan_d;
  logic go_13_2_bufchan_r;
  assign go_13_2_r = ((! go_13_2_bufchan_d[0]) || go_13_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_d <= 1'd0;
    else if (go_13_2_r) go_13_2_bufchan_d <= go_13_2_d;
  Go_t go_13_2_bufchan_buf;
  assign go_13_2_bufchan_r = (! go_13_2_bufchan_buf[0]);
  assign go_13_2_argbuf_d = (go_13_2_bufchan_buf[0] ? go_13_2_bufchan_buf :
                             go_13_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_buf <= 1'd0;
    else
      if ((go_13_2_argbuf_r && go_13_2_bufchan_buf[0]))
        go_13_2_bufchan_buf <= 1'd0;
      else if (((! go_13_2_argbuf_r) && (! go_13_2_bufchan_buf[0])))
        go_13_2_bufchan_buf <= go_13_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int) : [(go_13_2_argbuf,Go),
                                                                                                                    (m2aeH_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                    (m3aeI_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                    (is_zaeJ_1_1_argbuf,MyDTInt_Bool),
                                                                                                                    (op_addaeK_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                    (lizzieLet12_1_1_argbuf,Pointer_CTf'_f'_Int)] > (call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int) */
  assign \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d  = \TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_dc ((& {go_13_2_argbuf_d[0],
                                                                                                                                                                                                                                                  m2aeH_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                  m3aeI_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                  is_zaeJ_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                  op_addaeK_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                  lizzieLet12_1_1_argbuf_d[0]}), go_13_2_argbuf_d, m2aeH_1_1_argbuf_d, m3aeI_1_1_argbuf_d, is_zaeJ_1_1_argbuf_d, op_addaeK_1_1_argbuf_d, lizzieLet12_1_1_argbuf_d);
  assign {go_13_2_argbuf_r,
          m2aeH_1_1_argbuf_r,
          m3aeI_1_1_argbuf_r,
          is_zaeJ_1_1_argbuf_r,
          op_addaeK_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r} = {6 {(\call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_r  && \call_f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf'_f'_Int_1_d [0])}};
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lf_f_Intsbos) : [(go_14_1,Go)] > (go_14_1Lf_f_Intsbos,CTf_f_Int) */
  assign go_14_1Lf_f_Intsbos_d = Lf_f_Intsbos_dc((& {go_14_1_d[0]}), go_14_1_d);
  assign {go_14_1_r} = {1 {(go_14_1Lf_f_Intsbos_r && go_14_1Lf_f_Intsbos_d[0])}};
  
  /* buf (Ty CTf_f_Int) : (go_14_1Lf_f_Intsbos,CTf_f_Int) > (lizzieLet45_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t go_14_1Lf_f_Intsbos_bufchan_d;
  logic go_14_1Lf_f_Intsbos_bufchan_r;
  assign go_14_1Lf_f_Intsbos_r = ((! go_14_1Lf_f_Intsbos_bufchan_d[0]) || go_14_1Lf_f_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Intsbos_bufchan_d <= {163'd0, 1'd0};
    else
      if (go_14_1Lf_f_Intsbos_r)
        go_14_1Lf_f_Intsbos_bufchan_d <= go_14_1Lf_f_Intsbos_d;
  CTf_f_Int_t go_14_1Lf_f_Intsbos_bufchan_buf;
  assign go_14_1Lf_f_Intsbos_bufchan_r = (! go_14_1Lf_f_Intsbos_bufchan_buf[0]);
  assign lizzieLet45_1_argbuf_d = (go_14_1Lf_f_Intsbos_bufchan_buf[0] ? go_14_1Lf_f_Intsbos_bufchan_buf :
                                   go_14_1Lf_f_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Intsbos_bufchan_buf <= {163'd0, 1'd0};
    else
      if ((lizzieLet45_1_argbuf_r && go_14_1Lf_f_Intsbos_bufchan_buf[0]))
        go_14_1Lf_f_Intsbos_bufchan_buf <= {163'd0, 1'd0};
      else if (((! lizzieLet45_1_argbuf_r) && (! go_14_1Lf_f_Intsbos_bufchan_buf[0])))
        go_14_1Lf_f_Intsbos_bufchan_buf <= go_14_1Lf_f_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_14_2,Go) > (go_14_2_argbuf,Go) */
  Go_t go_14_2_bufchan_d;
  logic go_14_2_bufchan_r;
  assign go_14_2_r = ((! go_14_2_bufchan_d[0]) || go_14_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_d <= 1'd0;
    else if (go_14_2_r) go_14_2_bufchan_d <= go_14_2_d;
  Go_t go_14_2_bufchan_buf;
  assign go_14_2_bufchan_r = (! go_14_2_bufchan_buf[0]);
  assign go_14_2_argbuf_d = (go_14_2_bufchan_buf[0] ? go_14_2_bufchan_buf :
                             go_14_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_buf <= 1'd0;
    else
      if ((go_14_2_argbuf_r && go_14_2_bufchan_buf[0]))
        go_14_2_bufchan_buf <= 1'd0;
      else if (((! go_14_2_argbuf_r) && (! go_14_2_bufchan_buf[0])))
        go_14_2_bufchan_buf <= go_14_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) : [(go_14_2_argbuf,Go),
                                                                                                                                      (m1ae3_1_1_argbuf,Pointer_MaskQTree),
                                                                                                                                      (m2ae4_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                      (m3ae5_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                      (is_zae6_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                      (op_addae7_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                      (lizzieLet27_1_1_argbuf,Pointer_CTf_f_Int)] > (call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int) */
  assign call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d = TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_dc((& {go_14_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                m1ae3_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                m2ae4_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                m3ae5_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                is_zae6_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                op_addae7_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                lizzieLet27_1_1_argbuf_d[0]}), go_14_2_argbuf_d, m1ae3_1_1_argbuf_d, m2ae4_1_1_argbuf_d, m3ae5_1_1_argbuf_d, is_zae6_1_1_argbuf_d, op_addae7_1_1_argbuf_d, lizzieLet27_1_1_argbuf_d);
  assign {go_14_2_argbuf_r,
          m1ae3_1_1_argbuf_r,
          m2ae4_1_1_argbuf_r,
          m3ae5_1_1_argbuf_r,
          is_zae6_1_1_argbuf_r,
          op_addae7_1_1_argbuf_r,
          lizzieLet27_1_1_argbuf_r} = {7 {(call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_r && call_f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Pointer_CTf_f_Int_1_d[0])}};
  
  /* fork (Ty C4) : (go_15_goMux_choice,C4) > [(go_15_goMux_choice_1,C4),
                                          (go_15_goMux_choice_2,C4)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_15_goMux_choice_1,C4) [(lizzieLet28_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet29_1_argbuf,Int#),
                                           (lizzieLet28_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet28_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet29_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet28_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet28_1_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet28_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz_Int) : (go_15_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_7_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_7_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C6) : (go_16_goMux_choice,C6) > [(go_16_goMux_choice_1,C6),
                                          (go_16_goMux_choice_2,C6)] */
  logic [1:0] go_16_goMux_choice_emitted;
  logic [1:0] go_16_goMux_choice_done;
  assign go_16_goMux_choice_1_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[0]))};
  assign go_16_goMux_choice_2_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[1]))};
  assign go_16_goMux_choice_done = (go_16_goMux_choice_emitted | ({go_16_goMux_choice_2_d[0],
                                                                   go_16_goMux_choice_1_d[0]} & {go_16_goMux_choice_2_r,
                                                                                                 go_16_goMux_choice_1_r}));
  assign go_16_goMux_choice_r = (& go_16_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_goMux_choice_emitted <= 2'd0;
    else
      go_16_goMux_choice_emitted <= (go_16_goMux_choice_r ? 2'd0 :
                                     go_16_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Int) : (go_16_goMux_choice_1,C6) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet6_5MQVal_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [5:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet6_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_1_d[0])};
  assign go_16_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet6_5MQVal_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_16_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTf'''''''''_f'''''''''_Int) : (go_16_goMux_choice_2,C6) [(lizzieLet6_6MQNone_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                          (sc_0_11_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                          (lizzieLet6_6MQVal_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                          (lizzieLet6_4MQNode_4QNone_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                          (lizzieLet6_4MQNode_4QVal_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                          (lizzieLet6_4MQNode_4QError_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [5:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet6_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   sc_0_11_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet6_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet6_4MQNode_4QNone_Int_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet6_4MQNode_4QVal_Int_1_argbuf_d};
      3'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet6_4MQNode_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_2_d[0])};
  assign go_16_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_4MQNode_4QError_Int_1_argbuf_r,
          lizzieLet6_4MQNode_4QVal_Int_1_argbuf_r,
          lizzieLet6_4MQNode_4QNone_Int_1_argbuf_r,
          lizzieLet6_6MQVal_1_argbuf_r,
          sc_0_11_1_argbuf_r,
          lizzieLet6_6MQNone_1_argbuf_r} = (go_16_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                            6'd0);
  
  /* fork (Ty C11) : (go_17_goMux_choice,C11) > [(go_17_goMux_choice_1,C11),
                                            (go_17_goMux_choice_2,C11)] */
  logic [1:0] go_17_goMux_choice_emitted;
  logic [1:0] go_17_goMux_choice_done;
  assign go_17_goMux_choice_1_d = {go_17_goMux_choice_d[4:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[0]))};
  assign go_17_goMux_choice_2_d = {go_17_goMux_choice_d[4:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[1]))};
  assign go_17_goMux_choice_done = (go_17_goMux_choice_emitted | ({go_17_goMux_choice_2_d[0],
                                                                   go_17_goMux_choice_1_d[0]} & {go_17_goMux_choice_2_r,
                                                                                                 go_17_goMux_choice_1_r}));
  assign go_17_goMux_choice_r = (& go_17_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_goMux_choice_emitted <= 2'd0;
    else
      go_17_goMux_choice_emitted <= (go_17_goMux_choice_r ? 2'd0 :
                                     go_17_goMux_choice_done);
  
  /* mux (Ty C11,
     Ty Pointer_QTree_Int) : (go_17_goMux_choice_1,C11) [(lizzieLet13_7QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet5_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet6_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet9_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet10_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet11_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [10:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd1,
                                                                   lizzieLet13_7QNone_Int_1_argbuf_d};
      4'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd2,
                                                                   contRet_0_2_1_argbuf_d};
      4'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd4,
                                                                   lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_d};
      4'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd8,
                                                                   lizzieLet5_1_1_argbuf_d};
      4'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd16,
                                                                   lizzieLet6_1_1_argbuf_d};
      4'd5:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd32,
                                                                   lizzieLet7_1_1_argbuf_d};
      4'd6:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd64,
                                                                   lizzieLet8_1_1_argbuf_d};
      4'd7:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd128,
                                                                   lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_d};
      4'd8:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd256,
                                                                   lizzieLet9_1_1_argbuf_d};
      4'd9:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd512,
                                                                   lizzieLet10_1_1_argbuf_d};
      4'd10:
        {srtarg_0_2_goMux_mux_onehot,
         srtarg_0_2_goMux_mux_mux} = {11'd1024, lizzieLet11_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {11'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_1_d[0])};
  assign go_17_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet11_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r,
          lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet13_7QNone_Int_1_argbuf_r} = (go_17_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                                11'd0);
  
  /* mux (Ty C11,
     Ty Pointer_CTf'_f'_Int) : (go_17_goMux_choice_2,C11) [(lizzieLet13_9QNone_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (sc_0_15_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (es_2_3MyFalse_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (es_2_3MyTrue_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QVal_Int_7QError_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_5QNode_Int_7QError_Int_1_argbuf,Pointer_CTf'_f'_Int),
                                                           (lizzieLet13_9QError_Int_1_argbuf,Pointer_CTf'_f'_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTf'_f'_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [10:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd1,
                                                                   lizzieLet13_9QNone_Int_1_argbuf_d};
      4'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd2,
                                                                   sc_0_15_1_argbuf_d};
      4'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd4,
                                                                   lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_d};
      4'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd8,
                                                                   es_2_3MyFalse_1_argbuf_d};
      4'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd16,
                                                                   es_2_3MyTrue_1_argbuf_d};
      4'd5:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd32,
                                                                   lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd64,
                                                                   lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_d};
      4'd7:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd128,
                                                                   lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_d};
      4'd8:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd256,
                                                                   lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_d};
      4'd9:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd512,
                                                                   lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_d};
      4'd10:
        {scfarg_0_2_goMux_mux_onehot,
         scfarg_0_2_goMux_mux_mux} = {11'd1024,
                                      lizzieLet13_9QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {11'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_2_d[0])};
  assign go_17_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet13_9QError_Int_1_argbuf_r,
          lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_r,
          lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_r,
          lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_r,
          lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_r,
          lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_r,
          es_2_3MyTrue_1_argbuf_r,
          es_2_3MyFalse_1_argbuf_r,
          lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_r,
          sc_0_15_1_argbuf_r,
          lizzieLet13_9QNone_Int_1_argbuf_r} = (go_17_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                11'd0);
  
  /* fork (Ty C16) : (go_18_goMux_choice,C16) > [(go_18_goMux_choice_1,C16),
                                            (go_18_goMux_choice_2,C16)] */
  logic [1:0] go_18_goMux_choice_emitted;
  logic [1:0] go_18_goMux_choice_done;
  assign go_18_goMux_choice_1_d = {go_18_goMux_choice_d[4:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[0]))};
  assign go_18_goMux_choice_2_d = {go_18_goMux_choice_d[4:1],
                                   (go_18_goMux_choice_d[0] && (! go_18_goMux_choice_emitted[1]))};
  assign go_18_goMux_choice_done = (go_18_goMux_choice_emitted | ({go_18_goMux_choice_2_d[0],
                                                                   go_18_goMux_choice_1_d[0]} & {go_18_goMux_choice_2_r,
                                                                                                 go_18_goMux_choice_1_r}));
  assign go_18_goMux_choice_r = (& go_18_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_18_goMux_choice_emitted <= 2'd0;
    else
      go_18_goMux_choice_emitted <= (go_18_goMux_choice_r ? 2'd0 :
                                     go_18_goMux_choice_done);
  
  /* mux (Ty C16,
     Ty Pointer_QTree_Int) : (go_18_goMux_choice_1,C16) [(lizzieLet13_1_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_3_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet14_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet15_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet16_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet17_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet18_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet19_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet20_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet21_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet22_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet19_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet23_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet24_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet25_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet26_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_3_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_3_goMux_mux_mux;
  logic [15:0] srtarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd1,
                                                                   lizzieLet13_1_1_argbuf_d};
      4'd1:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd2,
                                                                   contRet_0_3_1_argbuf_d};
      4'd2:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd4,
                                                                   lizzieLet14_1_1_argbuf_d};
      4'd3:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd8,
                                                                   lizzieLet15_1_1_argbuf_d};
      4'd4:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd16,
                                                                   lizzieLet16_1_1_argbuf_d};
      4'd5:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd32,
                                                                   lizzieLet17_1_1_argbuf_d};
      4'd6:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd64,
                                                                   lizzieLet18_1_1_argbuf_d};
      4'd7:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd128,
                                                                   lizzieLet19_1_argbuf_d};
      4'd8:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd256,
                                                                   lizzieLet20_1_1_argbuf_d};
      4'd9:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd512,
                                                                   lizzieLet21_1_1_argbuf_d};
      4'd10:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd1024, lizzieLet22_1_1_argbuf_d};
      4'd11:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd2048, lizzieLet19_1_1_argbuf_d};
      4'd12:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd4096, lizzieLet23_1_1_argbuf_d};
      4'd13:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd8192, lizzieLet24_1_1_argbuf_d};
      4'd14:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd16384, lizzieLet25_1_1_argbuf_d};
      4'd15:
        {srtarg_0_3_goMux_mux_onehot,
         srtarg_0_3_goMux_mux_mux} = {16'd32768, lizzieLet26_1_1_argbuf_d};
      default:
        {srtarg_0_3_goMux_mux_onehot, srtarg_0_3_goMux_mux_mux} = {16'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_3_goMux_mux_d = {srtarg_0_3_goMux_mux_mux[16:1],
                                   (srtarg_0_3_goMux_mux_mux[0] && go_18_goMux_choice_1_d[0])};
  assign go_18_goMux_choice_1_r = (srtarg_0_3_goMux_mux_d[0] && srtarg_0_3_goMux_mux_r);
  assign {lizzieLet26_1_1_argbuf_r,
          lizzieLet25_1_1_argbuf_r,
          lizzieLet24_1_1_argbuf_r,
          lizzieLet23_1_1_argbuf_r,
          lizzieLet19_1_1_argbuf_r,
          lizzieLet22_1_1_argbuf_r,
          lizzieLet21_1_1_argbuf_r,
          lizzieLet20_1_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_1_argbuf_r,
          lizzieLet17_1_1_argbuf_r,
          lizzieLet16_1_1_argbuf_r,
          lizzieLet15_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r,
          contRet_0_3_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r} = (go_18_goMux_choice_1_r ? srtarg_0_3_goMux_mux_onehot :
                                       16'd0);
  
  /* mux (Ty C16,
     Ty Pointer_CTf_f_Int) : (go_18_goMux_choice_2,C16) [(lizzieLet24_10MQNone_1_argbuf,Pointer_CTf_f_Int),
                                                         (sc_0_19_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_10MQVal_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_6_1_1MyFalse_1_argbuf,Pointer_CTf_f_Int),
                                                         (es_6_1_1MyTrue_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int),
                                                         (lizzieLet24_5MQNode_3QError_Int_1_argbuf,Pointer_CTf_f_Int)] > (scfarg_0_3_goMux_mux,Pointer_CTf_f_Int) */
  logic [16:0] scfarg_0_3_goMux_mux_mux;
  logic [15:0] scfarg_0_3_goMux_mux_onehot;
  always_comb
    unique case (go_18_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd1,
                                                                   lizzieLet24_10MQNone_1_argbuf_d};
      4'd1:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd2,
                                                                   sc_0_19_1_argbuf_d};
      4'd2:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd4,
                                                                   lizzieLet24_10MQVal_1_argbuf_d};
      4'd3:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd8,
                                                                   lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_d};
      4'd4:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd16,
                                                                   lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_d};
      4'd5:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd32,
                                                                   lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd64,
                                                                   lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_d};
      4'd7:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd128,
                                                                   lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_d};
      4'd8:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd256,
                                                                   es_6_1_1MyFalse_1_argbuf_d};
      4'd9:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd512,
                                                                   es_6_1_1MyTrue_1_argbuf_d};
      4'd10:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd1024,
                                      lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_d};
      4'd11:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd2048,
                                      lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_d};
      4'd12:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd4096,
                                      lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_d};
      4'd13:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd8192,
                                      lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_d};
      4'd14:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd16384,
                                      lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_d};
      4'd15:
        {scfarg_0_3_goMux_mux_onehot,
         scfarg_0_3_goMux_mux_mux} = {16'd32768,
                                      lizzieLet24_5MQNode_3QError_Int_1_argbuf_d};
      default:
        {scfarg_0_3_goMux_mux_onehot, scfarg_0_3_goMux_mux_mux} = {16'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_3_goMux_mux_d = {scfarg_0_3_goMux_mux_mux[16:1],
                                   (scfarg_0_3_goMux_mux_mux[0] && go_18_goMux_choice_2_d[0])};
  assign go_18_goMux_choice_2_r = (scfarg_0_3_goMux_mux_d[0] && scfarg_0_3_goMux_mux_r);
  assign {lizzieLet24_5MQNode_3QError_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_r,
          es_6_1_1MyTrue_1_argbuf_r,
          es_6_1_1MyFalse_1_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_r,
          lizzieLet24_10MQVal_1_argbuf_r,
          sc_0_19_1_argbuf_r,
          lizzieLet24_10MQNone_1_argbuf_r} = (go_18_goMux_choice_2_r ? scfarg_0_3_goMux_mux_onehot :
                                              16'd0);
  
  /* buf (Ty MyDTInt_Int_Int) : (go_1Dcon_$fNumInt_$c+,MyDTInt_Int_Int) > (es_5_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  logic \go_1Dcon_$fNumInt_$c+_bufchan_r ;
  assign \go_1Dcon_$fNumInt_$c+_r  = ((! \go_1Dcon_$fNumInt_$c+_bufchan_d [0]) || \go_1Dcon_$fNumInt_$c+_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_$fNumInt_$c+_r )
        \go_1Dcon_$fNumInt_$c+_bufchan_d  <= \go_1Dcon_$fNumInt_$c+_d ;
  MyDTInt_Int_Int_t \go_1Dcon_$fNumInt_$c+_bufchan_buf ;
  assign \go_1Dcon_$fNumInt_$c+_bufchan_r  = (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]);
  assign es_5_1_argbuf_d = (\go_1Dcon_$fNumInt_$c+_bufchan_buf [0] ? \go_1Dcon_$fNumInt_$c+_bufchan_buf  :
                            \go_1Dcon_$fNumInt_$c+_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
    else
      if ((es_5_1_argbuf_r && \go_1Dcon_$fNumInt_$c+_bufchan_buf [0]))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
      else if (((! es_5_1_argbuf_r) && (! \go_1Dcon_$fNumInt_$c+_bufchan_buf [0])))
        \go_1Dcon_$fNumInt_$c+_bufchan_buf  <= \go_1Dcon_$fNumInt_$c+_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_main1) : [(go_2,Go)] > (go_2Dcon_main1,MyDTInt_Bool) */
  assign go_2Dcon_main1_d = Dcon_main1_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_main1_r && go_2Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_2Dcon_main1,MyDTInt_Bool) > (es_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_2Dcon_main1_bufchan_d;
  logic go_2Dcon_main1_bufchan_r;
  assign go_2Dcon_main1_r = ((! go_2Dcon_main1_bufchan_d[0]) || go_2Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_main1_r) go_2Dcon_main1_bufchan_d <= go_2Dcon_main1_d;
  MyDTInt_Bool_t go_2Dcon_main1_bufchan_buf;
  assign go_2Dcon_main1_bufchan_r = (! go_2Dcon_main1_bufchan_buf[0]);
  assign es_4_1_argbuf_d = (go_2Dcon_main1_bufchan_buf[0] ? go_2Dcon_main1_bufchan_buf :
                            go_2Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_4_1_argbuf_r && go_2Dcon_main1_bufchan_buf[0]))
        go_2Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! go_2Dcon_main1_bufchan_buf[0])))
        go_2Dcon_main1_bufchan_buf <= go_2Dcon_main1_bufchan_d;
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(go_3_argbuf,Go),
                                                                                                                  (m1a8v_0,Pointer_MaskQTree),
                                                                                                                  (m2a8w_1,Pointer_QTree_Int),
                                                                                                                  (m3a8x_2,Pointer_QTree_Int),
                                                                                                                  (es_4_1_argbuf,MyDTInt_Bool),
                                                                                                                  (es_5_1_argbuf,MyDTInt_Int_Int)] > (f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d = TupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {go_3_argbuf_d[0],
                                                                                                                                                                                                                                   m1a8v_0_d[0],
                                                                                                                                                                                                                                   m2a8w_1_d[0],
                                                                                                                                                                                                                                   m3a8x_2_d[0],
                                                                                                                                                                                                                                   es_4_1_argbuf_d[0],
                                                                                                                                                                                                                                   es_5_1_argbuf_d[0]}), go_3_argbuf_d, m1a8v_0_d, m2a8w_1_d, m3a8x_2_d, es_4_1_argbuf_d, es_5_1_argbuf_d);
  assign {go_3_argbuf_r,
          m1a8v_0_r,
          m2a8w_1_r,
          m3a8x_2_r,
          es_4_1_argbuf_r,
          es_5_1_argbuf_r} = {6 {(f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r && f_f_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_4,Go) > (go_4_argbuf,Go) */
  Go_t go_4_bufchan_d;
  logic go_4_bufchan_r;
  assign go_4_r = ((! go_4_bufchan_d[0]) || go_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_d <= 1'd0;
    else if (go_4_r) go_4_bufchan_d <= go_4_d;
  Go_t go_4_bufchan_buf;
  assign go_4_bufchan_r = (! go_4_bufchan_buf[0]);
  assign go_4_argbuf_d = (go_4_bufchan_buf[0] ? go_4_bufchan_buf :
                          go_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_bufchan_buf <= 1'd0;
    else
      if ((go_4_argbuf_r && go_4_bufchan_buf[0]))
        go_4_bufchan_buf <= 1'd0;
      else if (((! go_4_argbuf_r) && (! go_4_bufchan_buf[0])))
        go_4_bufchan_buf <= go_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_4_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_4_argbuf_d[0],
                                                                                     es_0_1_argbuf_d[0]}), go_4_argbuf_d, es_0_1_argbuf_d);
  assign {go_4_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  && \$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon L$wnnz_Intsbos) : [(go_6_1,Go)] > (go_6_1L$wnnz_Intsbos,CT$wnnz_Int) */
  assign go_6_1L$wnnz_Intsbos_d = L$wnnz_Intsbos_dc((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(go_6_1L$wnnz_Intsbos_r && go_6_1L$wnnz_Intsbos_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (go_6_1L$wnnz_Intsbos,CT$wnnz_Int) > (lizzieLet0_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_bufchan_d;
  logic go_6_1L$wnnz_Intsbos_bufchan_r;
  assign go_6_1L$wnnz_Intsbos_r = ((! go_6_1L$wnnz_Intsbos_bufchan_d[0]) || go_6_1L$wnnz_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wnnz_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_6_1L$wnnz_Intsbos_r)
        go_6_1L$wnnz_Intsbos_bufchan_d <= go_6_1L$wnnz_Intsbos_d;
  CT$wnnz_Int_t go_6_1L$wnnz_Intsbos_bufchan_buf;
  assign go_6_1L$wnnz_Intsbos_bufchan_r = (! go_6_1L$wnnz_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_6_1L$wnnz_Intsbos_bufchan_buf[0] ? go_6_1L$wnnz_Intsbos_bufchan_buf :
                                  go_6_1L$wnnz_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_6_1L$wnnz_Intsbos_bufchan_buf[0]))
        go_6_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_6_1L$wnnz_Intsbos_bufchan_buf[0])))
        go_6_1L$wnnz_Intsbos_bufchan_buf <= go_6_1L$wnnz_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : [(go_6_2_argbuf,Go),
                                                               (wsjQ_1_argbuf,Pointer_QTree_Int),
                                                               (lizzieLet30_1_argbuf,Pointer_CT$wnnz_Int)] > (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) */
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_dc((& {go_6_2_argbuf_d[0],
                                                                                                                                    wsjQ_1_argbuf_d[0],
                                                                                                                                    lizzieLet30_1_argbuf_d[0]}), go_6_2_argbuf_d, wsjQ_1_argbuf_d, lizzieLet30_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          wsjQ_1_argbuf_r,
          lizzieLet30_1_argbuf_r} = {3 {(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0])}};
  
  /* fork (Ty C5) : (go_8_goMux_choice,C5) > [(go_8_goMux_choice_1,C5),
                                         (go_8_goMux_choice_2,C5)] */
  logic [1:0] go_8_goMux_choice_emitted;
  logic [1:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 2'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 2'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_8_goMux_choice_1,C5) [(call_$wnnz_Int_goMux2,Pointer_QTree_Int),
                                                       (q2a86_1_1_argbuf,Pointer_QTree_Int),
                                                       (q3a87_2_1_argbuf,Pointer_QTree_Int),
                                                       (q4a88_3_1_argbuf,Pointer_QTree_Int),
                                                       (q1a85_1_argbuf,Pointer_QTree_Int)] > (wsjQ_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wsjQ_1_goMux_mux_mux;
  logic [4:0] wsjQ_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux2_d};
      3'd1:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd2,
                                                           q2a86_1_1_argbuf_d};
      3'd2:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd4,
                                                           q3a87_2_1_argbuf_d};
      3'd3:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd8,
                                                           q4a88_3_1_argbuf_d};
      3'd4:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd16,
                                                           q1a85_1_argbuf_d};
      default:
        {wsjQ_1_goMux_mux_onehot, wsjQ_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wsjQ_1_goMux_mux_d = {wsjQ_1_goMux_mux_mux[16:1],
                               (wsjQ_1_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (wsjQ_1_goMux_mux_d[0] && wsjQ_1_goMux_mux_r);
  assign {q1a85_1_argbuf_r,
          q4a88_3_1_argbuf_r,
          q3a87_2_1_argbuf_r,
          q2a86_1_1_argbuf_r,
          call_$wnnz_Int_goMux2_r} = (go_8_goMux_choice_1_r ? wsjQ_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz_Int) : (go_8_goMux_choice_2,C5) [(call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int),
                                                         (sca2_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca1_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca0_1_argbuf,Pointer_CT$wnnz_Int),
                                                         (sca3_1_argbuf,Pointer_CT$wnnz_Int)] > (sc_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_Int_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_Int_goMux3_r} = (go_8_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                      5'd0);
  
  /* fork (Ty C5) : (go_9_goMux_choice,C5) > [(go_9_goMux_choice_1,C5),
                                         (go_9_goMux_choice_2,C5),
                                         (go_9_goMux_choice_3,C5)] */
  logic [2:0] go_9_goMux_choice_emitted;
  logic [2:0] go_9_goMux_choice_done;
  assign go_9_goMux_choice_1_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[0]))};
  assign go_9_goMux_choice_2_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[1]))};
  assign go_9_goMux_choice_3_d = {go_9_goMux_choice_d[3:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[2]))};
  assign go_9_goMux_choice_done = (go_9_goMux_choice_emitted | ({go_9_goMux_choice_3_d[0],
                                                                 go_9_goMux_choice_2_d[0],
                                                                 go_9_goMux_choice_1_d[0]} & {go_9_goMux_choice_3_r,
                                                                                              go_9_goMux_choice_2_r,
                                                                                              go_9_goMux_choice_1_r}));
  assign go_9_goMux_choice_r = (& go_9_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_goMux_choice_emitted <= 3'd0;
    else
      go_9_goMux_choice_emitted <= (go_9_goMux_choice_r ? 3'd0 :
                                    go_9_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_9_goMux_choice_1,C5) [(call_f'''''''''_f'''''''''_Int_goMux2,Pointer_MaskQTree),
                                                       (q3aeA_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2aez_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1aey_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet6_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree)] > (q4aew_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] q4aew_goMux_mux_mux;
  logic [4:0] q4aew_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_1_d[3:1])
      3'd0:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd1,
                                                         \call_f'''''''''_f'''''''''_Int_goMux2_d };
      3'd1:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd2,
                                                         q3aeA_1_1_argbuf_d};
      3'd2:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd4,
                                                         q2aez_2_1_argbuf_d};
      3'd3:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd8,
                                                         q1aey_3_1_argbuf_d};
      3'd4:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd16,
                                                         lizzieLet6_4MQNode_8QNode_Int_1_argbuf_d};
      default:
        {q4aew_goMux_mux_onehot, q4aew_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign q4aew_goMux_mux_d = {q4aew_goMux_mux_mux[16:1],
                              (q4aew_goMux_mux_mux[0] && go_9_goMux_choice_1_d[0])};
  assign go_9_goMux_choice_1_r = (q4aew_goMux_mux_d[0] && q4aew_goMux_mux_r);
  assign {lizzieLet6_4MQNode_8QNode_Int_1_argbuf_r,
          q1aey_3_1_argbuf_r,
          q2aez_2_1_argbuf_r,
          q3aeA_1_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Int_goMux2_r } = (go_9_goMux_choice_1_r ? q4aew_goMux_mux_onehot :
                                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_9_goMux_choice_2,C5) [(call_f'''''''''_f'''''''''_Int_goMux3,Pointer_QTree_Int),
                                                       (t3aeF_1_1_argbuf,Pointer_QTree_Int),
                                                       (t2aeE_2_1_argbuf,Pointer_QTree_Int),
                                                       (t1aeD_3_1_argbuf,Pointer_QTree_Int),
                                                       (t4aeG_1_argbuf,Pointer_QTree_Int)] > (q4'aex_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] \q4'aex_goMux_mux_mux ;
  logic [4:0] \q4'aex_goMux_mux_onehot ;
  always_comb
    unique case (go_9_goMux_choice_2_d[3:1])
      3'd0:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd1,
                                                               \call_f'''''''''_f'''''''''_Int_goMux3_d };
      3'd1:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd2,
                                                               t3aeF_1_1_argbuf_d};
      3'd2:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd4,
                                                               t2aeE_2_1_argbuf_d};
      3'd3:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd8,
                                                               t1aeD_3_1_argbuf_d};
      3'd4:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd16,
                                                               t4aeG_1_argbuf_d};
      default:
        {\q4'aex_goMux_mux_onehot , \q4'aex_goMux_mux_mux } = {5'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign \q4'aex_goMux_mux_d  = {\q4'aex_goMux_mux_mux [16:1],
                                 (\q4'aex_goMux_mux_mux [0] && go_9_goMux_choice_2_d[0])};
  assign go_9_goMux_choice_2_r = (\q4'aex_goMux_mux_d [0] && \q4'aex_goMux_mux_r );
  assign {t4aeG_1_argbuf_r,
          t1aeD_3_1_argbuf_r,
          t2aeE_2_1_argbuf_r,
          t3aeF_1_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Int_goMux3_r } = (go_9_goMux_choice_2_r ? \q4'aex_goMux_mux_onehot  :
                                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf'''''''''_f'''''''''_Int) : (go_9_goMux_choice_3,C5) [(call_f'''''''''_f'''''''''_Int_goMux4,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                         (sca2_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                         (sca1_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                         (sca0_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                         (sca3_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int)] > (sc_0_1_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f'''''''''_f'''''''''_Int_goMux4_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_9_goMux_choice_3_d[0])};
  assign go_9_goMux_choice_3_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f'''''''''_f'''''''''_Int_goMux4_r } = (go_9_goMux_choice_3_r ? sc_0_1_goMux_mux_onehot :
                                                        5'd0);
  
  /* buf (Ty MyDTInt_Bool) : (is_zae6_2_2,MyDTInt_Bool) > (is_zae6_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zae6_2_2_bufchan_d;
  logic is_zae6_2_2_bufchan_r;
  assign is_zae6_2_2_r = ((! is_zae6_2_2_bufchan_d[0]) || is_zae6_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_2_2_bufchan_d <= 1'd0;
    else if (is_zae6_2_2_r) is_zae6_2_2_bufchan_d <= is_zae6_2_2_d;
  MyDTInt_Bool_t is_zae6_2_2_bufchan_buf;
  assign is_zae6_2_2_bufchan_r = (! is_zae6_2_2_bufchan_buf[0]);
  assign is_zae6_2_2_argbuf_d = (is_zae6_2_2_bufchan_buf[0] ? is_zae6_2_2_bufchan_buf :
                                 is_zae6_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_zae6_2_2_argbuf_r && is_zae6_2_2_bufchan_buf[0]))
        is_zae6_2_2_bufchan_buf <= 1'd0;
      else if (((! is_zae6_2_2_argbuf_r) && (! is_zae6_2_2_bufchan_buf[0])))
        is_zae6_2_2_bufchan_buf <= is_zae6_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zae6_2_destruct,MyDTInt_Bool) > [(is_zae6_2_1,MyDTInt_Bool),
                                                              (is_zae6_2_2,MyDTInt_Bool)] */
  logic [1:0] is_zae6_2_destruct_emitted;
  logic [1:0] is_zae6_2_destruct_done;
  assign is_zae6_2_1_d = (is_zae6_2_destruct_d[0] && (! is_zae6_2_destruct_emitted[0]));
  assign is_zae6_2_2_d = (is_zae6_2_destruct_d[0] && (! is_zae6_2_destruct_emitted[1]));
  assign is_zae6_2_destruct_done = (is_zae6_2_destruct_emitted | ({is_zae6_2_2_d[0],
                                                                   is_zae6_2_1_d[0]} & {is_zae6_2_2_r,
                                                                                        is_zae6_2_1_r}));
  assign is_zae6_2_destruct_r = (& is_zae6_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_2_destruct_emitted <= 2'd0;
    else
      is_zae6_2_destruct_emitted <= (is_zae6_2_destruct_r ? 2'd0 :
                                     is_zae6_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zae6_3_2,MyDTInt_Bool) > (is_zae6_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zae6_3_2_bufchan_d;
  logic is_zae6_3_2_bufchan_r;
  assign is_zae6_3_2_r = ((! is_zae6_3_2_bufchan_d[0]) || is_zae6_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_3_2_bufchan_d <= 1'd0;
    else if (is_zae6_3_2_r) is_zae6_3_2_bufchan_d <= is_zae6_3_2_d;
  MyDTInt_Bool_t is_zae6_3_2_bufchan_buf;
  assign is_zae6_3_2_bufchan_r = (! is_zae6_3_2_bufchan_buf[0]);
  assign is_zae6_3_2_argbuf_d = (is_zae6_3_2_bufchan_buf[0] ? is_zae6_3_2_bufchan_buf :
                                 is_zae6_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_zae6_3_2_argbuf_r && is_zae6_3_2_bufchan_buf[0]))
        is_zae6_3_2_bufchan_buf <= 1'd0;
      else if (((! is_zae6_3_2_argbuf_r) && (! is_zae6_3_2_bufchan_buf[0])))
        is_zae6_3_2_bufchan_buf <= is_zae6_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zae6_3_destruct,MyDTInt_Bool) > [(is_zae6_3_1,MyDTInt_Bool),
                                                              (is_zae6_3_2,MyDTInt_Bool)] */
  logic [1:0] is_zae6_3_destruct_emitted;
  logic [1:0] is_zae6_3_destruct_done;
  assign is_zae6_3_1_d = (is_zae6_3_destruct_d[0] && (! is_zae6_3_destruct_emitted[0]));
  assign is_zae6_3_2_d = (is_zae6_3_destruct_d[0] && (! is_zae6_3_destruct_emitted[1]));
  assign is_zae6_3_destruct_done = (is_zae6_3_destruct_emitted | ({is_zae6_3_2_d[0],
                                                                   is_zae6_3_1_d[0]} & {is_zae6_3_2_r,
                                                                                        is_zae6_3_1_r}));
  assign is_zae6_3_destruct_r = (& is_zae6_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_3_destruct_emitted <= 2'd0;
    else
      is_zae6_3_destruct_emitted <= (is_zae6_3_destruct_r ? 2'd0 :
                                     is_zae6_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zae6_4_destruct,MyDTInt_Bool) > (is_zae6_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zae6_4_destruct_bufchan_d;
  logic is_zae6_4_destruct_bufchan_r;
  assign is_zae6_4_destruct_r = ((! is_zae6_4_destruct_bufchan_d[0]) || is_zae6_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_zae6_4_destruct_r)
        is_zae6_4_destruct_bufchan_d <= is_zae6_4_destruct_d;
  MyDTInt_Bool_t is_zae6_4_destruct_bufchan_buf;
  assign is_zae6_4_destruct_bufchan_r = (! is_zae6_4_destruct_bufchan_buf[0]);
  assign is_zae6_4_1_argbuf_d = (is_zae6_4_destruct_bufchan_buf[0] ? is_zae6_4_destruct_bufchan_buf :
                                 is_zae6_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zae6_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_zae6_4_1_argbuf_r && is_zae6_4_destruct_bufchan_buf[0]))
        is_zae6_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_zae6_4_1_argbuf_r) && (! is_zae6_4_destruct_bufchan_buf[0])))
        is_zae6_4_destruct_bufchan_buf <= is_zae6_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_zaeJ_2_2,MyDTInt_Bool) > (is_zaeJ_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaeJ_2_2_bufchan_d;
  logic is_zaeJ_2_2_bufchan_r;
  assign is_zaeJ_2_2_r = ((! is_zaeJ_2_2_bufchan_d[0]) || is_zaeJ_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_2_2_bufchan_d <= 1'd0;
    else if (is_zaeJ_2_2_r) is_zaeJ_2_2_bufchan_d <= is_zaeJ_2_2_d;
  MyDTInt_Bool_t is_zaeJ_2_2_bufchan_buf;
  assign is_zaeJ_2_2_bufchan_r = (! is_zaeJ_2_2_bufchan_buf[0]);
  assign is_zaeJ_2_2_argbuf_d = (is_zaeJ_2_2_bufchan_buf[0] ? is_zaeJ_2_2_bufchan_buf :
                                 is_zaeJ_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_zaeJ_2_2_argbuf_r && is_zaeJ_2_2_bufchan_buf[0]))
        is_zaeJ_2_2_bufchan_buf <= 1'd0;
      else if (((! is_zaeJ_2_2_argbuf_r) && (! is_zaeJ_2_2_bufchan_buf[0])))
        is_zaeJ_2_2_bufchan_buf <= is_zaeJ_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zaeJ_2_destruct,MyDTInt_Bool) > [(is_zaeJ_2_1,MyDTInt_Bool),
                                                              (is_zaeJ_2_2,MyDTInt_Bool)] */
  logic [1:0] is_zaeJ_2_destruct_emitted;
  logic [1:0] is_zaeJ_2_destruct_done;
  assign is_zaeJ_2_1_d = (is_zaeJ_2_destruct_d[0] && (! is_zaeJ_2_destruct_emitted[0]));
  assign is_zaeJ_2_2_d = (is_zaeJ_2_destruct_d[0] && (! is_zaeJ_2_destruct_emitted[1]));
  assign is_zaeJ_2_destruct_done = (is_zaeJ_2_destruct_emitted | ({is_zaeJ_2_2_d[0],
                                                                   is_zaeJ_2_1_d[0]} & {is_zaeJ_2_2_r,
                                                                                        is_zaeJ_2_1_r}));
  assign is_zaeJ_2_destruct_r = (& is_zaeJ_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_2_destruct_emitted <= 2'd0;
    else
      is_zaeJ_2_destruct_emitted <= (is_zaeJ_2_destruct_r ? 2'd0 :
                                     is_zaeJ_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zaeJ_3_2,MyDTInt_Bool) > (is_zaeJ_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaeJ_3_2_bufchan_d;
  logic is_zaeJ_3_2_bufchan_r;
  assign is_zaeJ_3_2_r = ((! is_zaeJ_3_2_bufchan_d[0]) || is_zaeJ_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_3_2_bufchan_d <= 1'd0;
    else if (is_zaeJ_3_2_r) is_zaeJ_3_2_bufchan_d <= is_zaeJ_3_2_d;
  MyDTInt_Bool_t is_zaeJ_3_2_bufchan_buf;
  assign is_zaeJ_3_2_bufchan_r = (! is_zaeJ_3_2_bufchan_buf[0]);
  assign is_zaeJ_3_2_argbuf_d = (is_zaeJ_3_2_bufchan_buf[0] ? is_zaeJ_3_2_bufchan_buf :
                                 is_zaeJ_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_zaeJ_3_2_argbuf_r && is_zaeJ_3_2_bufchan_buf[0]))
        is_zaeJ_3_2_bufchan_buf <= 1'd0;
      else if (((! is_zaeJ_3_2_argbuf_r) && (! is_zaeJ_3_2_bufchan_buf[0])))
        is_zaeJ_3_2_bufchan_buf <= is_zaeJ_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_zaeJ_3_destruct,MyDTInt_Bool) > [(is_zaeJ_3_1,MyDTInt_Bool),
                                                              (is_zaeJ_3_2,MyDTInt_Bool)] */
  logic [1:0] is_zaeJ_3_destruct_emitted;
  logic [1:0] is_zaeJ_3_destruct_done;
  assign is_zaeJ_3_1_d = (is_zaeJ_3_destruct_d[0] && (! is_zaeJ_3_destruct_emitted[0]));
  assign is_zaeJ_3_2_d = (is_zaeJ_3_destruct_d[0] && (! is_zaeJ_3_destruct_emitted[1]));
  assign is_zaeJ_3_destruct_done = (is_zaeJ_3_destruct_emitted | ({is_zaeJ_3_2_d[0],
                                                                   is_zaeJ_3_1_d[0]} & {is_zaeJ_3_2_r,
                                                                                        is_zaeJ_3_1_r}));
  assign is_zaeJ_3_destruct_r = (& is_zaeJ_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_3_destruct_emitted <= 2'd0;
    else
      is_zaeJ_3_destruct_emitted <= (is_zaeJ_3_destruct_r ? 2'd0 :
                                     is_zaeJ_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_zaeJ_4_destruct,MyDTInt_Bool) > (is_zaeJ_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_zaeJ_4_destruct_bufchan_d;
  logic is_zaeJ_4_destruct_bufchan_r;
  assign is_zaeJ_4_destruct_r = ((! is_zaeJ_4_destruct_bufchan_d[0]) || is_zaeJ_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_zaeJ_4_destruct_r)
        is_zaeJ_4_destruct_bufchan_d <= is_zaeJ_4_destruct_d;
  MyDTInt_Bool_t is_zaeJ_4_destruct_bufchan_buf;
  assign is_zaeJ_4_destruct_bufchan_r = (! is_zaeJ_4_destruct_bufchan_buf[0]);
  assign is_zaeJ_4_1_argbuf_d = (is_zaeJ_4_destruct_bufchan_buf[0] ? is_zaeJ_4_destruct_bufchan_buf :
                                 is_zaeJ_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_zaeJ_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_zaeJ_4_1_argbuf_r && is_zaeJ_4_destruct_bufchan_buf[0]))
        is_zaeJ_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_zaeJ_4_1_argbuf_r) && (! is_zaeJ_4_destruct_bufchan_buf[0])))
        is_zaeJ_4_destruct_bufchan_buf <= is_zaeJ_4_destruct_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet13_1QNode_Int,QTree_Int) > [(q1aeR_destruct,Pointer_QTree_Int),
                                                                  (q2aeS_destruct,Pointer_QTree_Int),
                                                                  (q3aeT_destruct,Pointer_QTree_Int),
                                                                  (q4aeU_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet13_1QNode_Int_emitted;
  logic [3:0] lizzieLet13_1QNode_Int_done;
  assign q1aeR_destruct_d = {lizzieLet13_1QNode_Int_d[18:3],
                             (lizzieLet13_1QNode_Int_d[0] && (! lizzieLet13_1QNode_Int_emitted[0]))};
  assign q2aeS_destruct_d = {lizzieLet13_1QNode_Int_d[34:19],
                             (lizzieLet13_1QNode_Int_d[0] && (! lizzieLet13_1QNode_Int_emitted[1]))};
  assign q3aeT_destruct_d = {lizzieLet13_1QNode_Int_d[50:35],
                             (lizzieLet13_1QNode_Int_d[0] && (! lizzieLet13_1QNode_Int_emitted[2]))};
  assign q4aeU_destruct_d = {lizzieLet13_1QNode_Int_d[66:51],
                             (lizzieLet13_1QNode_Int_d[0] && (! lizzieLet13_1QNode_Int_emitted[3]))};
  assign lizzieLet13_1QNode_Int_done = (lizzieLet13_1QNode_Int_emitted | ({q4aeU_destruct_d[0],
                                                                           q3aeT_destruct_d[0],
                                                                           q2aeS_destruct_d[0],
                                                                           q1aeR_destruct_d[0]} & {q4aeU_destruct_r,
                                                                                                   q3aeT_destruct_r,
                                                                                                   q2aeS_destruct_r,
                                                                                                   q1aeR_destruct_r}));
  assign lizzieLet13_1QNode_Int_r = (& lizzieLet13_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet13_1QNode_Int_emitted <= (lizzieLet13_1QNode_Int_r ? 4'd0 :
                                         lizzieLet13_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet13_1QVal_Int,QTree_Int) > [(v1aeL_destruct,Int)] */
  assign v1aeL_destruct_d = {lizzieLet13_1QVal_Int_d[34:3],
                             lizzieLet13_1QVal_Int_d[0]};
  assign lizzieLet13_1QVal_Int_r = v1aeL_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet13_2,QTree_Int) (lizzieLet13_1,QTree_Int) > [(_162,QTree_Int),
                                                                              (lizzieLet13_1QVal_Int,QTree_Int),
                                                                              (lizzieLet13_1QNode_Int,QTree_Int),
                                                                              (_161,QTree_Int)] */
  logic [3:0] lizzieLet13_1_onehotd;
  always_comb
    if ((lizzieLet13_2_d[0] && lizzieLet13_1_d[0]))
      unique case (lizzieLet13_2_d[2:1])
        2'd0: lizzieLet13_1_onehotd = 4'd1;
        2'd1: lizzieLet13_1_onehotd = 4'd2;
        2'd2: lizzieLet13_1_onehotd = 4'd4;
        2'd3: lizzieLet13_1_onehotd = 4'd8;
        default: lizzieLet13_1_onehotd = 4'd0;
      endcase
    else lizzieLet13_1_onehotd = 4'd0;
  assign _162_d = {lizzieLet13_1_d[66:1], lizzieLet13_1_onehotd[0]};
  assign lizzieLet13_1QVal_Int_d = {lizzieLet13_1_d[66:1],
                                    lizzieLet13_1_onehotd[1]};
  assign lizzieLet13_1QNode_Int_d = {lizzieLet13_1_d[66:1],
                                     lizzieLet13_1_onehotd[2]};
  assign _161_d = {lizzieLet13_1_d[66:1], lizzieLet13_1_onehotd[3]};
  assign lizzieLet13_1_r = (| (lizzieLet13_1_onehotd & {_161_r,
                                                        lizzieLet13_1QNode_Int_r,
                                                        lizzieLet13_1QVal_Int_r,
                                                        _162_r}));
  assign lizzieLet13_2_r = lizzieLet13_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet13_3,QTree_Int) (go_10_goMux_data,Go) > [(lizzieLet13_3QNone_Int,Go),
                                                                   (lizzieLet13_3QVal_Int,Go),
                                                                   (lizzieLet13_3QNode_Int,Go),
                                                                   (lizzieLet13_3QError_Int,Go)] */
  logic [3:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet13_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet13_3_d[2:1])
        2'd0: go_10_goMux_data_onehotd = 4'd1;
        2'd1: go_10_goMux_data_onehotd = 4'd2;
        2'd2: go_10_goMux_data_onehotd = 4'd4;
        2'd3: go_10_goMux_data_onehotd = 4'd8;
        default: go_10_goMux_data_onehotd = 4'd0;
      endcase
    else go_10_goMux_data_onehotd = 4'd0;
  assign lizzieLet13_3QNone_Int_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet13_3QVal_Int_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet13_3QNode_Int_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet13_3QError_Int_d = go_10_goMux_data_onehotd[3];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet13_3QError_Int_r,
                                                              lizzieLet13_3QNode_Int_r,
                                                              lizzieLet13_3QVal_Int_r,
                                                              lizzieLet13_3QNone_Int_r}));
  assign lizzieLet13_3_r = go_10_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet13_3QError_Int,Go) > [(lizzieLet13_3QError_Int_1,Go),
                                               (lizzieLet13_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet13_3QError_Int_emitted;
  logic [1:0] lizzieLet13_3QError_Int_done;
  assign lizzieLet13_3QError_Int_1_d = (lizzieLet13_3QError_Int_d[0] && (! lizzieLet13_3QError_Int_emitted[0]));
  assign lizzieLet13_3QError_Int_2_d = (lizzieLet13_3QError_Int_d[0] && (! lizzieLet13_3QError_Int_emitted[1]));
  assign lizzieLet13_3QError_Int_done = (lizzieLet13_3QError_Int_emitted | ({lizzieLet13_3QError_Int_2_d[0],
                                                                             lizzieLet13_3QError_Int_1_d[0]} & {lizzieLet13_3QError_Int_2_r,
                                                                                                                lizzieLet13_3QError_Int_1_r}));
  assign lizzieLet13_3QError_Int_r = (& lizzieLet13_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet13_3QError_Int_emitted <= (lizzieLet13_3QError_Int_r ? 2'd0 :
                                          lizzieLet13_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_3QError_Int_1,Go)] > (lizzieLet13_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_3QError_Int_1_d[0]}), lizzieLet13_3QError_Int_1_d);
  assign {lizzieLet13_3QError_Int_1_r} = {1 {(lizzieLet13_3QError_Int_1QError_Int_r && lizzieLet13_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet23_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_3QError_Int_1QError_Int_r = ((! lizzieLet13_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet13_3QError_Int_1QError_Int_r)
        lizzieLet13_3QError_Int_1QError_Int_bufchan_d <= lizzieLet13_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet13_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet13_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet13_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet13_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet13_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_3QError_Int_2,Go) > (lizzieLet13_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet13_3QError_Int_2_bufchan_d;
  logic lizzieLet13_3QError_Int_2_bufchan_r;
  assign lizzieLet13_3QError_Int_2_r = ((! lizzieLet13_3QError_Int_2_bufchan_d[0]) || lizzieLet13_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_3QError_Int_2_r)
        lizzieLet13_3QError_Int_2_bufchan_d <= lizzieLet13_3QError_Int_2_d;
  Go_t lizzieLet13_3QError_Int_2_bufchan_buf;
  assign lizzieLet13_3QError_Int_2_bufchan_r = (! lizzieLet13_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet13_3QError_Int_2_argbuf_d = (lizzieLet13_3QError_Int_2_bufchan_buf[0] ? lizzieLet13_3QError_Int_2_bufchan_buf :
                                               lizzieLet13_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_3QError_Int_2_argbuf_r && lizzieLet13_3QError_Int_2_bufchan_buf[0]))
        lizzieLet13_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_3QError_Int_2_argbuf_r) && (! lizzieLet13_3QError_Int_2_bufchan_buf[0])))
        lizzieLet13_3QError_Int_2_bufchan_buf <= lizzieLet13_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_3QNone_Int,Go) > (lizzieLet13_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet13_3QNone_Int_bufchan_d;
  logic lizzieLet13_3QNone_Int_bufchan_r;
  assign lizzieLet13_3QNone_Int_r = ((! lizzieLet13_3QNone_Int_bufchan_d[0]) || lizzieLet13_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_3QNone_Int_r)
        lizzieLet13_3QNone_Int_bufchan_d <= lizzieLet13_3QNone_Int_d;
  Go_t lizzieLet13_3QNone_Int_bufchan_buf;
  assign lizzieLet13_3QNone_Int_bufchan_r = (! lizzieLet13_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_3QNone_Int_1_argbuf_d = (lizzieLet13_3QNone_Int_bufchan_buf[0] ? lizzieLet13_3QNone_Int_bufchan_buf :
                                              lizzieLet13_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_3QNone_Int_1_argbuf_r && lizzieLet13_3QNone_Int_bufchan_buf[0]))
        lizzieLet13_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_3QNone_Int_1_argbuf_r) && (! lizzieLet13_3QNone_Int_bufchan_buf[0])))
        lizzieLet13_3QNone_Int_bufchan_buf <= lizzieLet13_3QNone_Int_bufchan_d;
  
  /* mergectrl (Ty C11,Ty Go) : [(lizzieLet13_3QNone_Int_1_argbuf,Go),
                            (lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf,Go),
                            (lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf,Go),
                            (es_2_1MyFalse_1_argbuf,Go),
                            (es_2_1MyTrue_2_argbuf,Go),
                            (lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf,Go),
                            (lizzieLet13_5QVal_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf,Go),
                            (lizzieLet13_5QNode_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet13_3QError_Int_2_argbuf,Go)] > (go_17_goMux_choice,C11) (go_17_goMux_data,Go) */
  logic [10:0] lizzieLet13_3QNone_Int_1_argbuf_select_d;
  assign lizzieLet13_3QNone_Int_1_argbuf_select_d = ((| lizzieLet13_3QNone_Int_1_argbuf_select_q) ? lizzieLet13_3QNone_Int_1_argbuf_select_q :
                                                     (lizzieLet13_3QNone_Int_1_argbuf_d[0] ? 11'd1 :
                                                      (\lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_d [0] ? 11'd2 :
                                                       (lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_d[0] ? 11'd4 :
                                                        (es_2_1MyFalse_1_argbuf_d[0] ? 11'd8 :
                                                         (es_2_1MyTrue_2_argbuf_d[0] ? 11'd16 :
                                                          (lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_d[0] ? 11'd32 :
                                                           (lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_d[0] ? 11'd64 :
                                                            (lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_d[0] ? 11'd128 :
                                                             (lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_d[0] ? 11'd256 :
                                                              (lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_d[0] ? 11'd512 :
                                                               (lizzieLet13_3QError_Int_2_argbuf_d[0] ? 11'd1024 :
                                                                11'd0))))))))))));
  logic [10:0] lizzieLet13_3QNone_Int_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_3QNone_Int_1_argbuf_select_q <= 11'd0;
    else
      lizzieLet13_3QNone_Int_1_argbuf_select_q <= (lizzieLet13_3QNone_Int_1_argbuf_done ? 11'd0 :
                                                   lizzieLet13_3QNone_Int_1_argbuf_select_d);
  logic [1:0] lizzieLet13_3QNone_Int_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_3QNone_Int_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet13_3QNone_Int_1_argbuf_emit_q <= (lizzieLet13_3QNone_Int_1_argbuf_done ? 2'd0 :
                                                 lizzieLet13_3QNone_Int_1_argbuf_emit_d);
  logic [1:0] lizzieLet13_3QNone_Int_1_argbuf_emit_d;
  assign lizzieLet13_3QNone_Int_1_argbuf_emit_d = (lizzieLet13_3QNone_Int_1_argbuf_emit_q | ({go_17_goMux_choice_d[0],
                                                                                              go_17_goMux_data_d[0]} & {go_17_goMux_choice_r,
                                                                                                                        go_17_goMux_data_r}));
  logic lizzieLet13_3QNone_Int_1_argbuf_done;
  assign lizzieLet13_3QNone_Int_1_argbuf_done = (& lizzieLet13_3QNone_Int_1_argbuf_emit_d);
  assign {lizzieLet13_3QError_Int_2_argbuf_r,
          lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_r,
          es_2_1MyTrue_2_argbuf_r,
          es_2_1MyFalse_1_argbuf_r,
          lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_r,
          \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_r ,
          lizzieLet13_3QNone_Int_1_argbuf_r} = (lizzieLet13_3QNone_Int_1_argbuf_done ? lizzieLet13_3QNone_Int_1_argbuf_select_d :
                                                11'd0);
  assign go_17_goMux_data_d = ((lizzieLet13_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_3QNone_Int_1_argbuf_d :
                               ((lizzieLet13_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_d  :
                                ((lizzieLet13_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_d :
                                 ((lizzieLet13_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? es_2_1MyFalse_1_argbuf_d :
                                  ((lizzieLet13_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? es_2_1MyTrue_2_argbuf_d :
                                   ((lizzieLet13_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_d :
                                    ((lizzieLet13_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_d :
                                     ((lizzieLet13_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_d :
                                      ((lizzieLet13_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_d :
                                       ((lizzieLet13_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_d :
                                        ((lizzieLet13_3QNone_Int_1_argbuf_select_d[10] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet13_3QError_Int_2_argbuf_d :
                                         1'd0)))))))))));
  assign go_17_goMux_choice_d = ((lizzieLet13_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C1_11_dc(1'd1) :
                                 ((lizzieLet13_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C2_11_dc(1'd1) :
                                  ((lizzieLet13_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C3_11_dc(1'd1) :
                                   ((lizzieLet13_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C4_11_dc(1'd1) :
                                    ((lizzieLet13_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C5_11_dc(1'd1) :
                                     ((lizzieLet13_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C6_11_dc(1'd1) :
                                      ((lizzieLet13_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C7_11_dc(1'd1) :
                                       ((lizzieLet13_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C8_11_dc(1'd1) :
                                        ((lizzieLet13_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C9_11_dc(1'd1) :
                                         ((lizzieLet13_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C10_11_dc(1'd1) :
                                          ((lizzieLet13_3QNone_Int_1_argbuf_select_d[10] && (! lizzieLet13_3QNone_Int_1_argbuf_emit_q[1])) ? C11_11_dc(1'd1) :
                                           {4'd0, 1'd0})))))))))));
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet13_4,QTree_Int) (is_zaeJ_goMux_mux,MyDTInt_Bool) > [(_160,MyDTInt_Bool),
                                                                                        (lizzieLet13_4QVal_Int,MyDTInt_Bool),
                                                                                        (lizzieLet13_4QNode_Int,MyDTInt_Bool),
                                                                                        (_159,MyDTInt_Bool)] */
  logic [3:0] is_zaeJ_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_4_d[0] && is_zaeJ_goMux_mux_d[0]))
      unique case (lizzieLet13_4_d[2:1])
        2'd0: is_zaeJ_goMux_mux_onehotd = 4'd1;
        2'd1: is_zaeJ_goMux_mux_onehotd = 4'd2;
        2'd2: is_zaeJ_goMux_mux_onehotd = 4'd4;
        2'd3: is_zaeJ_goMux_mux_onehotd = 4'd8;
        default: is_zaeJ_goMux_mux_onehotd = 4'd0;
      endcase
    else is_zaeJ_goMux_mux_onehotd = 4'd0;
  assign _160_d = is_zaeJ_goMux_mux_onehotd[0];
  assign lizzieLet13_4QVal_Int_d = is_zaeJ_goMux_mux_onehotd[1];
  assign lizzieLet13_4QNode_Int_d = is_zaeJ_goMux_mux_onehotd[2];
  assign _159_d = is_zaeJ_goMux_mux_onehotd[3];
  assign is_zaeJ_goMux_mux_r = (| (is_zaeJ_goMux_mux_onehotd & {_159_r,
                                                                lizzieLet13_4QNode_Int_r,
                                                                lizzieLet13_4QVal_Int_r,
                                                                _160_r}));
  assign lizzieLet13_4_r = is_zaeJ_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet13_5,QTree_Int) (readPointer_QTree_Intm3aeI_1_argbuf_rwb,QTree_Int) > [(_158,QTree_Int),
                                                                                                        (lizzieLet13_5QVal_Int,QTree_Int),
                                                                                                        (lizzieLet13_5QNode_Int,QTree_Int),
                                                                                                        (_157,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet13_5_d[0] && readPointer_QTree_Intm3aeI_1_argbuf_rwb_d[0]))
      unique case (lizzieLet13_5_d[2:1])
        2'd0: readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd = 4'd0;
  assign _158_d = {readPointer_QTree_Intm3aeI_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet13_5QVal_Int_d = {readPointer_QTree_Intm3aeI_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet13_5QNode_Int_d = {readPointer_QTree_Intm3aeI_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd[2]};
  assign _157_d = {readPointer_QTree_Intm3aeI_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intm3aeI_1_argbuf_rwb_r = (| (readPointer_QTree_Intm3aeI_1_argbuf_rwb_onehotd & {_157_r,
                                                                                                            lizzieLet13_5QNode_Int_r,
                                                                                                            lizzieLet13_5QVal_Int_r,
                                                                                                            _158_r}));
  assign lizzieLet13_5_r = readPointer_QTree_Intm3aeI_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet13_5QNode_Int,QTree_Int) > [(lizzieLet13_5QNode_Int_1,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_2,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_3,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_4,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_5,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_6,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_7,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_8,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_9,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_10,QTree_Int),
                                                            (lizzieLet13_5QNode_Int_11,QTree_Int)] */
  logic [10:0] lizzieLet13_5QNode_Int_emitted;
  logic [10:0] lizzieLet13_5QNode_Int_done;
  assign lizzieLet13_5QNode_Int_1_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[0]))};
  assign lizzieLet13_5QNode_Int_2_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[1]))};
  assign lizzieLet13_5QNode_Int_3_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[2]))};
  assign lizzieLet13_5QNode_Int_4_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[3]))};
  assign lizzieLet13_5QNode_Int_5_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[4]))};
  assign lizzieLet13_5QNode_Int_6_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[5]))};
  assign lizzieLet13_5QNode_Int_7_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[6]))};
  assign lizzieLet13_5QNode_Int_8_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[7]))};
  assign lizzieLet13_5QNode_Int_9_d = {lizzieLet13_5QNode_Int_d[66:1],
                                       (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[8]))};
  assign lizzieLet13_5QNode_Int_10_d = {lizzieLet13_5QNode_Int_d[66:1],
                                        (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[9]))};
  assign lizzieLet13_5QNode_Int_11_d = {lizzieLet13_5QNode_Int_d[66:1],
                                        (lizzieLet13_5QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_emitted[10]))};
  assign lizzieLet13_5QNode_Int_done = (lizzieLet13_5QNode_Int_emitted | ({lizzieLet13_5QNode_Int_11_d[0],
                                                                           lizzieLet13_5QNode_Int_10_d[0],
                                                                           lizzieLet13_5QNode_Int_9_d[0],
                                                                           lizzieLet13_5QNode_Int_8_d[0],
                                                                           lizzieLet13_5QNode_Int_7_d[0],
                                                                           lizzieLet13_5QNode_Int_6_d[0],
                                                                           lizzieLet13_5QNode_Int_5_d[0],
                                                                           lizzieLet13_5QNode_Int_4_d[0],
                                                                           lizzieLet13_5QNode_Int_3_d[0],
                                                                           lizzieLet13_5QNode_Int_2_d[0],
                                                                           lizzieLet13_5QNode_Int_1_d[0]} & {lizzieLet13_5QNode_Int_11_r,
                                                                                                             lizzieLet13_5QNode_Int_10_r,
                                                                                                             lizzieLet13_5QNode_Int_9_r,
                                                                                                             lizzieLet13_5QNode_Int_8_r,
                                                                                                             lizzieLet13_5QNode_Int_7_r,
                                                                                                             lizzieLet13_5QNode_Int_6_r,
                                                                                                             lizzieLet13_5QNode_Int_5_r,
                                                                                                             lizzieLet13_5QNode_Int_4_r,
                                                                                                             lizzieLet13_5QNode_Int_3_r,
                                                                                                             lizzieLet13_5QNode_Int_2_r,
                                                                                                             lizzieLet13_5QNode_Int_1_r}));
  assign lizzieLet13_5QNode_Int_r = (& lizzieLet13_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_5QNode_Int_emitted <= 11'd0;
    else
      lizzieLet13_5QNode_Int_emitted <= (lizzieLet13_5QNode_Int_r ? 11'd0 :
                                         lizzieLet13_5QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_10,QTree_Int) (q3aeT_destruct,Pointer_QTree_Int) > [(_156,Pointer_QTree_Int),
                                                                                                           (_155,Pointer_QTree_Int),
                                                                                                           (lizzieLet13_5QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                           (_154,Pointer_QTree_Int)] */
  logic [3:0] q3aeT_destruct_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_10_d[0] && q3aeT_destruct_d[0]))
      unique case (lizzieLet13_5QNode_Int_10_d[2:1])
        2'd0: q3aeT_destruct_onehotd = 4'd1;
        2'd1: q3aeT_destruct_onehotd = 4'd2;
        2'd2: q3aeT_destruct_onehotd = 4'd4;
        2'd3: q3aeT_destruct_onehotd = 4'd8;
        default: q3aeT_destruct_onehotd = 4'd0;
      endcase
    else q3aeT_destruct_onehotd = 4'd0;
  assign _156_d = {q3aeT_destruct_d[16:1],
                   q3aeT_destruct_onehotd[0]};
  assign _155_d = {q3aeT_destruct_d[16:1],
                   q3aeT_destruct_onehotd[1]};
  assign lizzieLet13_5QNode_Int_10QNode_Int_d = {q3aeT_destruct_d[16:1],
                                                 q3aeT_destruct_onehotd[2]};
  assign _154_d = {q3aeT_destruct_d[16:1],
                   q3aeT_destruct_onehotd[3]};
  assign q3aeT_destruct_r = (| (q3aeT_destruct_onehotd & {_154_r,
                                                          lizzieLet13_5QNode_Int_10QNode_Int_r,
                                                          _155_r,
                                                          _156_r}));
  assign lizzieLet13_5QNode_Int_10_r = q3aeT_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_11,QTree_Int) (q4aeU_destruct,Pointer_QTree_Int) > [(_153,Pointer_QTree_Int),
                                                                                                           (_152,Pointer_QTree_Int),
                                                                                                           (lizzieLet13_5QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                           (_151,Pointer_QTree_Int)] */
  logic [3:0] q4aeU_destruct_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_11_d[0] && q4aeU_destruct_d[0]))
      unique case (lizzieLet13_5QNode_Int_11_d[2:1])
        2'd0: q4aeU_destruct_onehotd = 4'd1;
        2'd1: q4aeU_destruct_onehotd = 4'd2;
        2'd2: q4aeU_destruct_onehotd = 4'd4;
        2'd3: q4aeU_destruct_onehotd = 4'd8;
        default: q4aeU_destruct_onehotd = 4'd0;
      endcase
    else q4aeU_destruct_onehotd = 4'd0;
  assign _153_d = {q4aeU_destruct_d[16:1],
                   q4aeU_destruct_onehotd[0]};
  assign _152_d = {q4aeU_destruct_d[16:1],
                   q4aeU_destruct_onehotd[1]};
  assign lizzieLet13_5QNode_Int_11QNode_Int_d = {q4aeU_destruct_d[16:1],
                                                 q4aeU_destruct_onehotd[2]};
  assign _151_d = {q4aeU_destruct_d[16:1],
                   q4aeU_destruct_onehotd[3]};
  assign q4aeU_destruct_r = (| (q4aeU_destruct_onehotd & {_151_r,
                                                          lizzieLet13_5QNode_Int_11QNode_Int_r,
                                                          _152_r,
                                                          _153_r}));
  assign lizzieLet13_5QNode_Int_11_r = q4aeU_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_11QNode_Int,Pointer_QTree_Int) > (lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_11QNode_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_11QNode_Int_r = ((! lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_11QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QNode_Int_11QNode_Int_r)
        lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d <= lizzieLet13_5QNode_Int_11QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_11QNode_Int_bufchan_r = (! lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf :
                                                          lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_r && lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QNode_Int_11QNode_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_11QNode_Int_bufchan_buf <= lizzieLet13_5QNode_Int_11QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet13_5QNode_Int_1QNode_Int,QTree_Int) > [(t1aeW_destruct,Pointer_QTree_Int),
                                                                             (t2aeX_destruct,Pointer_QTree_Int),
                                                                             (t3aeY_destruct,Pointer_QTree_Int),
                                                                             (t4aeZ_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet13_5QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet13_5QNode_Int_1QNode_Int_done;
  assign t1aeW_destruct_d = {lizzieLet13_5QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet13_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_1QNode_Int_emitted[0]))};
  assign t2aeX_destruct_d = {lizzieLet13_5QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet13_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_1QNode_Int_emitted[1]))};
  assign t3aeY_destruct_d = {lizzieLet13_5QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet13_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_1QNode_Int_emitted[2]))};
  assign t4aeZ_destruct_d = {lizzieLet13_5QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet13_5QNode_Int_1QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet13_5QNode_Int_1QNode_Int_done = (lizzieLet13_5QNode_Int_1QNode_Int_emitted | ({t4aeZ_destruct_d[0],
                                                                                                 t3aeY_destruct_d[0],
                                                                                                 t2aeX_destruct_d[0],
                                                                                                 t1aeW_destruct_d[0]} & {t4aeZ_destruct_r,
                                                                                                                         t3aeY_destruct_r,
                                                                                                                         t2aeX_destruct_r,
                                                                                                                         t1aeW_destruct_r}));
  assign lizzieLet13_5QNode_Int_1QNode_Int_r = (& lizzieLet13_5QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet13_5QNode_Int_1QNode_Int_emitted <= (lizzieLet13_5QNode_Int_1QNode_Int_r ? 4'd0 :
                                                    lizzieLet13_5QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet13_5QNode_Int_2,QTree_Int) (lizzieLet13_5QNode_Int_1,QTree_Int) > [(_150,QTree_Int),
                                                                                                    (_149,QTree_Int),
                                                                                                    (lizzieLet13_5QNode_Int_1QNode_Int,QTree_Int),
                                                                                                    (_148,QTree_Int)] */
  logic [3:0] lizzieLet13_5QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_2_d[0] && lizzieLet13_5QNode_Int_1_d[0]))
      unique case (lizzieLet13_5QNode_Int_2_d[2:1])
        2'd0: lizzieLet13_5QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet13_5QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet13_5QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet13_5QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet13_5QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet13_5QNode_Int_1_onehotd = 4'd0;
  assign _150_d = {lizzieLet13_5QNode_Int_1_d[66:1],
                   lizzieLet13_5QNode_Int_1_onehotd[0]};
  assign _149_d = {lizzieLet13_5QNode_Int_1_d[66:1],
                   lizzieLet13_5QNode_Int_1_onehotd[1]};
  assign lizzieLet13_5QNode_Int_1QNode_Int_d = {lizzieLet13_5QNode_Int_1_d[66:1],
                                                lizzieLet13_5QNode_Int_1_onehotd[2]};
  assign _148_d = {lizzieLet13_5QNode_Int_1_d[66:1],
                   lizzieLet13_5QNode_Int_1_onehotd[3]};
  assign lizzieLet13_5QNode_Int_1_r = (| (lizzieLet13_5QNode_Int_1_onehotd & {_148_r,
                                                                              lizzieLet13_5QNode_Int_1QNode_Int_r,
                                                                              _149_r,
                                                                              _150_r}));
  assign lizzieLet13_5QNode_Int_2_r = lizzieLet13_5QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet13_5QNode_Int_3,QTree_Int) (lizzieLet13_3QNode_Int,Go) > [(lizzieLet13_5QNode_Int_3QNone_Int,Go),
                                                                                    (lizzieLet13_5QNode_Int_3QVal_Int,Go),
                                                                                    (lizzieLet13_5QNode_Int_3QNode_Int,Go),
                                                                                    (lizzieLet13_5QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet13_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_3_d[0] && lizzieLet13_3QNode_Int_d[0]))
      unique case (lizzieLet13_5QNode_Int_3_d[2:1])
        2'd0: lizzieLet13_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet13_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet13_5QNode_Int_3QNone_Int_d = lizzieLet13_3QNode_Int_onehotd[0];
  assign lizzieLet13_5QNode_Int_3QVal_Int_d = lizzieLet13_3QNode_Int_onehotd[1];
  assign lizzieLet13_5QNode_Int_3QNode_Int_d = lizzieLet13_3QNode_Int_onehotd[2];
  assign lizzieLet13_5QNode_Int_3QError_Int_d = lizzieLet13_3QNode_Int_onehotd[3];
  assign lizzieLet13_3QNode_Int_r = (| (lizzieLet13_3QNode_Int_onehotd & {lizzieLet13_5QNode_Int_3QError_Int_r,
                                                                          lizzieLet13_5QNode_Int_3QNode_Int_r,
                                                                          lizzieLet13_5QNode_Int_3QVal_Int_r,
                                                                          lizzieLet13_5QNode_Int_3QNone_Int_r}));
  assign lizzieLet13_5QNode_Int_3_r = lizzieLet13_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet13_5QNode_Int_3QError_Int,Go) > [(lizzieLet13_5QNode_Int_3QError_Int_1,Go),
                                                          (lizzieLet13_5QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet13_5QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet13_5QNode_Int_3QError_Int_done;
  assign lizzieLet13_5QNode_Int_3QError_Int_1_d = (lizzieLet13_5QNode_Int_3QError_Int_d[0] && (! lizzieLet13_5QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet13_5QNode_Int_3QError_Int_2_d = (lizzieLet13_5QNode_Int_3QError_Int_d[0] && (! lizzieLet13_5QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet13_5QNode_Int_3QError_Int_done = (lizzieLet13_5QNode_Int_3QError_Int_emitted | ({lizzieLet13_5QNode_Int_3QError_Int_2_d[0],
                                                                                                   lizzieLet13_5QNode_Int_3QError_Int_1_d[0]} & {lizzieLet13_5QNode_Int_3QError_Int_2_r,
                                                                                                                                                 lizzieLet13_5QNode_Int_3QError_Int_1_r}));
  assign lizzieLet13_5QNode_Int_3QError_Int_r = (& lizzieLet13_5QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QNode_Int_3QError_Int_emitted <= (lizzieLet13_5QNode_Int_3QError_Int_r ? 2'd0 :
                                                     lizzieLet13_5QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_5QNode_Int_3QError_Int_1,Go)] > (lizzieLet13_5QNode_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_5QNode_Int_3QError_Int_1_d[0]}), lizzieLet13_5QNode_Int_3QError_Int_1_d);
  assign {lizzieLet13_5QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_r && lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_5QNode_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet22_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_r = ((! lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_r)
        lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet13_5QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QNode_Int_3QError_Int_2,Go) > (lizzieLet13_5QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QError_Int_2_r = ((! lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_3QError_Int_2_r)
        lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet13_5QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf :
                                                          lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_r && lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet13_5QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QNode_Int_3QNode_Int,Go) > (lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QNode_Int_r = ((! lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_3QNode_Int_r)
        lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d <= lizzieLet13_5QNode_Int_3QNode_Int_d;
  Go_t lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet13_5QNode_Int_3QNode_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QNode_Int_3QNone_Int,Go) > (lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QNone_Int_r = ((! lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_3QNone_Int_r)
        lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d <= lizzieLet13_5QNode_Int_3QNone_Int_d;
  Go_t lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet13_5QNode_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet13_5QNode_Int_3QVal_Int,Go) > [(lizzieLet13_5QNode_Int_3QVal_Int_1,Go),
                                                        (lizzieLet13_5QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet13_5QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet13_5QNode_Int_3QVal_Int_done;
  assign lizzieLet13_5QNode_Int_3QVal_Int_1_d = (lizzieLet13_5QNode_Int_3QVal_Int_d[0] && (! lizzieLet13_5QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet13_5QNode_Int_3QVal_Int_2_d = (lizzieLet13_5QNode_Int_3QVal_Int_d[0] && (! lizzieLet13_5QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet13_5QNode_Int_3QVal_Int_done = (lizzieLet13_5QNode_Int_3QVal_Int_emitted | ({lizzieLet13_5QNode_Int_3QVal_Int_2_d[0],
                                                                                               lizzieLet13_5QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet13_5QNode_Int_3QVal_Int_2_r,
                                                                                                                                           lizzieLet13_5QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet13_5QNode_Int_3QVal_Int_r = (& lizzieLet13_5QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QNode_Int_3QVal_Int_emitted <= (lizzieLet13_5QNode_Int_3QVal_Int_r ? 2'd0 :
                                                   lizzieLet13_5QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_5QNode_Int_3QVal_Int_1,Go)] > (lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_5QNode_Int_3QVal_Int_1_d[0]}), lizzieLet13_5QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet13_5QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_r && lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet20_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_r = ((! lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_r)
        lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet13_5QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QNode_Int_3QVal_Int_2,Go) > (lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet13_5QNode_Int_3QVal_Int_2_r = ((! lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_3QVal_Int_2_r)
        lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet13_5QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf :
                                                        lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet13_5QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet13_5QNode_Int_4,QTree_Int) (lizzieLet13_4QNode_Int,MyDTInt_Bool) > [(_147,MyDTInt_Bool),
                                                                                                        (_146,MyDTInt_Bool),
                                                                                                        (lizzieLet13_5QNode_Int_4QNode_Int,MyDTInt_Bool),
                                                                                                        (_145,MyDTInt_Bool)] */
  logic [3:0] lizzieLet13_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_4_d[0] && lizzieLet13_4QNode_Int_d[0]))
      unique case (lizzieLet13_5QNode_Int_4_d[2:1])
        2'd0: lizzieLet13_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet13_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_4QNode_Int_onehotd = 4'd0;
  assign _147_d = lizzieLet13_4QNode_Int_onehotd[0];
  assign _146_d = lizzieLet13_4QNode_Int_onehotd[1];
  assign lizzieLet13_5QNode_Int_4QNode_Int_d = lizzieLet13_4QNode_Int_onehotd[2];
  assign _145_d = lizzieLet13_4QNode_Int_onehotd[3];
  assign lizzieLet13_4QNode_Int_r = (| (lizzieLet13_4QNode_Int_onehotd & {_145_r,
                                                                          lizzieLet13_5QNode_Int_4QNode_Int_r,
                                                                          _146_r,
                                                                          _147_r}));
  assign lizzieLet13_5QNode_Int_4_r = lizzieLet13_4QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet13_5QNode_Int_4QNode_Int,MyDTInt_Bool) > [(lizzieLet13_5QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                                                             (lizzieLet13_5QNode_Int_4QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet13_5QNode_Int_4QNode_Int_emitted;
  logic [1:0] lizzieLet13_5QNode_Int_4QNode_Int_done;
  assign lizzieLet13_5QNode_Int_4QNode_Int_1_d = (lizzieLet13_5QNode_Int_4QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_4QNode_Int_emitted[0]));
  assign lizzieLet13_5QNode_Int_4QNode_Int_2_d = (lizzieLet13_5QNode_Int_4QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_4QNode_Int_emitted[1]));
  assign lizzieLet13_5QNode_Int_4QNode_Int_done = (lizzieLet13_5QNode_Int_4QNode_Int_emitted | ({lizzieLet13_5QNode_Int_4QNode_Int_2_d[0],
                                                                                                 lizzieLet13_5QNode_Int_4QNode_Int_1_d[0]} & {lizzieLet13_5QNode_Int_4QNode_Int_2_r,
                                                                                                                                              lizzieLet13_5QNode_Int_4QNode_Int_1_r}));
  assign lizzieLet13_5QNode_Int_4QNode_Int_r = (& lizzieLet13_5QNode_Int_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_4QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QNode_Int_4QNode_Int_emitted <= (lizzieLet13_5QNode_Int_4QNode_Int_r ? 2'd0 :
                                                    lizzieLet13_5QNode_Int_4QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_5QNode_Int_4QNode_Int_2,MyDTInt_Bool) > (lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d;
  logic lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_r;
  assign lizzieLet13_5QNode_Int_4QNode_Int_2_r = ((! lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d[0]) || lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_4QNode_Int_2_r)
        lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d <= lizzieLet13_5QNode_Int_4QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf;
  assign lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_r = (! lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_d = (lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf[0] ? lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_r && lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_4QNode_Int_2_argbuf_r) && (! lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_buf <= lizzieLet13_5QNode_Int_4QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_5,QTree_Int) (lizzieLet13_6QNode_Int,Pointer_QTree_Int) > [(lizzieLet13_5QNode_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                                  (_144,Pointer_QTree_Int),
                                                                                                                  (_143,Pointer_QTree_Int),
                                                                                                                  (_142,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet13_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_5_d[0] && lizzieLet13_6QNode_Int_d[0]))
      unique case (lizzieLet13_5QNode_Int_5_d[2:1])
        2'd0: lizzieLet13_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet13_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_6QNode_Int_onehotd = 4'd0;
  assign lizzieLet13_5QNode_Int_5QNone_Int_d = {lizzieLet13_6QNode_Int_d[16:1],
                                                lizzieLet13_6QNode_Int_onehotd[0]};
  assign _144_d = {lizzieLet13_6QNode_Int_d[16:1],
                   lizzieLet13_6QNode_Int_onehotd[1]};
  assign _143_d = {lizzieLet13_6QNode_Int_d[16:1],
                   lizzieLet13_6QNode_Int_onehotd[2]};
  assign _142_d = {lizzieLet13_6QNode_Int_d[16:1],
                   lizzieLet13_6QNode_Int_onehotd[3]};
  assign lizzieLet13_6QNode_Int_r = (| (lizzieLet13_6QNode_Int_onehotd & {_142_r,
                                                                          _143_r,
                                                                          _144_r,
                                                                          lizzieLet13_5QNode_Int_5QNone_Int_r}));
  assign lizzieLet13_5QNode_Int_5_r = lizzieLet13_6QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_5QNone_Int_r = ((! lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QNode_Int_5QNone_Int_r)
        lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d <= lizzieLet13_5QNode_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet13_5QNode_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet13_5QNode_Int_6,QTree_Int) (lizzieLet13_8QNode_Int,MyDTInt_Int_Int) > [(_141,MyDTInt_Int_Int),
                                                                                                              (_140,MyDTInt_Int_Int),
                                                                                                              (lizzieLet13_5QNode_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                              (_139,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet13_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_6_d[0] && lizzieLet13_8QNode_Int_d[0]))
      unique case (lizzieLet13_5QNode_Int_6_d[2:1])
        2'd0: lizzieLet13_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet13_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_8QNode_Int_onehotd = 4'd0;
  assign _141_d = lizzieLet13_8QNode_Int_onehotd[0];
  assign _140_d = lizzieLet13_8QNode_Int_onehotd[1];
  assign lizzieLet13_5QNode_Int_6QNode_Int_d = lizzieLet13_8QNode_Int_onehotd[2];
  assign _139_d = lizzieLet13_8QNode_Int_onehotd[3];
  assign lizzieLet13_8QNode_Int_r = (| (lizzieLet13_8QNode_Int_onehotd & {_139_r,
                                                                          lizzieLet13_5QNode_Int_6QNode_Int_r,
                                                                          _140_r,
                                                                          _141_r}));
  assign lizzieLet13_5QNode_Int_6_r = lizzieLet13_8QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet13_5QNode_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet13_5QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                   (lizzieLet13_5QNode_Int_6QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet13_5QNode_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet13_5QNode_Int_6QNode_Int_done;
  assign lizzieLet13_5QNode_Int_6QNode_Int_1_d = (lizzieLet13_5QNode_Int_6QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet13_5QNode_Int_6QNode_Int_2_d = (lizzieLet13_5QNode_Int_6QNode_Int_d[0] && (! lizzieLet13_5QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet13_5QNode_Int_6QNode_Int_done = (lizzieLet13_5QNode_Int_6QNode_Int_emitted | ({lizzieLet13_5QNode_Int_6QNode_Int_2_d[0],
                                                                                                 lizzieLet13_5QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet13_5QNode_Int_6QNode_Int_2_r,
                                                                                                                                              lizzieLet13_5QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet13_5QNode_Int_6QNode_Int_r = (& lizzieLet13_5QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QNode_Int_6QNode_Int_emitted <= (lizzieLet13_5QNode_Int_6QNode_Int_r ? 2'd0 :
                                                    lizzieLet13_5QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet13_5QNode_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet13_5QNode_Int_6QNode_Int_2_r = ((! lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QNode_Int_6QNode_Int_2_r)
        lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet13_5QNode_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet13_5QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QNode_Int_7,QTree_Int) (lizzieLet13_9QNode_Int,Pointer_CTf'_f'_Int) > [(lizzieLet13_5QNode_Int_7QNone_Int,Pointer_CTf'_f'_Int),
                                                                                                                      (lizzieLet13_5QNode_Int_7QVal_Int,Pointer_CTf'_f'_Int),
                                                                                                                      (lizzieLet13_5QNode_Int_7QNode_Int,Pointer_CTf'_f'_Int),
                                                                                                                      (lizzieLet13_5QNode_Int_7QError_Int,Pointer_CTf'_f'_Int)] */
  logic [3:0] lizzieLet13_9QNode_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_7_d[0] && lizzieLet13_9QNode_Int_d[0]))
      unique case (lizzieLet13_5QNode_Int_7_d[2:1])
        2'd0: lizzieLet13_9QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_9QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_9QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_9QNode_Int_onehotd = 4'd8;
        default: lizzieLet13_9QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_9QNode_Int_onehotd = 4'd0;
  assign lizzieLet13_5QNode_Int_7QNone_Int_d = {lizzieLet13_9QNode_Int_d[16:1],
                                                lizzieLet13_9QNode_Int_onehotd[0]};
  assign lizzieLet13_5QNode_Int_7QVal_Int_d = {lizzieLet13_9QNode_Int_d[16:1],
                                               lizzieLet13_9QNode_Int_onehotd[1]};
  assign lizzieLet13_5QNode_Int_7QNode_Int_d = {lizzieLet13_9QNode_Int_d[16:1],
                                                lizzieLet13_9QNode_Int_onehotd[2]};
  assign lizzieLet13_5QNode_Int_7QError_Int_d = {lizzieLet13_9QNode_Int_d[16:1],
                                                 lizzieLet13_9QNode_Int_onehotd[3]};
  assign lizzieLet13_9QNode_Int_r = (| (lizzieLet13_9QNode_Int_onehotd & {lizzieLet13_5QNode_Int_7QError_Int_r,
                                                                          lizzieLet13_5QNode_Int_7QNode_Int_r,
                                                                          lizzieLet13_5QNode_Int_7QVal_Int_r,
                                                                          lizzieLet13_5QNode_Int_7QNone_Int_r}));
  assign lizzieLet13_5QNode_Int_7_r = lizzieLet13_9QNode_Int_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QNode_Int_7QError_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QNode_Int_7QError_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QError_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_7QError_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_7QError_Int_r = ((! lizzieLet13_5QNode_Int_7QError_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QNode_Int_7QError_Int_r)
        lizzieLet13_5QNode_Int_7QError_Int_bufchan_d <= lizzieLet13_5QNode_Int_7QError_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_7QError_Int_bufchan_r = (! lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf :
                                                          lizzieLet13_5QNode_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_r && lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QNode_Int_7QError_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_7QError_Int_bufchan_buf <= lizzieLet13_5QNode_Int_7QError_Int_bufchan_d;
  
  /* dcon (Ty CTf'_f'_Int,
      Dcon Lcall_f'_f'_Int3) : [(lizzieLet13_5QNode_Int_7QNode_Int,Pointer_CTf'_f'_Int),
                                (lizzieLet13_5QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                (t1aeW_destruct,Pointer_QTree_Int),
                                (lizzieLet13_5QNode_Int_4QNode_Int_1,MyDTInt_Bool),
                                (lizzieLet13_5QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                (lizzieLet13_5QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                (t2aeX_destruct,Pointer_QTree_Int),
                                (lizzieLet13_5QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                (t3aeY_destruct,Pointer_QTree_Int)] > (lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3,CTf'_f'_Int) */
  assign \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_d  = \Lcall_f'_f'_Int3_dc ((& {lizzieLet13_5QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                  lizzieLet13_5QNode_Int_8QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                  t1aeW_destruct_d[0],
                                                                                                                                                                                                                                                                                                  lizzieLet13_5QNode_Int_4QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                  lizzieLet13_5QNode_Int_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                  lizzieLet13_5QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                  t2aeX_destruct_d[0],
                                                                                                                                                                                                                                                                                                  lizzieLet13_5QNode_Int_10QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                  t3aeY_destruct_d[0]}), lizzieLet13_5QNode_Int_7QNode_Int_d, lizzieLet13_5QNode_Int_8QNode_Int_d, t1aeW_destruct_d, lizzieLet13_5QNode_Int_4QNode_Int_1_d, lizzieLet13_5QNode_Int_6QNode_Int_1_d, lizzieLet13_5QNode_Int_9QNode_Int_d, t2aeX_destruct_d, lizzieLet13_5QNode_Int_10QNode_Int_d, t3aeY_destruct_d);
  assign {lizzieLet13_5QNode_Int_7QNode_Int_r,
          lizzieLet13_5QNode_Int_8QNode_Int_r,
          t1aeW_destruct_r,
          lizzieLet13_5QNode_Int_4QNode_Int_1_r,
          lizzieLet13_5QNode_Int_6QNode_Int_1_r,
          lizzieLet13_5QNode_Int_9QNode_Int_r,
          t2aeX_destruct_r,
          lizzieLet13_5QNode_Int_10QNode_Int_r,
          t3aeY_destruct_r} = {9 {(\lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_r  && \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_d [0])}};
  
  /* buf (Ty CTf'_f'_Int) : (lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3,CTf'_f'_Int) > (lizzieLet21_1_argbuf,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d ;
  logic \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_r ;
  assign \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_r  = ((! \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d [0]) || \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                                                                                               1'd0};
    else
      if (\lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_r )
        \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d  <= \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_d ;
  \CTf'_f'_Int_t  \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf ;
  assign \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_r  = (! \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf [0]);
  assign lizzieLet21_1_argbuf_d = (\lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf [0] ? \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf  :
                                   \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf [0]))
        \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                                                                                                   1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf [0])))
        \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_buf  <= \lizzieLet13_5QNode_Int_7QNode_Int_1lizzieLet13_5QNode_Int_8QNode_Int_1t1aeW_1lizzieLet13_5QNode_Int_4QNode_Int_1lizzieLet13_5QNode_Int_6QNode_Int_1lizzieLet13_5QNode_Int_9QNode_Int_1t2aeX_1lizzieLet13_5QNode_Int_10QNode_Int_1t3aeY_1Lcall_f'_f'_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QNode_Int_7QNone_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_7QNone_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_7QNone_Int_r = ((! lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QNode_Int_7QNone_Int_r)
        lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d <= lizzieLet13_5QNode_Int_7QNone_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_7QNone_Int_bufchan_r = (! lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf :
                                                         lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_r && lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QNode_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_7QNone_Int_bufchan_buf <= lizzieLet13_5QNode_Int_7QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QNode_Int_7QVal_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d;
  logic lizzieLet13_5QNode_Int_7QVal_Int_bufchan_r;
  assign lizzieLet13_5QNode_Int_7QVal_Int_r = ((! lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d[0]) || lizzieLet13_5QNode_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QNode_Int_7QVal_Int_r)
        lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d <= lizzieLet13_5QNode_Int_7QVal_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet13_5QNode_Int_7QVal_Int_bufchan_r = (! lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_d = (lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf :
                                                        lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_r && lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QNode_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet13_5QNode_Int_7QVal_Int_bufchan_buf <= lizzieLet13_5QNode_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_8,QTree_Int) (q1aeR_destruct,Pointer_QTree_Int) > [(_138,Pointer_QTree_Int),
                                                                                                          (_137,Pointer_QTree_Int),
                                                                                                          (lizzieLet13_5QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                          (_136,Pointer_QTree_Int)] */
  logic [3:0] q1aeR_destruct_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_8_d[0] && q1aeR_destruct_d[0]))
      unique case (lizzieLet13_5QNode_Int_8_d[2:1])
        2'd0: q1aeR_destruct_onehotd = 4'd1;
        2'd1: q1aeR_destruct_onehotd = 4'd2;
        2'd2: q1aeR_destruct_onehotd = 4'd4;
        2'd3: q1aeR_destruct_onehotd = 4'd8;
        default: q1aeR_destruct_onehotd = 4'd0;
      endcase
    else q1aeR_destruct_onehotd = 4'd0;
  assign _138_d = {q1aeR_destruct_d[16:1],
                   q1aeR_destruct_onehotd[0]};
  assign _137_d = {q1aeR_destruct_d[16:1],
                   q1aeR_destruct_onehotd[1]};
  assign lizzieLet13_5QNode_Int_8QNode_Int_d = {q1aeR_destruct_d[16:1],
                                                q1aeR_destruct_onehotd[2]};
  assign _136_d = {q1aeR_destruct_d[16:1],
                   q1aeR_destruct_onehotd[3]};
  assign q1aeR_destruct_r = (| (q1aeR_destruct_onehotd & {_136_r,
                                                          lizzieLet13_5QNode_Int_8QNode_Int_r,
                                                          _137_r,
                                                          _138_r}));
  assign lizzieLet13_5QNode_Int_8_r = q1aeR_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QNode_Int_9,QTree_Int) (q2aeS_destruct,Pointer_QTree_Int) > [(_135,Pointer_QTree_Int),
                                                                                                          (_134,Pointer_QTree_Int),
                                                                                                          (lizzieLet13_5QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                          (_133,Pointer_QTree_Int)] */
  logic [3:0] q2aeS_destruct_onehotd;
  always_comb
    if ((lizzieLet13_5QNode_Int_9_d[0] && q2aeS_destruct_d[0]))
      unique case (lizzieLet13_5QNode_Int_9_d[2:1])
        2'd0: q2aeS_destruct_onehotd = 4'd1;
        2'd1: q2aeS_destruct_onehotd = 4'd2;
        2'd2: q2aeS_destruct_onehotd = 4'd4;
        2'd3: q2aeS_destruct_onehotd = 4'd8;
        default: q2aeS_destruct_onehotd = 4'd0;
      endcase
    else q2aeS_destruct_onehotd = 4'd0;
  assign _135_d = {q2aeS_destruct_d[16:1],
                   q2aeS_destruct_onehotd[0]};
  assign _134_d = {q2aeS_destruct_d[16:1],
                   q2aeS_destruct_onehotd[1]};
  assign lizzieLet13_5QNode_Int_9QNode_Int_d = {q2aeS_destruct_d[16:1],
                                                q2aeS_destruct_onehotd[2]};
  assign _133_d = {q2aeS_destruct_d[16:1],
                   q2aeS_destruct_onehotd[3]};
  assign q2aeS_destruct_r = (| (q2aeS_destruct_onehotd & {_133_r,
                                                          lizzieLet13_5QNode_Int_9QNode_Int_r,
                                                          _134_r,
                                                          _135_r}));
  assign lizzieLet13_5QNode_Int_9_r = q2aeS_destruct_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet13_5QVal_Int,QTree_Int) > [(lizzieLet13_5QVal_Int_1,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_2,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_3,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_4,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_5,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_6,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_7,QTree_Int),
                                                           (lizzieLet13_5QVal_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet13_5QVal_Int_emitted;
  logic [7:0] lizzieLet13_5QVal_Int_done;
  assign lizzieLet13_5QVal_Int_1_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[0]))};
  assign lizzieLet13_5QVal_Int_2_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[1]))};
  assign lizzieLet13_5QVal_Int_3_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[2]))};
  assign lizzieLet13_5QVal_Int_4_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[3]))};
  assign lizzieLet13_5QVal_Int_5_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[4]))};
  assign lizzieLet13_5QVal_Int_6_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[5]))};
  assign lizzieLet13_5QVal_Int_7_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[6]))};
  assign lizzieLet13_5QVal_Int_8_d = {lizzieLet13_5QVal_Int_d[66:1],
                                      (lizzieLet13_5QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_emitted[7]))};
  assign lizzieLet13_5QVal_Int_done = (lizzieLet13_5QVal_Int_emitted | ({lizzieLet13_5QVal_Int_8_d[0],
                                                                         lizzieLet13_5QVal_Int_7_d[0],
                                                                         lizzieLet13_5QVal_Int_6_d[0],
                                                                         lizzieLet13_5QVal_Int_5_d[0],
                                                                         lizzieLet13_5QVal_Int_4_d[0],
                                                                         lizzieLet13_5QVal_Int_3_d[0],
                                                                         lizzieLet13_5QVal_Int_2_d[0],
                                                                         lizzieLet13_5QVal_Int_1_d[0]} & {lizzieLet13_5QVal_Int_8_r,
                                                                                                          lizzieLet13_5QVal_Int_7_r,
                                                                                                          lizzieLet13_5QVal_Int_6_r,
                                                                                                          lizzieLet13_5QVal_Int_5_r,
                                                                                                          lizzieLet13_5QVal_Int_4_r,
                                                                                                          lizzieLet13_5QVal_Int_3_r,
                                                                                                          lizzieLet13_5QVal_Int_2_r,
                                                                                                          lizzieLet13_5QVal_Int_1_r}));
  assign lizzieLet13_5QVal_Int_r = (& lizzieLet13_5QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_5QVal_Int_emitted <= 8'd0;
    else
      lizzieLet13_5QVal_Int_emitted <= (lizzieLet13_5QVal_Int_r ? 8'd0 :
                                        lizzieLet13_5QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet13_5QVal_Int_1QVal_Int,QTree_Int) > [(vaeM_destruct,Int)] */
  assign vaeM_destruct_d = {lizzieLet13_5QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet13_5QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet13_5QVal_Int_1QVal_Int_r = vaeM_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet13_5QVal_Int_2,QTree_Int) (lizzieLet13_5QVal_Int_1,QTree_Int) > [(_132,QTree_Int),
                                                                                                  (lizzieLet13_5QVal_Int_1QVal_Int,QTree_Int),
                                                                                                  (_131,QTree_Int),
                                                                                                  (_130,QTree_Int)] */
  logic [3:0] lizzieLet13_5QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_2_d[0] && lizzieLet13_5QVal_Int_1_d[0]))
      unique case (lizzieLet13_5QVal_Int_2_d[2:1])
        2'd0: lizzieLet13_5QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet13_5QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet13_5QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet13_5QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet13_5QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet13_5QVal_Int_1_onehotd = 4'd0;
  assign _132_d = {lizzieLet13_5QVal_Int_1_d[66:1],
                   lizzieLet13_5QVal_Int_1_onehotd[0]};
  assign lizzieLet13_5QVal_Int_1QVal_Int_d = {lizzieLet13_5QVal_Int_1_d[66:1],
                                              lizzieLet13_5QVal_Int_1_onehotd[1]};
  assign _131_d = {lizzieLet13_5QVal_Int_1_d[66:1],
                   lizzieLet13_5QVal_Int_1_onehotd[2]};
  assign _130_d = {lizzieLet13_5QVal_Int_1_d[66:1],
                   lizzieLet13_5QVal_Int_1_onehotd[3]};
  assign lizzieLet13_5QVal_Int_1_r = (| (lizzieLet13_5QVal_Int_1_onehotd & {_130_r,
                                                                            _131_r,
                                                                            lizzieLet13_5QVal_Int_1QVal_Int_r,
                                                                            _132_r}));
  assign lizzieLet13_5QVal_Int_2_r = lizzieLet13_5QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet13_5QVal_Int_3,QTree_Int) (lizzieLet13_3QVal_Int,Go) > [(lizzieLet13_5QVal_Int_3QNone_Int,Go),
                                                                                  (lizzieLet13_5QVal_Int_3QVal_Int,Go),
                                                                                  (lizzieLet13_5QVal_Int_3QNode_Int,Go),
                                                                                  (lizzieLet13_5QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet13_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_3_d[0] && lizzieLet13_3QVal_Int_d[0]))
      unique case (lizzieLet13_5QVal_Int_3_d[2:1])
        2'd0: lizzieLet13_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet13_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet13_5QVal_Int_3QNone_Int_d = lizzieLet13_3QVal_Int_onehotd[0];
  assign lizzieLet13_5QVal_Int_3QVal_Int_d = lizzieLet13_3QVal_Int_onehotd[1];
  assign lizzieLet13_5QVal_Int_3QNode_Int_d = lizzieLet13_3QVal_Int_onehotd[2];
  assign lizzieLet13_5QVal_Int_3QError_Int_d = lizzieLet13_3QVal_Int_onehotd[3];
  assign lizzieLet13_3QVal_Int_r = (| (lizzieLet13_3QVal_Int_onehotd & {lizzieLet13_5QVal_Int_3QError_Int_r,
                                                                        lizzieLet13_5QVal_Int_3QNode_Int_r,
                                                                        lizzieLet13_5QVal_Int_3QVal_Int_r,
                                                                        lizzieLet13_5QVal_Int_3QNone_Int_r}));
  assign lizzieLet13_5QVal_Int_3_r = lizzieLet13_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet13_5QVal_Int_3QError_Int,Go) > [(lizzieLet13_5QVal_Int_3QError_Int_1,Go),
                                                         (lizzieLet13_5QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet13_5QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet13_5QVal_Int_3QError_Int_done;
  assign lizzieLet13_5QVal_Int_3QError_Int_1_d = (lizzieLet13_5QVal_Int_3QError_Int_d[0] && (! lizzieLet13_5QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet13_5QVal_Int_3QError_Int_2_d = (lizzieLet13_5QVal_Int_3QError_Int_d[0] && (! lizzieLet13_5QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet13_5QVal_Int_3QError_Int_done = (lizzieLet13_5QVal_Int_3QError_Int_emitted | ({lizzieLet13_5QVal_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet13_5QVal_Int_3QError_Int_1_d[0]} & {lizzieLet13_5QVal_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet13_5QVal_Int_3QError_Int_1_r}));
  assign lizzieLet13_5QVal_Int_3QError_Int_r = (& lizzieLet13_5QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QVal_Int_3QError_Int_emitted <= (lizzieLet13_5QVal_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet13_5QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_5QVal_Int_3QError_Int_1,Go)] > (lizzieLet13_5QVal_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_5QVal_Int_3QError_Int_1_d[0]}), lizzieLet13_5QVal_Int_3QError_Int_1_d);
  assign {lizzieLet13_5QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_r && lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_5QVal_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet18_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_r = ((! lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_r)
        lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet13_5QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QVal_Int_3QError_Int_2,Go) > (lizzieLet13_5QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QError_Int_2_r = ((! lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_3QError_Int_2_r)
        lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet13_5QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_r && lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet13_5QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet13_5QVal_Int_3QNode_Int,Go) > [(lizzieLet13_5QVal_Int_3QNode_Int_1,Go),
                                                        (lizzieLet13_5QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet13_5QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet13_5QVal_Int_3QNode_Int_done;
  assign lizzieLet13_5QVal_Int_3QNode_Int_1_d = (lizzieLet13_5QVal_Int_3QNode_Int_d[0] && (! lizzieLet13_5QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet13_5QVal_Int_3QNode_Int_2_d = (lizzieLet13_5QVal_Int_3QNode_Int_d[0] && (! lizzieLet13_5QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet13_5QVal_Int_3QNode_Int_done = (lizzieLet13_5QVal_Int_3QNode_Int_emitted | ({lizzieLet13_5QVal_Int_3QNode_Int_2_d[0],
                                                                                               lizzieLet13_5QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet13_5QVal_Int_3QNode_Int_2_r,
                                                                                                                                           lizzieLet13_5QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet13_5QVal_Int_3QNode_Int_r = (& lizzieLet13_5QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QVal_Int_3QNode_Int_emitted <= (lizzieLet13_5QVal_Int_3QNode_Int_r ? 2'd0 :
                                                   lizzieLet13_5QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_5QVal_Int_3QNode_Int_1,Go)] > (lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_5QVal_Int_3QNode_Int_1_d[0]}), lizzieLet13_5QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet13_5QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_r && lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int,QTree_Int) > (lizzieLet17_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_r = ((! lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_r)
        lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_r = (! lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= lizzieLet13_5QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QVal_Int_3QNode_Int_2,Go) > (lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QNode_Int_2_r = ((! lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_3QNode_Int_2_r)
        lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet13_5QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf :
                                                        lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet13_5QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_5QVal_Int_3QNone_Int,Go) > (lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QNone_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QNone_Int_r = ((! lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_3QNone_Int_r)
        lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d <= lizzieLet13_5QVal_Int_3QNone_Int_d;
  Go_t lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QNone_Int_bufchan_r = (! lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf :
                                                        lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QNone_Int_bufchan_buf <= lizzieLet13_5QVal_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet13_5QVal_Int_3QVal_Int,Go) > [(lizzieLet13_5QVal_Int_3QVal_Int_1,Go),
                                                       (lizzieLet13_5QVal_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet13_5QVal_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet13_5QVal_Int_3QVal_Int_done;
  assign lizzieLet13_5QVal_Int_3QVal_Int_1_d = (lizzieLet13_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_3QVal_Int_emitted[0]));
  assign lizzieLet13_5QVal_Int_3QVal_Int_2_d = (lizzieLet13_5QVal_Int_3QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_3QVal_Int_emitted[1]));
  assign lizzieLet13_5QVal_Int_3QVal_Int_done = (lizzieLet13_5QVal_Int_3QVal_Int_emitted | ({lizzieLet13_5QVal_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet13_5QVal_Int_3QVal_Int_1_d[0]} & {lizzieLet13_5QVal_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet13_5QVal_Int_3QVal_Int_1_r}));
  assign lizzieLet13_5QVal_Int_3QVal_Int_r = (& lizzieLet13_5QVal_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QVal_Int_3QVal_Int_emitted <= (lizzieLet13_5QVal_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet13_5QVal_Int_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet13_5QVal_Int_3QVal_Int_1,Go) > (lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d;
  logic lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_r;
  assign lizzieLet13_5QVal_Int_3QVal_Int_1_r = ((! lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d[0]) || lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_3QVal_Int_1_r)
        lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d <= lizzieLet13_5QVal_Int_3QVal_Int_1_d;
  Go_t lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf;
  assign lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_r = (! lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf[0] ? lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf :
                                                       lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_buf <= lizzieLet13_5QVal_Int_3QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf,Go),
                                          (lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_d[0],
                                                                                             es_1_1_argbuf_d[0]}), lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_d, lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_d, es_1_1_argbuf_d);
  assign {lizzieLet13_5QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_r,
          es_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet13_5QVal_Int_4,QTree_Int) (lizzieLet13_4QVal_Int,MyDTInt_Bool) > [(_129,MyDTInt_Bool),
                                                                                                      (lizzieLet13_5QVal_Int_4QVal_Int,MyDTInt_Bool),
                                                                                                      (_128,MyDTInt_Bool),
                                                                                                      (_127,MyDTInt_Bool)] */
  logic [3:0] lizzieLet13_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_4_d[0] && lizzieLet13_4QVal_Int_d[0]))
      unique case (lizzieLet13_5QVal_Int_4_d[2:1])
        2'd0: lizzieLet13_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet13_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_4QVal_Int_onehotd = 4'd0;
  assign _129_d = lizzieLet13_4QVal_Int_onehotd[0];
  assign lizzieLet13_5QVal_Int_4QVal_Int_d = lizzieLet13_4QVal_Int_onehotd[1];
  assign _128_d = lizzieLet13_4QVal_Int_onehotd[2];
  assign _127_d = lizzieLet13_4QVal_Int_onehotd[3];
  assign lizzieLet13_4QVal_Int_r = (| (lizzieLet13_4QVal_Int_onehotd & {_127_r,
                                                                        _128_r,
                                                                        lizzieLet13_5QVal_Int_4QVal_Int_r,
                                                                        _129_r}));
  assign lizzieLet13_5QVal_Int_4_r = lizzieLet13_4QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_5QVal_Int_4QVal_Int,MyDTInt_Bool) > (lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_4QVal_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_4QVal_Int_r = ((! lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_4QVal_Int_r)
        lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d <= lizzieLet13_5QVal_Int_4QVal_Int_d;
  MyDTInt_Bool_t lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_4QVal_Int_bufchan_r = (! lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf :
                                                       lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_4QVal_Int_bufchan_buf <= lizzieLet13_5QVal_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_5QVal_Int_5,QTree_Int) (lizzieLet13_6QVal_Int,Pointer_QTree_Int) > [(lizzieLet13_5QVal_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                                (_126,Pointer_QTree_Int),
                                                                                                                (_125,Pointer_QTree_Int),
                                                                                                                (_124,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet13_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_5_d[0] && lizzieLet13_6QVal_Int_d[0]))
      unique case (lizzieLet13_5QVal_Int_5_d[2:1])
        2'd0: lizzieLet13_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet13_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_6QVal_Int_onehotd = 4'd0;
  assign lizzieLet13_5QVal_Int_5QNone_Int_d = {lizzieLet13_6QVal_Int_d[16:1],
                                               lizzieLet13_6QVal_Int_onehotd[0]};
  assign _126_d = {lizzieLet13_6QVal_Int_d[16:1],
                   lizzieLet13_6QVal_Int_onehotd[1]};
  assign _125_d = {lizzieLet13_6QVal_Int_d[16:1],
                   lizzieLet13_6QVal_Int_onehotd[2]};
  assign _124_d = {lizzieLet13_6QVal_Int_d[16:1],
                   lizzieLet13_6QVal_Int_onehotd[3]};
  assign lizzieLet13_6QVal_Int_r = (| (lizzieLet13_6QVal_Int_onehotd & {_124_r,
                                                                        _125_r,
                                                                        _126_r,
                                                                        lizzieLet13_5QVal_Int_5QNone_Int_r}));
  assign lizzieLet13_5QVal_Int_5_r = lizzieLet13_6QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_5QVal_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_5QNone_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_5QNone_Int_r = ((! lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QVal_Int_5QNone_Int_r)
        lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d <= lizzieLet13_5QVal_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_5QNone_Int_bufchan_r = (! lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf :
                                                        lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_r && lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QVal_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_5QNone_Int_bufchan_buf <= lizzieLet13_5QVal_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet13_5QVal_Int_6,QTree_Int) (lizzieLet13_8QVal_Int,MyDTInt_Int_Int) > [(_123,MyDTInt_Int_Int),
                                                                                                            (lizzieLet13_5QVal_Int_6QVal_Int,MyDTInt_Int_Int),
                                                                                                            (_122,MyDTInt_Int_Int),
                                                                                                            (_121,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet13_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_6_d[0] && lizzieLet13_8QVal_Int_d[0]))
      unique case (lizzieLet13_5QVal_Int_6_d[2:1])
        2'd0: lizzieLet13_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet13_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_8QVal_Int_onehotd = 4'd0;
  assign _123_d = lizzieLet13_8QVal_Int_onehotd[0];
  assign lizzieLet13_5QVal_Int_6QVal_Int_d = lizzieLet13_8QVal_Int_onehotd[1];
  assign _122_d = lizzieLet13_8QVal_Int_onehotd[2];
  assign _121_d = lizzieLet13_8QVal_Int_onehotd[3];
  assign lizzieLet13_8QVal_Int_r = (| (lizzieLet13_8QVal_Int_onehotd & {_121_r,
                                                                        _122_r,
                                                                        lizzieLet13_5QVal_Int_6QVal_Int_r,
                                                                        _123_r}));
  assign lizzieLet13_5QVal_Int_6_r = lizzieLet13_8QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet13_5QVal_Int_6QVal_Int,MyDTInt_Int_Int) > [(lizzieLet13_5QVal_Int_6QVal_Int_1,MyDTInt_Int_Int),
                                                                                 (lizzieLet13_5QVal_Int_6QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet13_5QVal_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet13_5QVal_Int_6QVal_Int_done;
  assign lizzieLet13_5QVal_Int_6QVal_Int_1_d = (lizzieLet13_5QVal_Int_6QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_6QVal_Int_emitted[0]));
  assign lizzieLet13_5QVal_Int_6QVal_Int_2_d = (lizzieLet13_5QVal_Int_6QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_6QVal_Int_emitted[1]));
  assign lizzieLet13_5QVal_Int_6QVal_Int_done = (lizzieLet13_5QVal_Int_6QVal_Int_emitted | ({lizzieLet13_5QVal_Int_6QVal_Int_2_d[0],
                                                                                             lizzieLet13_5QVal_Int_6QVal_Int_1_d[0]} & {lizzieLet13_5QVal_Int_6QVal_Int_2_r,
                                                                                                                                        lizzieLet13_5QVal_Int_6QVal_Int_1_r}));
  assign lizzieLet13_5QVal_Int_6QVal_Int_r = (& lizzieLet13_5QVal_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QVal_Int_6QVal_Int_emitted <= (lizzieLet13_5QVal_Int_6QVal_Int_r ? 2'd0 :
                                                  lizzieLet13_5QVal_Int_6QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet13_5QVal_Int_6QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d;
  logic lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_r;
  assign lizzieLet13_5QVal_Int_6QVal_Int_1_r = ((! lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d[0]) || lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_5QVal_Int_6QVal_Int_1_r)
        lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d <= lizzieLet13_5QVal_Int_6QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf;
  assign lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_r = (! lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf[0] ? lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf :
                                                       lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_buf <= lizzieLet13_5QVal_Int_6QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf,Int),
                                              (vaeM_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_d[0],
                                                                                                        vaeM_1_argbuf_d[0]}), lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_d, lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_d, vaeM_1_argbuf_d);
  assign {lizzieLet13_5QVal_Int_6QVal_Int_1_argbuf_r,
          lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_r,
          vaeM_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QVal_Int_7,QTree_Int) (lizzieLet13_9QVal_Int,Pointer_CTf'_f'_Int) > [(lizzieLet13_5QVal_Int_7QNone_Int,Pointer_CTf'_f'_Int),
                                                                                                                    (lizzieLet13_5QVal_Int_7QVal_Int,Pointer_CTf'_f'_Int),
                                                                                                                    (lizzieLet13_5QVal_Int_7QNode_Int,Pointer_CTf'_f'_Int),
                                                                                                                    (lizzieLet13_5QVal_Int_7QError_Int,Pointer_CTf'_f'_Int)] */
  logic [3:0] lizzieLet13_9QVal_Int_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_7_d[0] && lizzieLet13_9QVal_Int_d[0]))
      unique case (lizzieLet13_5QVal_Int_7_d[2:1])
        2'd0: lizzieLet13_9QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet13_9QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet13_9QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet13_9QVal_Int_onehotd = 4'd8;
        default: lizzieLet13_9QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet13_9QVal_Int_onehotd = 4'd0;
  assign lizzieLet13_5QVal_Int_7QNone_Int_d = {lizzieLet13_9QVal_Int_d[16:1],
                                               lizzieLet13_9QVal_Int_onehotd[0]};
  assign lizzieLet13_5QVal_Int_7QVal_Int_d = {lizzieLet13_9QVal_Int_d[16:1],
                                              lizzieLet13_9QVal_Int_onehotd[1]};
  assign lizzieLet13_5QVal_Int_7QNode_Int_d = {lizzieLet13_9QVal_Int_d[16:1],
                                               lizzieLet13_9QVal_Int_onehotd[2]};
  assign lizzieLet13_5QVal_Int_7QError_Int_d = {lizzieLet13_9QVal_Int_d[16:1],
                                                lizzieLet13_9QVal_Int_onehotd[3]};
  assign lizzieLet13_9QVal_Int_r = (| (lizzieLet13_9QVal_Int_onehotd & {lizzieLet13_5QVal_Int_7QError_Int_r,
                                                                        lizzieLet13_5QVal_Int_7QNode_Int_r,
                                                                        lizzieLet13_5QVal_Int_7QVal_Int_r,
                                                                        lizzieLet13_5QVal_Int_7QNone_Int_r}));
  assign lizzieLet13_5QVal_Int_7_r = lizzieLet13_9QVal_Int_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QVal_Int_7QError_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QVal_Int_7QError_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QError_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_7QError_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_7QError_Int_r = ((! lizzieLet13_5QVal_Int_7QError_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_7QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QVal_Int_7QError_Int_r)
        lizzieLet13_5QVal_Int_7QError_Int_bufchan_d <= lizzieLet13_5QVal_Int_7QError_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_7QError_Int_bufchan_r = (! lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf :
                                                         lizzieLet13_5QVal_Int_7QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_r && lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QVal_Int_7QError_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_7QError_Int_bufchan_buf <= lizzieLet13_5QVal_Int_7QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QVal_Int_7QNode_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_7QNode_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_7QNode_Int_r = ((! lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_7QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QVal_Int_7QNode_Int_r)
        lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d <= lizzieLet13_5QVal_Int_7QNode_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_7QNode_Int_bufchan_r = (! lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf :
                                                        lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_r && lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QVal_Int_7QNode_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_7QNode_Int_bufchan_buf <= lizzieLet13_5QVal_Int_7QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_5QVal_Int_7QNone_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d;
  logic lizzieLet13_5QVal_Int_7QNone_Int_bufchan_r;
  assign lizzieLet13_5QVal_Int_7QNone_Int_r = ((! lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d[0]) || lizzieLet13_5QVal_Int_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_5QVal_Int_7QNone_Int_r)
        lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d <= lizzieLet13_5QVal_Int_7QNone_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf;
  assign lizzieLet13_5QVal_Int_7QNone_Int_bufchan_r = (! lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf[0] ? lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf :
                                                        lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_r && lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_5QVal_Int_7QNone_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_7QNone_Int_bufchan_buf <= lizzieLet13_5QVal_Int_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet13_5QVal_Int_8,QTree_Int) (v1aeL_destruct,Int) > [(_120,Int),
                                                                             (lizzieLet13_5QVal_Int_8QVal_Int,Int),
                                                                             (_119,Int),
                                                                             (_118,Int)] */
  logic [3:0] v1aeL_destruct_onehotd;
  always_comb
    if ((lizzieLet13_5QVal_Int_8_d[0] && v1aeL_destruct_d[0]))
      unique case (lizzieLet13_5QVal_Int_8_d[2:1])
        2'd0: v1aeL_destruct_onehotd = 4'd1;
        2'd1: v1aeL_destruct_onehotd = 4'd2;
        2'd2: v1aeL_destruct_onehotd = 4'd4;
        2'd3: v1aeL_destruct_onehotd = 4'd8;
        default: v1aeL_destruct_onehotd = 4'd0;
      endcase
    else v1aeL_destruct_onehotd = 4'd0;
  assign _120_d = {v1aeL_destruct_d[32:1],
                   v1aeL_destruct_onehotd[0]};
  assign lizzieLet13_5QVal_Int_8QVal_Int_d = {v1aeL_destruct_d[32:1],
                                              v1aeL_destruct_onehotd[1]};
  assign _119_d = {v1aeL_destruct_d[32:1],
                   v1aeL_destruct_onehotd[2]};
  assign _118_d = {v1aeL_destruct_d[32:1],
                   v1aeL_destruct_onehotd[3]};
  assign v1aeL_destruct_r = (| (v1aeL_destruct_onehotd & {_118_r,
                                                          _119_r,
                                                          lizzieLet13_5QVal_Int_8QVal_Int_r,
                                                          _120_r}));
  assign lizzieLet13_5QVal_Int_8_r = v1aeL_destruct_r;
  
  /* fork (Ty Int) : (lizzieLet13_5QVal_Int_8QVal_Int,Int) > [(lizzieLet13_5QVal_Int_8QVal_Int_1,Int),
                                                         (lizzieLet13_5QVal_Int_8QVal_Int_2,Int)] */
  logic [1:0] lizzieLet13_5QVal_Int_8QVal_Int_emitted;
  logic [1:0] lizzieLet13_5QVal_Int_8QVal_Int_done;
  assign lizzieLet13_5QVal_Int_8QVal_Int_1_d = {lizzieLet13_5QVal_Int_8QVal_Int_d[32:1],
                                                (lizzieLet13_5QVal_Int_8QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_8QVal_Int_emitted[0]))};
  assign lizzieLet13_5QVal_Int_8QVal_Int_2_d = {lizzieLet13_5QVal_Int_8QVal_Int_d[32:1],
                                                (lizzieLet13_5QVal_Int_8QVal_Int_d[0] && (! lizzieLet13_5QVal_Int_8QVal_Int_emitted[1]))};
  assign lizzieLet13_5QVal_Int_8QVal_Int_done = (lizzieLet13_5QVal_Int_8QVal_Int_emitted | ({lizzieLet13_5QVal_Int_8QVal_Int_2_d[0],
                                                                                             lizzieLet13_5QVal_Int_8QVal_Int_1_d[0]} & {lizzieLet13_5QVal_Int_8QVal_Int_2_r,
                                                                                                                                        lizzieLet13_5QVal_Int_8QVal_Int_1_r}));
  assign lizzieLet13_5QVal_Int_8QVal_Int_r = (& lizzieLet13_5QVal_Int_8QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_8QVal_Int_emitted <= 2'd0;
    else
      lizzieLet13_5QVal_Int_8QVal_Int_emitted <= (lizzieLet13_5QVal_Int_8QVal_Int_r ? 2'd0 :
                                                  lizzieLet13_5QVal_Int_8QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet13_5QVal_Int_8QVal_Int_1,Int) > (lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d;
  logic lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_r;
  assign lizzieLet13_5QVal_Int_8QVal_Int_1_r = ((! lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d[0]) || lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet13_5QVal_Int_8QVal_Int_1_r)
        lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d <= lizzieLet13_5QVal_Int_8QVal_Int_1_d;
  Int_t lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf;
  assign lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_r = (! lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_d = (lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf[0] ? lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf :
                                                       lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_r && lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf[0]))
        lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet13_5QVal_Int_8QVal_Int_1_argbuf_r) && (! lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf[0])))
        lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_buf <= lizzieLet13_5QVal_Int_8QVal_Int_1_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_6,QTree_Int) (m2aeH_2,Pointer_QTree_Int) > [(_117,Pointer_QTree_Int),
                                                                                        (lizzieLet13_6QVal_Int,Pointer_QTree_Int),
                                                                                        (lizzieLet13_6QNode_Int,Pointer_QTree_Int),
                                                                                        (_116,Pointer_QTree_Int)] */
  logic [3:0] m2aeH_2_onehotd;
  always_comb
    if ((lizzieLet13_6_d[0] && m2aeH_2_d[0]))
      unique case (lizzieLet13_6_d[2:1])
        2'd0: m2aeH_2_onehotd = 4'd1;
        2'd1: m2aeH_2_onehotd = 4'd2;
        2'd2: m2aeH_2_onehotd = 4'd4;
        2'd3: m2aeH_2_onehotd = 4'd8;
        default: m2aeH_2_onehotd = 4'd0;
      endcase
    else m2aeH_2_onehotd = 4'd0;
  assign _117_d = {m2aeH_2_d[16:1], m2aeH_2_onehotd[0]};
  assign lizzieLet13_6QVal_Int_d = {m2aeH_2_d[16:1],
                                    m2aeH_2_onehotd[1]};
  assign lizzieLet13_6QNode_Int_d = {m2aeH_2_d[16:1],
                                     m2aeH_2_onehotd[2]};
  assign _116_d = {m2aeH_2_d[16:1], m2aeH_2_onehotd[3]};
  assign m2aeH_2_r = (| (m2aeH_2_onehotd & {_116_r,
                                            lizzieLet13_6QNode_Int_r,
                                            lizzieLet13_6QVal_Int_r,
                                            _117_r}));
  assign lizzieLet13_6_r = m2aeH_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_7,QTree_Int) (m3aeI_2,Pointer_QTree_Int) > [(lizzieLet13_7QNone_Int,Pointer_QTree_Int),
                                                                                        (_115,Pointer_QTree_Int),
                                                                                        (_114,Pointer_QTree_Int),
                                                                                        (_113,Pointer_QTree_Int)] */
  logic [3:0] m3aeI_2_onehotd;
  always_comb
    if ((lizzieLet13_7_d[0] && m3aeI_2_d[0]))
      unique case (lizzieLet13_7_d[2:1])
        2'd0: m3aeI_2_onehotd = 4'd1;
        2'd1: m3aeI_2_onehotd = 4'd2;
        2'd2: m3aeI_2_onehotd = 4'd4;
        2'd3: m3aeI_2_onehotd = 4'd8;
        default: m3aeI_2_onehotd = 4'd0;
      endcase
    else m3aeI_2_onehotd = 4'd0;
  assign lizzieLet13_7QNone_Int_d = {m3aeI_2_d[16:1],
                                     m3aeI_2_onehotd[0]};
  assign _115_d = {m3aeI_2_d[16:1], m3aeI_2_onehotd[1]};
  assign _114_d = {m3aeI_2_d[16:1], m3aeI_2_onehotd[2]};
  assign _113_d = {m3aeI_2_d[16:1], m3aeI_2_onehotd[3]};
  assign m3aeI_2_r = (| (m3aeI_2_onehotd & {_113_r,
                                            _114_r,
                                            _115_r,
                                            lizzieLet13_7QNone_Int_r}));
  assign lizzieLet13_7_r = m3aeI_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_7QNone_Int,Pointer_QTree_Int) > (lizzieLet13_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_7QNone_Int_bufchan_d;
  logic lizzieLet13_7QNone_Int_bufchan_r;
  assign lizzieLet13_7QNone_Int_r = ((! lizzieLet13_7QNone_Int_bufchan_d[0]) || lizzieLet13_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_7QNone_Int_r)
        lizzieLet13_7QNone_Int_bufchan_d <= lizzieLet13_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet13_7QNone_Int_bufchan_buf;
  assign lizzieLet13_7QNone_Int_bufchan_r = (! lizzieLet13_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_7QNone_Int_1_argbuf_d = (lizzieLet13_7QNone_Int_bufchan_buf[0] ? lizzieLet13_7QNone_Int_bufchan_buf :
                                              lizzieLet13_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_7QNone_Int_1_argbuf_r && lizzieLet13_7QNone_Int_bufchan_buf[0]))
        lizzieLet13_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_7QNone_Int_1_argbuf_r) && (! lizzieLet13_7QNone_Int_bufchan_buf[0])))
        lizzieLet13_7QNone_Int_bufchan_buf <= lizzieLet13_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet13_8,QTree_Int) (op_addaeK_goMux_mux,MyDTInt_Int_Int) > [(_112,MyDTInt_Int_Int),
                                                                                                (lizzieLet13_8QVal_Int,MyDTInt_Int_Int),
                                                                                                (lizzieLet13_8QNode_Int,MyDTInt_Int_Int),
                                                                                                (_111,MyDTInt_Int_Int)] */
  logic [3:0] op_addaeK_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_8_d[0] && op_addaeK_goMux_mux_d[0]))
      unique case (lizzieLet13_8_d[2:1])
        2'd0: op_addaeK_goMux_mux_onehotd = 4'd1;
        2'd1: op_addaeK_goMux_mux_onehotd = 4'd2;
        2'd2: op_addaeK_goMux_mux_onehotd = 4'd4;
        2'd3: op_addaeK_goMux_mux_onehotd = 4'd8;
        default: op_addaeK_goMux_mux_onehotd = 4'd0;
      endcase
    else op_addaeK_goMux_mux_onehotd = 4'd0;
  assign _112_d = op_addaeK_goMux_mux_onehotd[0];
  assign lizzieLet13_8QVal_Int_d = op_addaeK_goMux_mux_onehotd[1];
  assign lizzieLet13_8QNode_Int_d = op_addaeK_goMux_mux_onehotd[2];
  assign _111_d = op_addaeK_goMux_mux_onehotd[3];
  assign op_addaeK_goMux_mux_r = (| (op_addaeK_goMux_mux_onehotd & {_111_r,
                                                                    lizzieLet13_8QNode_Int_r,
                                                                    lizzieLet13_8QVal_Int_r,
                                                                    _112_r}));
  assign lizzieLet13_8_r = op_addaeK_goMux_mux_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf'_f'_Int) : (lizzieLet13_9,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTf'_f'_Int) > [(lizzieLet13_9QNone_Int,Pointer_CTf'_f'_Int),
                                                                                                     (lizzieLet13_9QVal_Int,Pointer_CTf'_f'_Int),
                                                                                                     (lizzieLet13_9QNode_Int,Pointer_CTf'_f'_Int),
                                                                                                     (lizzieLet13_9QError_Int,Pointer_CTf'_f'_Int)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_9_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet13_9_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet13_9QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet13_9QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet13_9QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet13_9QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet13_9QError_Int_r,
                                                              lizzieLet13_9QNode_Int_r,
                                                              lizzieLet13_9QVal_Int_r,
                                                              lizzieLet13_9QNone_Int_r}));
  assign lizzieLet13_9_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_9QError_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_9QError_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QError_Int_bufchan_d;
  logic lizzieLet13_9QError_Int_bufchan_r;
  assign lizzieLet13_9QError_Int_r = ((! lizzieLet13_9QError_Int_bufchan_d[0]) || lizzieLet13_9QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_9QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_9QError_Int_r)
        lizzieLet13_9QError_Int_bufchan_d <= lizzieLet13_9QError_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QError_Int_bufchan_buf;
  assign lizzieLet13_9QError_Int_bufchan_r = (! lizzieLet13_9QError_Int_bufchan_buf[0]);
  assign lizzieLet13_9QError_Int_1_argbuf_d = (lizzieLet13_9QError_Int_bufchan_buf[0] ? lizzieLet13_9QError_Int_bufchan_buf :
                                               lizzieLet13_9QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_9QError_Int_1_argbuf_r && lizzieLet13_9QError_Int_bufchan_buf[0]))
        lizzieLet13_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_9QError_Int_1_argbuf_r) && (! lizzieLet13_9QError_Int_bufchan_buf[0])))
        lizzieLet13_9QError_Int_bufchan_buf <= lizzieLet13_9QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (lizzieLet13_9QNone_Int,Pointer_CTf'_f'_Int) > (lizzieLet13_9QNone_Int_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QNone_Int_bufchan_d;
  logic lizzieLet13_9QNone_Int_bufchan_r;
  assign lizzieLet13_9QNone_Int_r = ((! lizzieLet13_9QNone_Int_bufchan_d[0]) || lizzieLet13_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_9QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_9QNone_Int_r)
        lizzieLet13_9QNone_Int_bufchan_d <= lizzieLet13_9QNone_Int_d;
  \Pointer_CTf'_f'_Int_t  lizzieLet13_9QNone_Int_bufchan_buf;
  assign lizzieLet13_9QNone_Int_bufchan_r = (! lizzieLet13_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_9QNone_Int_1_argbuf_d = (lizzieLet13_9QNone_Int_bufchan_buf[0] ? lizzieLet13_9QNone_Int_bufchan_buf :
                                              lizzieLet13_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_9QNone_Int_1_argbuf_r && lizzieLet13_9QNone_Int_bufchan_buf[0]))
        lizzieLet13_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_9QNone_Int_1_argbuf_r) && (! lizzieLet13_9QNone_Int_bufchan_buf[0])))
        lizzieLet13_9QNone_Int_bufchan_buf <= lizzieLet13_9QNone_Int_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1Xt_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1Xt_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1Xt_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1Xt_1_Eq_r = ((! lizzieLet1_1wild1Xt_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1Xt_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xt_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1Xt_1_Eq_r)
        lizzieLet1_1wild1Xt_1_Eq_bufchan_d <= lizzieLet1_1wild1Xt_1_Eq_d;
  Bool_t lizzieLet1_1wild1Xt_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1Xt_1_Eq_bufchan_r = (! lizzieLet1_1wild1Xt_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1Xt_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1Xt_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1Xt_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1Xt_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1Xt_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1Xt_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1Xt_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1Xt_1_Eq_bufchan_buf <= lizzieLet1_1wild1Xt_1_Eq_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTf_f_Int) : (lizzieLet24_10,MaskQTree) (sc_0_3_goMux_mux,Pointer_CTf_f_Int) > [(lizzieLet24_10MQNone,Pointer_CTf_f_Int),
                                                                                                  (lizzieLet24_10MQVal,Pointer_CTf_f_Int),
                                                                                                  (lizzieLet24_10MQNode,Pointer_CTf_f_Int)] */
  logic [2:0] sc_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_10_d[0] && sc_0_3_goMux_mux_d[0]))
      unique case (lizzieLet24_10_d[2:1])
        2'd0: sc_0_3_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_3_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_3_goMux_mux_onehotd = 3'd4;
        default: sc_0_3_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_3_goMux_mux_onehotd = 3'd0;
  assign lizzieLet24_10MQNone_d = {sc_0_3_goMux_mux_d[16:1],
                                   sc_0_3_goMux_mux_onehotd[0]};
  assign lizzieLet24_10MQVal_d = {sc_0_3_goMux_mux_d[16:1],
                                  sc_0_3_goMux_mux_onehotd[1]};
  assign lizzieLet24_10MQNode_d = {sc_0_3_goMux_mux_d[16:1],
                                   sc_0_3_goMux_mux_onehotd[2]};
  assign sc_0_3_goMux_mux_r = (| (sc_0_3_goMux_mux_onehotd & {lizzieLet24_10MQNode_r,
                                                              lizzieLet24_10MQVal_r,
                                                              lizzieLet24_10MQNone_r}));
  assign lizzieLet24_10_r = sc_0_3_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_10MQNone,Pointer_CTf_f_Int) > (lizzieLet24_10MQNone_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_10MQNone_bufchan_d;
  logic lizzieLet24_10MQNone_bufchan_r;
  assign lizzieLet24_10MQNone_r = ((! lizzieLet24_10MQNone_bufchan_d[0]) || lizzieLet24_10MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_10MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet24_10MQNone_r)
        lizzieLet24_10MQNone_bufchan_d <= lizzieLet24_10MQNone_d;
  Pointer_CTf_f_Int_t lizzieLet24_10MQNone_bufchan_buf;
  assign lizzieLet24_10MQNone_bufchan_r = (! lizzieLet24_10MQNone_bufchan_buf[0]);
  assign lizzieLet24_10MQNone_1_argbuf_d = (lizzieLet24_10MQNone_bufchan_buf[0] ? lizzieLet24_10MQNone_bufchan_buf :
                                            lizzieLet24_10MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_10MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_10MQNone_1_argbuf_r && lizzieLet24_10MQNone_bufchan_buf[0]))
        lizzieLet24_10MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet24_10MQNone_1_argbuf_r) && (! lizzieLet24_10MQNone_bufchan_buf[0])))
        lizzieLet24_10MQNone_bufchan_buf <= lizzieLet24_10MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_10MQVal,Pointer_CTf_f_Int) > (lizzieLet24_10MQVal_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_10MQVal_bufchan_d;
  logic lizzieLet24_10MQVal_bufchan_r;
  assign lizzieLet24_10MQVal_r = ((! lizzieLet24_10MQVal_bufchan_d[0]) || lizzieLet24_10MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_10MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet24_10MQVal_r)
        lizzieLet24_10MQVal_bufchan_d <= lizzieLet24_10MQVal_d;
  Pointer_CTf_f_Int_t lizzieLet24_10MQVal_bufchan_buf;
  assign lizzieLet24_10MQVal_bufchan_r = (! lizzieLet24_10MQVal_bufchan_buf[0]);
  assign lizzieLet24_10MQVal_1_argbuf_d = (lizzieLet24_10MQVal_bufchan_buf[0] ? lizzieLet24_10MQVal_bufchan_buf :
                                           lizzieLet24_10MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_10MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_10MQVal_1_argbuf_r && lizzieLet24_10MQVal_bufchan_buf[0]))
        lizzieLet24_10MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet24_10MQVal_1_argbuf_r) && (! lizzieLet24_10MQVal_bufchan_buf[0])))
        lizzieLet24_10MQVal_bufchan_buf <= lizzieLet24_10MQVal_bufchan_d;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet24_1MQNode,MaskQTree) > [(q1ae8_destruct,Pointer_MaskQTree),
                                                            (q2ae9_destruct,Pointer_MaskQTree),
                                                            (q3aea_destruct,Pointer_MaskQTree),
                                                            (q4aeb_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_1MQNode_emitted;
  logic [3:0] lizzieLet24_1MQNode_done;
  assign q1ae8_destruct_d = {lizzieLet24_1MQNode_d[18:3],
                             (lizzieLet24_1MQNode_d[0] && (! lizzieLet24_1MQNode_emitted[0]))};
  assign q2ae9_destruct_d = {lizzieLet24_1MQNode_d[34:19],
                             (lizzieLet24_1MQNode_d[0] && (! lizzieLet24_1MQNode_emitted[1]))};
  assign q3aea_destruct_d = {lizzieLet24_1MQNode_d[50:35],
                             (lizzieLet24_1MQNode_d[0] && (! lizzieLet24_1MQNode_emitted[2]))};
  assign q4aeb_destruct_d = {lizzieLet24_1MQNode_d[66:51],
                             (lizzieLet24_1MQNode_d[0] && (! lizzieLet24_1MQNode_emitted[3]))};
  assign lizzieLet24_1MQNode_done = (lizzieLet24_1MQNode_emitted | ({q4aeb_destruct_d[0],
                                                                     q3aea_destruct_d[0],
                                                                     q2ae9_destruct_d[0],
                                                                     q1ae8_destruct_d[0]} & {q4aeb_destruct_r,
                                                                                             q3aea_destruct_r,
                                                                                             q2ae9_destruct_r,
                                                                                             q1ae8_destruct_r}));
  assign lizzieLet24_1MQNode_r = (& lizzieLet24_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_1MQNode_emitted <= 4'd0;
    else
      lizzieLet24_1MQNode_emitted <= (lizzieLet24_1MQNode_r ? 4'd0 :
                                      lizzieLet24_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet24_2,MaskQTree) (lizzieLet24_1,MaskQTree) > [(_110,MaskQTree),
                                                                              (_109,MaskQTree),
                                                                              (lizzieLet24_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet24_1_onehotd;
  always_comb
    if ((lizzieLet24_2_d[0] && lizzieLet24_1_d[0]))
      unique case (lizzieLet24_2_d[2:1])
        2'd0: lizzieLet24_1_onehotd = 3'd1;
        2'd1: lizzieLet24_1_onehotd = 3'd2;
        2'd2: lizzieLet24_1_onehotd = 3'd4;
        default: lizzieLet24_1_onehotd = 3'd0;
      endcase
    else lizzieLet24_1_onehotd = 3'd0;
  assign _110_d = {lizzieLet24_1_d[66:1], lizzieLet24_1_onehotd[0]};
  assign _109_d = {lizzieLet24_1_d[66:1], lizzieLet24_1_onehotd[1]};
  assign lizzieLet24_1MQNode_d = {lizzieLet24_1_d[66:1],
                                  lizzieLet24_1_onehotd[2]};
  assign lizzieLet24_1_r = (| (lizzieLet24_1_onehotd & {lizzieLet24_1MQNode_r,
                                                        _109_r,
                                                        _110_r}));
  assign lizzieLet24_2_r = lizzieLet24_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet24_3,MaskQTree) (go_11_goMux_data,Go) > [(lizzieLet24_3MQNone,Go),
                                                                   (lizzieLet24_3MQVal,Go),
                                                                   (lizzieLet24_3MQNode,Go)] */
  logic [2:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet24_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet24_3_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 3'd1;
        2'd1: go_11_goMux_data_onehotd = 3'd2;
        2'd2: go_11_goMux_data_onehotd = 3'd4;
        default: go_11_goMux_data_onehotd = 3'd0;
      endcase
    else go_11_goMux_data_onehotd = 3'd0;
  assign lizzieLet24_3MQNone_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet24_3MQVal_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet24_3MQNode_d = go_11_goMux_data_onehotd[2];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet24_3MQNode_r,
                                                              lizzieLet24_3MQVal_r,
                                                              lizzieLet24_3MQNone_r}));
  assign lizzieLet24_3_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet24_3MQNone,Go) > [(lizzieLet24_3MQNone_1,Go),
                                           (lizzieLet24_3MQNone_2,Go)] */
  logic [1:0] lizzieLet24_3MQNone_emitted;
  logic [1:0] lizzieLet24_3MQNone_done;
  assign lizzieLet24_3MQNone_1_d = (lizzieLet24_3MQNone_d[0] && (! lizzieLet24_3MQNone_emitted[0]));
  assign lizzieLet24_3MQNone_2_d = (lizzieLet24_3MQNone_d[0] && (! lizzieLet24_3MQNone_emitted[1]));
  assign lizzieLet24_3MQNone_done = (lizzieLet24_3MQNone_emitted | ({lizzieLet24_3MQNone_2_d[0],
                                                                     lizzieLet24_3MQNone_1_d[0]} & {lizzieLet24_3MQNone_2_r,
                                                                                                    lizzieLet24_3MQNone_1_r}));
  assign lizzieLet24_3MQNone_r = (& lizzieLet24_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQNone_emitted <= 2'd0;
    else
      lizzieLet24_3MQNone_emitted <= (lizzieLet24_3MQNone_r ? 2'd0 :
                                      lizzieLet24_3MQNone_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet24_3MQNone_1,Go)] > (lizzieLet24_3MQNone_1QNone_Int,QTree_Int) */
  assign lizzieLet24_3MQNone_1QNone_Int_d = QNone_Int_dc((& {lizzieLet24_3MQNone_1_d[0]}), lizzieLet24_3MQNone_1_d);
  assign {lizzieLet24_3MQNone_1_r} = {1 {(lizzieLet24_3MQNone_1QNone_Int_r && lizzieLet24_3MQNone_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_3MQNone_1QNone_Int,QTree_Int) > (lizzieLet25_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_3MQNone_1QNone_Int_bufchan_d;
  logic lizzieLet24_3MQNone_1QNone_Int_bufchan_r;
  assign lizzieLet24_3MQNone_1QNone_Int_r = ((! lizzieLet24_3MQNone_1QNone_Int_bufchan_d[0]) || lizzieLet24_3MQNone_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3MQNone_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet24_3MQNone_1QNone_Int_r)
        lizzieLet24_3MQNone_1QNone_Int_bufchan_d <= lizzieLet24_3MQNone_1QNone_Int_d;
  QTree_Int_t lizzieLet24_3MQNone_1QNone_Int_bufchan_buf;
  assign lizzieLet24_3MQNone_1QNone_Int_bufchan_r = (! lizzieLet24_3MQNone_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet24_3MQNone_1QNone_Int_bufchan_buf[0] ? lizzieLet24_3MQNone_1QNone_Int_bufchan_buf :
                                   lizzieLet24_3MQNone_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet24_3MQNone_1QNone_Int_bufchan_buf[0]))
        lizzieLet24_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet24_3MQNone_1QNone_Int_bufchan_buf[0])))
        lizzieLet24_3MQNone_1QNone_Int_bufchan_buf <= lizzieLet24_3MQNone_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3MQNone_2,Go) > (lizzieLet24_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet24_3MQNone_2_bufchan_d;
  logic lizzieLet24_3MQNone_2_bufchan_r;
  assign lizzieLet24_3MQNone_2_r = ((! lizzieLet24_3MQNone_2_bufchan_d[0]) || lizzieLet24_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3MQNone_2_r)
        lizzieLet24_3MQNone_2_bufchan_d <= lizzieLet24_3MQNone_2_d;
  Go_t lizzieLet24_3MQNone_2_bufchan_buf;
  assign lizzieLet24_3MQNone_2_bufchan_r = (! lizzieLet24_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet24_3MQNone_2_argbuf_d = (lizzieLet24_3MQNone_2_bufchan_buf[0] ? lizzieLet24_3MQNone_2_bufchan_buf :
                                           lizzieLet24_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3MQNone_2_argbuf_r && lizzieLet24_3MQNone_2_bufchan_buf[0]))
        lizzieLet24_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3MQNone_2_argbuf_r) && (! lizzieLet24_3MQNone_2_bufchan_buf[0])))
        lizzieLet24_3MQNone_2_bufchan_buf <= lizzieLet24_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C16,Ty Go) : [(lizzieLet24_3MQNone_2_argbuf,Go),
                            (lizzieLet60_3Lcall_f_f_Int0_1_argbuf,Go),
                            (lizzieLet24_3MQVal_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf,Go),
                            (es_6_1_2MyFalse_2_argbuf,Go),
                            (es_6_1_2MyTrue_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf,Go),
                            (lizzieLet24_5MQNode_4QError_Int_2_argbuf,Go)] > (go_18_goMux_choice,C16) (go_18_goMux_data,Go) */
  logic [15:0] lizzieLet24_3MQNone_2_argbuf_select_d;
  assign lizzieLet24_3MQNone_2_argbuf_select_d = ((| lizzieLet24_3MQNone_2_argbuf_select_q) ? lizzieLet24_3MQNone_2_argbuf_select_q :
                                                  (lizzieLet24_3MQNone_2_argbuf_d[0] ? 16'd1 :
                                                   (lizzieLet60_3Lcall_f_f_Int0_1_argbuf_d[0] ? 16'd2 :
                                                    (lizzieLet24_3MQVal_2_argbuf_d[0] ? 16'd4 :
                                                     (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_d[0] ? 16'd8 :
                                                      (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_d[0] ? 16'd16 :
                                                       (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_d[0] ? 16'd32 :
                                                        (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_d[0] ? 16'd64 :
                                                         (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_d[0] ? 16'd128 :
                                                          (es_6_1_2MyFalse_2_argbuf_d[0] ? 16'd256 :
                                                           (es_6_1_2MyTrue_2_argbuf_d[0] ? 16'd512 :
                                                            (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_d[0] ? 16'd1024 :
                                                             (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_d[0] ? 16'd2048 :
                                                              (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_d[0] ? 16'd4096 :
                                                               (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_d[0] ? 16'd8192 :
                                                                (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_d[0] ? 16'd16384 :
                                                                 (lizzieLet24_5MQNode_4QError_Int_2_argbuf_d[0] ? 16'd32768 :
                                                                  16'd0)))))))))))))))));
  logic [15:0] lizzieLet24_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3MQNone_2_argbuf_select_q <= 16'd0;
    else
      lizzieLet24_3MQNone_2_argbuf_select_q <= (lizzieLet24_3MQNone_2_argbuf_done ? 16'd0 :
                                                lizzieLet24_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet24_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet24_3MQNone_2_argbuf_emit_q <= (lizzieLet24_3MQNone_2_argbuf_done ? 2'd0 :
                                              lizzieLet24_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet24_3MQNone_2_argbuf_emit_d;
  assign lizzieLet24_3MQNone_2_argbuf_emit_d = (lizzieLet24_3MQNone_2_argbuf_emit_q | ({go_18_goMux_choice_d[0],
                                                                                        go_18_goMux_data_d[0]} & {go_18_goMux_choice_r,
                                                                                                                  go_18_goMux_data_r}));
  logic lizzieLet24_3MQNone_2_argbuf_done;
  assign lizzieLet24_3MQNone_2_argbuf_done = (& lizzieLet24_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet24_5MQNode_4QError_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_r,
          es_6_1_2MyTrue_2_argbuf_r,
          es_6_1_2MyFalse_2_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_r,
          lizzieLet24_3MQVal_2_argbuf_r,
          lizzieLet60_3Lcall_f_f_Int0_1_argbuf_r,
          lizzieLet24_3MQNone_2_argbuf_r} = (lizzieLet24_3MQNone_2_argbuf_done ? lizzieLet24_3MQNone_2_argbuf_select_d :
                                             16'd0);
  assign go_18_goMux_data_d = ((lizzieLet24_3MQNone_2_argbuf_select_d[0] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_3MQNone_2_argbuf_d :
                               ((lizzieLet24_3MQNone_2_argbuf_select_d[1] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet60_3Lcall_f_f_Int0_1_argbuf_d :
                                ((lizzieLet24_3MQNone_2_argbuf_select_d[2] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_3MQVal_2_argbuf_d :
                                 ((lizzieLet24_3MQNone_2_argbuf_select_d[3] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_d :
                                  ((lizzieLet24_3MQNone_2_argbuf_select_d[4] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_d :
                                   ((lizzieLet24_3MQNone_2_argbuf_select_d[5] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_d :
                                    ((lizzieLet24_3MQNone_2_argbuf_select_d[6] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_d :
                                     ((lizzieLet24_3MQNone_2_argbuf_select_d[7] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_d :
                                      ((lizzieLet24_3MQNone_2_argbuf_select_d[8] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? es_6_1_2MyFalse_2_argbuf_d :
                                       ((lizzieLet24_3MQNone_2_argbuf_select_d[9] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? es_6_1_2MyTrue_2_argbuf_d :
                                        ((lizzieLet24_3MQNone_2_argbuf_select_d[10] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_d :
                                         ((lizzieLet24_3MQNone_2_argbuf_select_d[11] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_d :
                                          ((lizzieLet24_3MQNone_2_argbuf_select_d[12] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_d :
                                           ((lizzieLet24_3MQNone_2_argbuf_select_d[13] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_d :
                                            ((lizzieLet24_3MQNone_2_argbuf_select_d[14] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_d :
                                             ((lizzieLet24_3MQNone_2_argbuf_select_d[15] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_5MQNode_4QError_Int_2_argbuf_d :
                                              1'd0))))))))))))))));
  assign go_18_goMux_choice_d = ((lizzieLet24_3MQNone_2_argbuf_select_d[0] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C1_16_dc(1'd1) :
                                 ((lizzieLet24_3MQNone_2_argbuf_select_d[1] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C2_16_dc(1'd1) :
                                  ((lizzieLet24_3MQNone_2_argbuf_select_d[2] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C3_16_dc(1'd1) :
                                   ((lizzieLet24_3MQNone_2_argbuf_select_d[3] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C4_16_dc(1'd1) :
                                    ((lizzieLet24_3MQNone_2_argbuf_select_d[4] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C5_16_dc(1'd1) :
                                     ((lizzieLet24_3MQNone_2_argbuf_select_d[5] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C6_16_dc(1'd1) :
                                      ((lizzieLet24_3MQNone_2_argbuf_select_d[6] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C7_16_dc(1'd1) :
                                       ((lizzieLet24_3MQNone_2_argbuf_select_d[7] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C8_16_dc(1'd1) :
                                        ((lizzieLet24_3MQNone_2_argbuf_select_d[8] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C9_16_dc(1'd1) :
                                         ((lizzieLet24_3MQNone_2_argbuf_select_d[9] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C10_16_dc(1'd1) :
                                          ((lizzieLet24_3MQNone_2_argbuf_select_d[10] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C11_16_dc(1'd1) :
                                           ((lizzieLet24_3MQNone_2_argbuf_select_d[11] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C12_16_dc(1'd1) :
                                            ((lizzieLet24_3MQNone_2_argbuf_select_d[12] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C13_16_dc(1'd1) :
                                             ((lizzieLet24_3MQNone_2_argbuf_select_d[13] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C14_16_dc(1'd1) :
                                              ((lizzieLet24_3MQNone_2_argbuf_select_d[14] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C15_16_dc(1'd1) :
                                               ((lizzieLet24_3MQNone_2_argbuf_select_d[15] && (! lizzieLet24_3MQNone_2_argbuf_emit_q[1])) ? C16_16_dc(1'd1) :
                                                {4'd0, 1'd0}))))))))))))))));
  
  /* fork (Ty Go) : (lizzieLet24_3MQVal,Go) > [(lizzieLet24_3MQVal_1,Go),
                                          (lizzieLet24_3MQVal_2,Go)] */
  logic [1:0] lizzieLet24_3MQVal_emitted;
  logic [1:0] lizzieLet24_3MQVal_done;
  assign lizzieLet24_3MQVal_1_d = (lizzieLet24_3MQVal_d[0] && (! lizzieLet24_3MQVal_emitted[0]));
  assign lizzieLet24_3MQVal_2_d = (lizzieLet24_3MQVal_d[0] && (! lizzieLet24_3MQVal_emitted[1]));
  assign lizzieLet24_3MQVal_done = (lizzieLet24_3MQVal_emitted | ({lizzieLet24_3MQVal_2_d[0],
                                                                   lizzieLet24_3MQVal_1_d[0]} & {lizzieLet24_3MQVal_2_r,
                                                                                                 lizzieLet24_3MQVal_1_r}));
  assign lizzieLet24_3MQVal_r = (& lizzieLet24_3MQVal_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQVal_emitted <= 2'd0;
    else
      lizzieLet24_3MQVal_emitted <= (lizzieLet24_3MQVal_r ? 2'd0 :
                                     lizzieLet24_3MQVal_done);
  
  /* buf (Ty Go) : (lizzieLet24_3MQVal_1,Go) > (lizzieLet24_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet24_3MQVal_1_bufchan_d;
  logic lizzieLet24_3MQVal_1_bufchan_r;
  assign lizzieLet24_3MQVal_1_r = ((! lizzieLet24_3MQVal_1_bufchan_d[0]) || lizzieLet24_3MQVal_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQVal_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3MQVal_1_r)
        lizzieLet24_3MQVal_1_bufchan_d <= lizzieLet24_3MQVal_1_d;
  Go_t lizzieLet24_3MQVal_1_bufchan_buf;
  assign lizzieLet24_3MQVal_1_bufchan_r = (! lizzieLet24_3MQVal_1_bufchan_buf[0]);
  assign lizzieLet24_3MQVal_1_argbuf_d = (lizzieLet24_3MQVal_1_bufchan_buf[0] ? lizzieLet24_3MQVal_1_bufchan_buf :
                                          lizzieLet24_3MQVal_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQVal_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3MQVal_1_argbuf_r && lizzieLet24_3MQVal_1_bufchan_buf[0]))
        lizzieLet24_3MQVal_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3MQVal_1_argbuf_r) && (! lizzieLet24_3MQVal_1_bufchan_buf[0])))
        lizzieLet24_3MQVal_1_bufchan_buf <= lizzieLet24_3MQVal_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) : [(lizzieLet24_3MQVal_1_argbuf,Go),
                                                                                              (lizzieLet24_7MQVal_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet24_8MQVal_1_argbuf,Pointer_QTree_Int),
                                                                                              (lizzieLet24_4MQVal_1_argbuf,MyDTInt_Bool),
                                                                                              (lizzieLet24_9MQVal_1_argbuf,MyDTInt_Int_Int)] > (f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int) */
  assign \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_dc((& {lizzieLet24_3MQVal_1_argbuf_d[0],
                                                                                                                                                                                               lizzieLet24_7MQVal_1_argbuf_d[0],
                                                                                                                                                                                               lizzieLet24_8MQVal_1_argbuf_d[0],
                                                                                                                                                                                               lizzieLet24_4MQVal_1_argbuf_d[0],
                                                                                                                                                                                               lizzieLet24_9MQVal_1_argbuf_d[0]}), lizzieLet24_3MQVal_1_argbuf_d, lizzieLet24_7MQVal_1_argbuf_d, lizzieLet24_8MQVal_1_argbuf_d, lizzieLet24_4MQVal_1_argbuf_d, lizzieLet24_9MQVal_1_argbuf_d);
  assign {lizzieLet24_3MQVal_1_argbuf_r,
          lizzieLet24_7MQVal_1_argbuf_r,
          lizzieLet24_8MQVal_1_argbuf_r,
          lizzieLet24_4MQVal_1_argbuf_r,
          lizzieLet24_9MQVal_1_argbuf_r} = {5 {(\f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_r  && \f'_f'_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_3MQVal_2,Go) > (lizzieLet24_3MQVal_2_argbuf,Go) */
  Go_t lizzieLet24_3MQVal_2_bufchan_d;
  logic lizzieLet24_3MQVal_2_bufchan_r;
  assign lizzieLet24_3MQVal_2_r = ((! lizzieLet24_3MQVal_2_bufchan_d[0]) || lizzieLet24_3MQVal_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQVal_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3MQVal_2_r)
        lizzieLet24_3MQVal_2_bufchan_d <= lizzieLet24_3MQVal_2_d;
  Go_t lizzieLet24_3MQVal_2_bufchan_buf;
  assign lizzieLet24_3MQVal_2_bufchan_r = (! lizzieLet24_3MQVal_2_bufchan_buf[0]);
  assign lizzieLet24_3MQVal_2_argbuf_d = (lizzieLet24_3MQVal_2_bufchan_buf[0] ? lizzieLet24_3MQVal_2_bufchan_buf :
                                          lizzieLet24_3MQVal_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_3MQVal_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3MQVal_2_argbuf_r && lizzieLet24_3MQVal_2_bufchan_buf[0]))
        lizzieLet24_3MQVal_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3MQVal_2_argbuf_r) && (! lizzieLet24_3MQVal_2_bufchan_buf[0])))
        lizzieLet24_3MQVal_2_bufchan_buf <= lizzieLet24_3MQVal_2_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty MyDTInt_Bool) : (lizzieLet24_4,MaskQTree) (is_zae6_goMux_mux,MyDTInt_Bool) > [(_108,MyDTInt_Bool),
                                                                                        (lizzieLet24_4MQVal,MyDTInt_Bool),
                                                                                        (lizzieLet24_4MQNode,MyDTInt_Bool)] */
  logic [2:0] is_zae6_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_4_d[0] && is_zae6_goMux_mux_d[0]))
      unique case (lizzieLet24_4_d[2:1])
        2'd0: is_zae6_goMux_mux_onehotd = 3'd1;
        2'd1: is_zae6_goMux_mux_onehotd = 3'd2;
        2'd2: is_zae6_goMux_mux_onehotd = 3'd4;
        default: is_zae6_goMux_mux_onehotd = 3'd0;
      endcase
    else is_zae6_goMux_mux_onehotd = 3'd0;
  assign _108_d = is_zae6_goMux_mux_onehotd[0];
  assign lizzieLet24_4MQVal_d = is_zae6_goMux_mux_onehotd[1];
  assign lizzieLet24_4MQNode_d = is_zae6_goMux_mux_onehotd[2];
  assign is_zae6_goMux_mux_r = (| (is_zae6_goMux_mux_onehotd & {lizzieLet24_4MQNode_r,
                                                                lizzieLet24_4MQVal_r,
                                                                _108_r}));
  assign lizzieLet24_4_r = is_zae6_goMux_mux_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet24_4MQVal,MyDTInt_Bool) > (lizzieLet24_4MQVal_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet24_4MQVal_bufchan_d;
  logic lizzieLet24_4MQVal_bufchan_r;
  assign lizzieLet24_4MQVal_r = ((! lizzieLet24_4MQVal_bufchan_d[0]) || lizzieLet24_4MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_4MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_4MQVal_r)
        lizzieLet24_4MQVal_bufchan_d <= lizzieLet24_4MQVal_d;
  MyDTInt_Bool_t lizzieLet24_4MQVal_bufchan_buf;
  assign lizzieLet24_4MQVal_bufchan_r = (! lizzieLet24_4MQVal_bufchan_buf[0]);
  assign lizzieLet24_4MQVal_1_argbuf_d = (lizzieLet24_4MQVal_bufchan_buf[0] ? lizzieLet24_4MQVal_bufchan_buf :
                                          lizzieLet24_4MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_4MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_4MQVal_1_argbuf_r && lizzieLet24_4MQVal_bufchan_buf[0]))
        lizzieLet24_4MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_4MQVal_1_argbuf_r) && (! lizzieLet24_4MQVal_bufchan_buf[0])))
        lizzieLet24_4MQVal_bufchan_buf <= lizzieLet24_4MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Int) : (lizzieLet24_5,MaskQTree) (readPointer_QTree_Intm2ae4_1_argbuf_rwb,QTree_Int) > [(_107,QTree_Int),
                                                                                                        (_106,QTree_Int),
                                                                                                        (lizzieLet24_5MQNode,QTree_Int)] */
  logic [2:0] readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet24_5_d[0] && readPointer_QTree_Intm2ae4_1_argbuf_rwb_d[0]))
      unique case (lizzieLet24_5_d[2:1])
        2'd0: readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd = 3'd0;
  assign _107_d = {readPointer_QTree_Intm2ae4_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd[0]};
  assign _106_d = {readPointer_QTree_Intm2ae4_1_argbuf_rwb_d[66:1],
                   readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet24_5MQNode_d = {readPointer_QTree_Intm2ae4_1_argbuf_rwb_d[66:1],
                                  readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Intm2ae4_1_argbuf_rwb_r = (| (readPointer_QTree_Intm2ae4_1_argbuf_rwb_onehotd & {lizzieLet24_5MQNode_r,
                                                                                                            _106_r,
                                                                                                            _107_r}));
  assign lizzieLet24_5_r = readPointer_QTree_Intm2ae4_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet24_5MQNode,QTree_Int) > [(lizzieLet24_5MQNode_1,QTree_Int),
                                                         (lizzieLet24_5MQNode_2,QTree_Int),
                                                         (lizzieLet24_5MQNode_3,QTree_Int),
                                                         (lizzieLet24_5MQNode_4,QTree_Int),
                                                         (lizzieLet24_5MQNode_5,QTree_Int),
                                                         (lizzieLet24_5MQNode_6,QTree_Int),
                                                         (lizzieLet24_5MQNode_7,QTree_Int),
                                                         (lizzieLet24_5MQNode_8,QTree_Int),
                                                         (lizzieLet24_5MQNode_9,QTree_Int),
                                                         (lizzieLet24_5MQNode_10,QTree_Int),
                                                         (lizzieLet24_5MQNode_11,QTree_Int)] */
  logic [10:0] lizzieLet24_5MQNode_emitted;
  logic [10:0] lizzieLet24_5MQNode_done;
  assign lizzieLet24_5MQNode_1_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[0]))};
  assign lizzieLet24_5MQNode_2_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[1]))};
  assign lizzieLet24_5MQNode_3_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[2]))};
  assign lizzieLet24_5MQNode_4_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[3]))};
  assign lizzieLet24_5MQNode_5_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[4]))};
  assign lizzieLet24_5MQNode_6_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[5]))};
  assign lizzieLet24_5MQNode_7_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[6]))};
  assign lizzieLet24_5MQNode_8_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[7]))};
  assign lizzieLet24_5MQNode_9_d = {lizzieLet24_5MQNode_d[66:1],
                                    (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[8]))};
  assign lizzieLet24_5MQNode_10_d = {lizzieLet24_5MQNode_d[66:1],
                                     (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[9]))};
  assign lizzieLet24_5MQNode_11_d = {lizzieLet24_5MQNode_d[66:1],
                                     (lizzieLet24_5MQNode_d[0] && (! lizzieLet24_5MQNode_emitted[10]))};
  assign lizzieLet24_5MQNode_done = (lizzieLet24_5MQNode_emitted | ({lizzieLet24_5MQNode_11_d[0],
                                                                     lizzieLet24_5MQNode_10_d[0],
                                                                     lizzieLet24_5MQNode_9_d[0],
                                                                     lizzieLet24_5MQNode_8_d[0],
                                                                     lizzieLet24_5MQNode_7_d[0],
                                                                     lizzieLet24_5MQNode_6_d[0],
                                                                     lizzieLet24_5MQNode_5_d[0],
                                                                     lizzieLet24_5MQNode_4_d[0],
                                                                     lizzieLet24_5MQNode_3_d[0],
                                                                     lizzieLet24_5MQNode_2_d[0],
                                                                     lizzieLet24_5MQNode_1_d[0]} & {lizzieLet24_5MQNode_11_r,
                                                                                                    lizzieLet24_5MQNode_10_r,
                                                                                                    lizzieLet24_5MQNode_9_r,
                                                                                                    lizzieLet24_5MQNode_8_r,
                                                                                                    lizzieLet24_5MQNode_7_r,
                                                                                                    lizzieLet24_5MQNode_6_r,
                                                                                                    lizzieLet24_5MQNode_5_r,
                                                                                                    lizzieLet24_5MQNode_4_r,
                                                                                                    lizzieLet24_5MQNode_3_r,
                                                                                                    lizzieLet24_5MQNode_2_r,
                                                                                                    lizzieLet24_5MQNode_1_r}));
  assign lizzieLet24_5MQNode_r = (& lizzieLet24_5MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_5MQNode_emitted <= 11'd0;
    else
      lizzieLet24_5MQNode_emitted <= (lizzieLet24_5MQNode_r ? 11'd0 :
                                      lizzieLet24_5MQNode_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_10,QTree_Int) (q3aea_destruct,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_10QNone_Int,Pointer_MaskQTree),
                                                                                                        (_105,Pointer_MaskQTree),
                                                                                                        (lizzieLet24_5MQNode_10QNode_Int,Pointer_MaskQTree),
                                                                                                        (_104,Pointer_MaskQTree)] */
  logic [3:0] q3aea_destruct_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_10_d[0] && q3aea_destruct_d[0]))
      unique case (lizzieLet24_5MQNode_10_d[2:1])
        2'd0: q3aea_destruct_onehotd = 4'd1;
        2'd1: q3aea_destruct_onehotd = 4'd2;
        2'd2: q3aea_destruct_onehotd = 4'd4;
        2'd3: q3aea_destruct_onehotd = 4'd8;
        default: q3aea_destruct_onehotd = 4'd0;
      endcase
    else q3aea_destruct_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_10QNone_Int_d = {q3aea_destruct_d[16:1],
                                              q3aea_destruct_onehotd[0]};
  assign _105_d = {q3aea_destruct_d[16:1],
                   q3aea_destruct_onehotd[1]};
  assign lizzieLet24_5MQNode_10QNode_Int_d = {q3aea_destruct_d[16:1],
                                              q3aea_destruct_onehotd[2]};
  assign _104_d = {q3aea_destruct_d[16:1],
                   q3aea_destruct_onehotd[3]};
  assign q3aea_destruct_r = (| (q3aea_destruct_onehotd & {_104_r,
                                                          lizzieLet24_5MQNode_10QNode_Int_r,
                                                          _105_r,
                                                          lizzieLet24_5MQNode_10QNone_Int_r}));
  assign lizzieLet24_5MQNode_10_r = q3aea_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_11,QTree_Int) (q4aeb_destruct,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_11QNone_Int,Pointer_MaskQTree),
                                                                                                        (_103,Pointer_MaskQTree),
                                                                                                        (lizzieLet24_5MQNode_11QNode_Int,Pointer_MaskQTree),
                                                                                                        (_102,Pointer_MaskQTree)] */
  logic [3:0] q4aeb_destruct_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_11_d[0] && q4aeb_destruct_d[0]))
      unique case (lizzieLet24_5MQNode_11_d[2:1])
        2'd0: q4aeb_destruct_onehotd = 4'd1;
        2'd1: q4aeb_destruct_onehotd = 4'd2;
        2'd2: q4aeb_destruct_onehotd = 4'd4;
        2'd3: q4aeb_destruct_onehotd = 4'd8;
        default: q4aeb_destruct_onehotd = 4'd0;
      endcase
    else q4aeb_destruct_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_11QNone_Int_d = {q4aeb_destruct_d[16:1],
                                              q4aeb_destruct_onehotd[0]};
  assign _103_d = {q4aeb_destruct_d[16:1],
                   q4aeb_destruct_onehotd[1]};
  assign lizzieLet24_5MQNode_11QNode_Int_d = {q4aeb_destruct_d[16:1],
                                              q4aeb_destruct_onehotd[2]};
  assign _102_d = {q4aeb_destruct_d[16:1],
                   q4aeb_destruct_onehotd[3]};
  assign q4aeb_destruct_r = (| (q4aeb_destruct_onehotd & {_102_r,
                                                          lizzieLet24_5MQNode_11QNode_Int_r,
                                                          _103_r,
                                                          lizzieLet24_5MQNode_11QNone_Int_r}));
  assign lizzieLet24_5MQNode_11_r = q4aeb_destruct_r;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet24_5MQNode_1QNode_Int,QTree_Int) > [(q1'aen_destruct,Pointer_QTree_Int),
                                                                          (q2'aeo_destruct,Pointer_QTree_Int),
                                                                          (q3'aep_destruct,Pointer_QTree_Int),
                                                                          (q4'aeq_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_1QNode_Int_emitted;
  logic [3:0] lizzieLet24_5MQNode_1QNode_Int_done;
  assign \q1'aen_destruct_d  = {lizzieLet24_5MQNode_1QNode_Int_d[18:3],
                                (lizzieLet24_5MQNode_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_1QNode_Int_emitted[0]))};
  assign \q2'aeo_destruct_d  = {lizzieLet24_5MQNode_1QNode_Int_d[34:19],
                                (lizzieLet24_5MQNode_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_1QNode_Int_emitted[1]))};
  assign \q3'aep_destruct_d  = {lizzieLet24_5MQNode_1QNode_Int_d[50:35],
                                (lizzieLet24_5MQNode_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_1QNode_Int_emitted[2]))};
  assign \q4'aeq_destruct_d  = {lizzieLet24_5MQNode_1QNode_Int_d[66:51],
                                (lizzieLet24_5MQNode_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_1QNode_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_1QNode_Int_done = (lizzieLet24_5MQNode_1QNode_Int_emitted | ({\q4'aeq_destruct_d [0],
                                                                                           \q3'aep_destruct_d [0],
                                                                                           \q2'aeo_destruct_d [0],
                                                                                           \q1'aen_destruct_d [0]} & {\q4'aeq_destruct_r ,
                                                                                                                      \q3'aep_destruct_r ,
                                                                                                                      \q2'aeo_destruct_r ,
                                                                                                                      \q1'aen_destruct_r }));
  assign lizzieLet24_5MQNode_1QNode_Int_r = (& lizzieLet24_5MQNode_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet24_5MQNode_1QNode_Int_emitted <= (lizzieLet24_5MQNode_1QNode_Int_r ? 4'd0 :
                                                 lizzieLet24_5MQNode_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet24_5MQNode_1QVal_Int,QTree_Int) > [(v1aeh_destruct,Int)] */
  assign v1aeh_destruct_d = {lizzieLet24_5MQNode_1QVal_Int_d[34:3],
                             lizzieLet24_5MQNode_1QVal_Int_d[0]};
  assign lizzieLet24_5MQNode_1QVal_Int_r = v1aeh_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet24_5MQNode_2,QTree_Int) (lizzieLet24_5MQNode_1,QTree_Int) > [(_101,QTree_Int),
                                                                                              (lizzieLet24_5MQNode_1QVal_Int,QTree_Int),
                                                                                              (lizzieLet24_5MQNode_1QNode_Int,QTree_Int),
                                                                                              (_100,QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_1_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_2_d[0] && lizzieLet24_5MQNode_1_d[0]))
      unique case (lizzieLet24_5MQNode_2_d[2:1])
        2'd0: lizzieLet24_5MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_1_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_1_onehotd = 4'd0;
  assign _101_d = {lizzieLet24_5MQNode_1_d[66:1],
                   lizzieLet24_5MQNode_1_onehotd[0]};
  assign lizzieLet24_5MQNode_1QVal_Int_d = {lizzieLet24_5MQNode_1_d[66:1],
                                            lizzieLet24_5MQNode_1_onehotd[1]};
  assign lizzieLet24_5MQNode_1QNode_Int_d = {lizzieLet24_5MQNode_1_d[66:1],
                                             lizzieLet24_5MQNode_1_onehotd[2]};
  assign _100_d = {lizzieLet24_5MQNode_1_d[66:1],
                   lizzieLet24_5MQNode_1_onehotd[3]};
  assign lizzieLet24_5MQNode_1_r = (| (lizzieLet24_5MQNode_1_onehotd & {_100_r,
                                                                        lizzieLet24_5MQNode_1QNode_Int_r,
                                                                        lizzieLet24_5MQNode_1QVal_Int_r,
                                                                        _101_r}));
  assign lizzieLet24_5MQNode_2_r = lizzieLet24_5MQNode_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_3,QTree_Int) (lizzieLet24_10MQNode,Pointer_CTf_f_Int) > [(lizzieLet24_5MQNode_3QNone_Int,Pointer_CTf_f_Int),
                                                                                                             (lizzieLet24_5MQNode_3QVal_Int,Pointer_CTf_f_Int),
                                                                                                             (lizzieLet24_5MQNode_3QNode_Int,Pointer_CTf_f_Int),
                                                                                                             (lizzieLet24_5MQNode_3QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet24_10MQNode_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_3_d[0] && lizzieLet24_10MQNode_d[0]))
      unique case (lizzieLet24_5MQNode_3_d[2:1])
        2'd0: lizzieLet24_10MQNode_onehotd = 4'd1;
        2'd1: lizzieLet24_10MQNode_onehotd = 4'd2;
        2'd2: lizzieLet24_10MQNode_onehotd = 4'd4;
        2'd3: lizzieLet24_10MQNode_onehotd = 4'd8;
        default: lizzieLet24_10MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet24_10MQNode_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_3QNone_Int_d = {lizzieLet24_10MQNode_d[16:1],
                                             lizzieLet24_10MQNode_onehotd[0]};
  assign lizzieLet24_5MQNode_3QVal_Int_d = {lizzieLet24_10MQNode_d[16:1],
                                            lizzieLet24_10MQNode_onehotd[1]};
  assign lizzieLet24_5MQNode_3QNode_Int_d = {lizzieLet24_10MQNode_d[16:1],
                                             lizzieLet24_10MQNode_onehotd[2]};
  assign lizzieLet24_5MQNode_3QError_Int_d = {lizzieLet24_10MQNode_d[16:1],
                                              lizzieLet24_10MQNode_onehotd[3]};
  assign lizzieLet24_10MQNode_r = (| (lizzieLet24_10MQNode_onehotd & {lizzieLet24_5MQNode_3QError_Int_r,
                                                                      lizzieLet24_5MQNode_3QNode_Int_r,
                                                                      lizzieLet24_5MQNode_3QVal_Int_r,
                                                                      lizzieLet24_5MQNode_3QNone_Int_r}));
  assign lizzieLet24_5MQNode_3_r = lizzieLet24_10MQNode_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_3QError_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_3QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_3QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_3QError_Int_r = ((! lizzieLet24_5MQNode_3QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_3QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_3QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet24_5MQNode_3QError_Int_r)
        lizzieLet24_5MQNode_3QError_Int_bufchan_d <= lizzieLet24_5MQNode_3QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_3QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_3QError_Int_bufchan_r = (! lizzieLet24_5MQNode_3QError_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_3QError_Int_1_argbuf_d = (lizzieLet24_5MQNode_3QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_3QError_Int_bufchan_buf :
                                                       lizzieLet24_5MQNode_3QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_3QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_5MQNode_3QError_Int_1_argbuf_r && lizzieLet24_5MQNode_3QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_3QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet24_5MQNode_3QError_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_3QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_3QError_Int_bufchan_buf <= lizzieLet24_5MQNode_3QError_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet24_5MQNode_4,QTree_Int) (lizzieLet24_3MQNode,Go) > [(lizzieLet24_5MQNode_4QNone_Int,Go),
                                                                              (lizzieLet24_5MQNode_4QVal_Int,Go),
                                                                              (lizzieLet24_5MQNode_4QNode_Int,Go),
                                                                              (lizzieLet24_5MQNode_4QError_Int,Go)] */
  logic [3:0] lizzieLet24_3MQNode_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_4_d[0] && lizzieLet24_3MQNode_d[0]))
      unique case (lizzieLet24_5MQNode_4_d[2:1])
        2'd0: lizzieLet24_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet24_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet24_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet24_3MQNode_onehotd = 4'd8;
        default: lizzieLet24_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet24_3MQNode_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_4QNone_Int_d = lizzieLet24_3MQNode_onehotd[0];
  assign lizzieLet24_5MQNode_4QVal_Int_d = lizzieLet24_3MQNode_onehotd[1];
  assign lizzieLet24_5MQNode_4QNode_Int_d = lizzieLet24_3MQNode_onehotd[2];
  assign lizzieLet24_5MQNode_4QError_Int_d = lizzieLet24_3MQNode_onehotd[3];
  assign lizzieLet24_3MQNode_r = (| (lizzieLet24_3MQNode_onehotd & {lizzieLet24_5MQNode_4QError_Int_r,
                                                                    lizzieLet24_5MQNode_4QNode_Int_r,
                                                                    lizzieLet24_5MQNode_4QVal_Int_r,
                                                                    lizzieLet24_5MQNode_4QNone_Int_r}));
  assign lizzieLet24_5MQNode_4_r = lizzieLet24_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_4QError_Int,Go) > [(lizzieLet24_5MQNode_4QError_Int_1,Go),
                                                       (lizzieLet24_5MQNode_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_4QError_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_4QError_Int_done;
  assign lizzieLet24_5MQNode_4QError_Int_1_d = (lizzieLet24_5MQNode_4QError_Int_d[0] && (! lizzieLet24_5MQNode_4QError_Int_emitted[0]));
  assign lizzieLet24_5MQNode_4QError_Int_2_d = (lizzieLet24_5MQNode_4QError_Int_d[0] && (! lizzieLet24_5MQNode_4QError_Int_emitted[1]));
  assign lizzieLet24_5MQNode_4QError_Int_done = (lizzieLet24_5MQNode_4QError_Int_emitted | ({lizzieLet24_5MQNode_4QError_Int_2_d[0],
                                                                                             lizzieLet24_5MQNode_4QError_Int_1_d[0]} & {lizzieLet24_5MQNode_4QError_Int_2_r,
                                                                                                                                        lizzieLet24_5MQNode_4QError_Int_1_r}));
  assign lizzieLet24_5MQNode_4QError_Int_r = (& lizzieLet24_5MQNode_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_4QError_Int_emitted <= (lizzieLet24_5MQNode_4QError_Int_r ? 2'd0 :
                                                  lizzieLet24_5MQNode_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_4QError_Int_1,Go)] > (lizzieLet24_5MQNode_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_4QError_Int_1_d[0]}), lizzieLet24_5MQNode_4QError_Int_1_d);
  assign {lizzieLet24_5MQNode_4QError_Int_1_r} = {1 {(lizzieLet24_5MQNode_4QError_Int_1QError_Int_r && lizzieLet24_5MQNode_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet42_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_4QError_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet24_5MQNode_4QError_Int_1QError_Int_r)
        lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet42_1_argbuf_d = (lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet42_1_argbuf_r && lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet42_1_argbuf_r) && (! lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_4QError_Int_2,Go) > (lizzieLet24_5MQNode_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_4QError_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_4QError_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_4QError_Int_2_r = ((! lizzieLet24_5MQNode_4QError_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_4QError_Int_2_r)
        lizzieLet24_5MQNode_4QError_Int_2_bufchan_d <= lizzieLet24_5MQNode_4QError_Int_2_d;
  Go_t lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_4QError_Int_2_bufchan_r = (! lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_4QError_Int_2_argbuf_d = (lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf :
                                                       lizzieLet24_5MQNode_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_4QError_Int_2_argbuf_r && lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_4QError_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_4QError_Int_2_bufchan_buf <= lizzieLet24_5MQNode_4QError_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_5,QTree_Int) (lizzieLet24_4MQNode,MyDTInt_Bool) > [(_99,MyDTInt_Bool),
                                                                                                  (lizzieLet24_5MQNode_5QVal_Int,MyDTInt_Bool),
                                                                                                  (lizzieLet24_5MQNode_5QNode_Int,MyDTInt_Bool),
                                                                                                  (_98,MyDTInt_Bool)] */
  logic [3:0] lizzieLet24_4MQNode_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_5_d[0] && lizzieLet24_4MQNode_d[0]))
      unique case (lizzieLet24_5MQNode_5_d[2:1])
        2'd0: lizzieLet24_4MQNode_onehotd = 4'd1;
        2'd1: lizzieLet24_4MQNode_onehotd = 4'd2;
        2'd2: lizzieLet24_4MQNode_onehotd = 4'd4;
        2'd3: lizzieLet24_4MQNode_onehotd = 4'd8;
        default: lizzieLet24_4MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet24_4MQNode_onehotd = 4'd0;
  assign _99_d = lizzieLet24_4MQNode_onehotd[0];
  assign lizzieLet24_5MQNode_5QVal_Int_d = lizzieLet24_4MQNode_onehotd[1];
  assign lizzieLet24_5MQNode_5QNode_Int_d = lizzieLet24_4MQNode_onehotd[2];
  assign _98_d = lizzieLet24_4MQNode_onehotd[3];
  assign lizzieLet24_4MQNode_r = (| (lizzieLet24_4MQNode_onehotd & {_98_r,
                                                                    lizzieLet24_5MQNode_5QNode_Int_r,
                                                                    lizzieLet24_5MQNode_5QVal_Int_r,
                                                                    _99_r}));
  assign lizzieLet24_5MQNode_5_r = lizzieLet24_4MQNode_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet24_5MQNode_6,QTree_Int) (lizzieLet24_6MQNode,QTree_Int) > [(lizzieLet24_5MQNode_6QNone_Int,QTree_Int),
                                                                                            (lizzieLet24_5MQNode_6QVal_Int,QTree_Int),
                                                                                            (lizzieLet24_5MQNode_6QNode_Int,QTree_Int),
                                                                                            (_97,QTree_Int)] */
  logic [3:0] lizzieLet24_6MQNode_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6_d[0] && lizzieLet24_6MQNode_d[0]))
      unique case (lizzieLet24_5MQNode_6_d[2:1])
        2'd0: lizzieLet24_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet24_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet24_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet24_6MQNode_onehotd = 4'd8;
        default: lizzieLet24_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet24_6MQNode_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNone_Int_d = {lizzieLet24_6MQNode_d[66:1],
                                             lizzieLet24_6MQNode_onehotd[0]};
  assign lizzieLet24_5MQNode_6QVal_Int_d = {lizzieLet24_6MQNode_d[66:1],
                                            lizzieLet24_6MQNode_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_d = {lizzieLet24_6MQNode_d[66:1],
                                             lizzieLet24_6MQNode_onehotd[2]};
  assign _97_d = {lizzieLet24_6MQNode_d[66:1],
                  lizzieLet24_6MQNode_onehotd[3]};
  assign lizzieLet24_6MQNode_r = (| (lizzieLet24_6MQNode_onehotd & {_97_r,
                                                                    lizzieLet24_5MQNode_6QNode_Int_r,
                                                                    lizzieLet24_5MQNode_6QVal_Int_r,
                                                                    lizzieLet24_5MQNode_6QNone_Int_r}));
  assign lizzieLet24_5MQNode_6_r = lizzieLet24_6MQNode_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int,QTree_Int) > [(lizzieLet24_5MQNode_6QNode_Int_1,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_2,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_3,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_4,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_5,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_6,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_7,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_8,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_9,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_10,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_11,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_12,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_13,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNode_Int_14,QTree_Int)] */
  logic [13:0] lizzieLet24_5MQNode_6QNode_Int_emitted;
  logic [13:0] lizzieLet24_5MQNode_6QNode_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_1_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[0]))};
  assign lizzieLet24_5MQNode_6QNode_Int_2_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[1]))};
  assign lizzieLet24_5MQNode_6QNode_Int_3_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[2]))};
  assign lizzieLet24_5MQNode_6QNode_Int_4_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_6QNode_Int_5_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[4]))};
  assign lizzieLet24_5MQNode_6QNode_Int_6_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[5]))};
  assign lizzieLet24_5MQNode_6QNode_Int_7_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[6]))};
  assign lizzieLet24_5MQNode_6QNode_Int_8_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[7]))};
  assign lizzieLet24_5MQNode_6QNode_Int_9_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[8]))};
  assign lizzieLet24_5MQNode_6QNode_Int_10_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                                (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[9]))};
  assign lizzieLet24_5MQNode_6QNode_Int_11_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                                (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[10]))};
  assign lizzieLet24_5MQNode_6QNode_Int_12_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                                (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[11]))};
  assign lizzieLet24_5MQNode_6QNode_Int_13_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                                (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[12]))};
  assign lizzieLet24_5MQNode_6QNode_Int_14_d = {lizzieLet24_5MQNode_6QNode_Int_d[66:1],
                                                (lizzieLet24_5MQNode_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_emitted[13]))};
  assign lizzieLet24_5MQNode_6QNode_Int_done = (lizzieLet24_5MQNode_6QNode_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_14_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_13_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_12_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_11_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_10_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_9_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_8_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_7_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_6_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_5_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_4_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_3_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_2_d[0],
                                                                                           lizzieLet24_5MQNode_6QNode_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_14_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_13_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_12_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_11_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_10_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_9_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_8_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_7_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_6_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_5_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_4_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_3_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_2_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNode_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_emitted <= 14'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_r ? 14'd0 :
                                                 lizzieLet24_5MQNode_6QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_10,QTree_Int) (lizzieLet24_5MQNode_9QNode_Int,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_6QNode_Int_10QNone_Int,Pointer_MaskQTree),
                                                                                                                                   (_96,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet24_5MQNode_6QNode_Int_10QNode_Int,Pointer_MaskQTree),
                                                                                                                                   (_95,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_9QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_10_d[0] && lizzieLet24_5MQNode_9QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_10_d[2:1])
        2'd0: lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_9QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_d = {lizzieLet24_5MQNode_9QNode_Int_d[16:1],
                                                         lizzieLet24_5MQNode_9QNode_Int_onehotd[0]};
  assign _96_d = {lizzieLet24_5MQNode_9QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_9QNode_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_d = {lizzieLet24_5MQNode_9QNode_Int_d[16:1],
                                                         lizzieLet24_5MQNode_9QNode_Int_onehotd[2]};
  assign _95_d = {lizzieLet24_5MQNode_9QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_9QNode_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_9QNode_Int_r = (| (lizzieLet24_5MQNode_9QNode_Int_onehotd & {_95_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_r,
                                                                                          _96_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_10_r = lizzieLet24_5MQNode_9QNode_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_10QNone_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_11,QTree_Int) (q1'aen_destruct,Pointer_QTree_Int) > [(lizzieLet24_5MQNode_6QNode_Int_11QNone_Int,Pointer_QTree_Int),
                                                                                                                    (_94,Pointer_QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_11QNode_Int,Pointer_QTree_Int),
                                                                                                                    (_93,Pointer_QTree_Int)] */
  logic [3:0] \q1'aen_destruct_onehotd ;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_11_d[0] && \q1'aen_destruct_d [0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_11_d[2:1])
        2'd0: \q1'aen_destruct_onehotd  = 4'd1;
        2'd1: \q1'aen_destruct_onehotd  = 4'd2;
        2'd2: \q1'aen_destruct_onehotd  = 4'd4;
        2'd3: \q1'aen_destruct_onehotd  = 4'd8;
        default: \q1'aen_destruct_onehotd  = 4'd0;
      endcase
    else \q1'aen_destruct_onehotd  = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_d = {\q1'aen_destruct_d [16:1],
                                                         \q1'aen_destruct_onehotd [0]};
  assign _94_d = {\q1'aen_destruct_d [16:1],
                  \q1'aen_destruct_onehotd [1]};
  assign lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_d = {\q1'aen_destruct_d [16:1],
                                                         \q1'aen_destruct_onehotd [2]};
  assign _93_d = {\q1'aen_destruct_d [16:1],
                  \q1'aen_destruct_onehotd [3]};
  assign \q1'aen_destruct_r  = (| (\q1'aen_destruct_onehotd  & {_93_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_r,
                                                                _94_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_11_r = \q1'aen_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_11QNone_Int,Pointer_QTree_Int) > (lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_12,QTree_Int) (q2'aeo_destruct,Pointer_QTree_Int) > [(lizzieLet24_5MQNode_6QNode_Int_12QNone_Int,Pointer_QTree_Int),
                                                                                                                    (_92,Pointer_QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_12QNode_Int,Pointer_QTree_Int),
                                                                                                                    (_91,Pointer_QTree_Int)] */
  logic [3:0] \q2'aeo_destruct_onehotd ;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_12_d[0] && \q2'aeo_destruct_d [0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_12_d[2:1])
        2'd0: \q2'aeo_destruct_onehotd  = 4'd1;
        2'd1: \q2'aeo_destruct_onehotd  = 4'd2;
        2'd2: \q2'aeo_destruct_onehotd  = 4'd4;
        2'd3: \q2'aeo_destruct_onehotd  = 4'd8;
        default: \q2'aeo_destruct_onehotd  = 4'd0;
      endcase
    else \q2'aeo_destruct_onehotd  = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_d = {\q2'aeo_destruct_d [16:1],
                                                         \q2'aeo_destruct_onehotd [0]};
  assign _92_d = {\q2'aeo_destruct_d [16:1],
                  \q2'aeo_destruct_onehotd [1]};
  assign lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_d = {\q2'aeo_destruct_d [16:1],
                                                         \q2'aeo_destruct_onehotd [2]};
  assign _91_d = {\q2'aeo_destruct_d [16:1],
                  \q2'aeo_destruct_onehotd [3]};
  assign \q2'aeo_destruct_r  = (| (\q2'aeo_destruct_onehotd  & {_91_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_r,
                                                                _92_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_12_r = \q2'aeo_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_12QNone_Int,Pointer_QTree_Int) > (lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_13,QTree_Int) (q3'aep_destruct,Pointer_QTree_Int) > [(lizzieLet24_5MQNode_6QNode_Int_13QNone_Int,Pointer_QTree_Int),
                                                                                                                    (_90,Pointer_QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_13QNode_Int,Pointer_QTree_Int),
                                                                                                                    (_89,Pointer_QTree_Int)] */
  logic [3:0] \q3'aep_destruct_onehotd ;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_13_d[0] && \q3'aep_destruct_d [0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_13_d[2:1])
        2'd0: \q3'aep_destruct_onehotd  = 4'd1;
        2'd1: \q3'aep_destruct_onehotd  = 4'd2;
        2'd2: \q3'aep_destruct_onehotd  = 4'd4;
        2'd3: \q3'aep_destruct_onehotd  = 4'd8;
        default: \q3'aep_destruct_onehotd  = 4'd0;
      endcase
    else \q3'aep_destruct_onehotd  = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_d = {\q3'aep_destruct_d [16:1],
                                                         \q3'aep_destruct_onehotd [0]};
  assign _90_d = {\q3'aep_destruct_d [16:1],
                  \q3'aep_destruct_onehotd [1]};
  assign lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_d = {\q3'aep_destruct_d [16:1],
                                                         \q3'aep_destruct_onehotd [2]};
  assign _89_d = {\q3'aep_destruct_d [16:1],
                  \q3'aep_destruct_onehotd [3]};
  assign \q3'aep_destruct_r  = (| (\q3'aep_destruct_onehotd  & {_89_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_r,
                                                                _90_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_13_r = \q3'aep_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_13QNone_Int,Pointer_QTree_Int) > (lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_14,QTree_Int) (q4'aeq_destruct,Pointer_QTree_Int) > [(lizzieLet24_5MQNode_6QNode_Int_14QNone_Int,Pointer_QTree_Int),
                                                                                                                    (_88,Pointer_QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int,Pointer_QTree_Int),
                                                                                                                    (_87,Pointer_QTree_Int)] */
  logic [3:0] \q4'aeq_destruct_onehotd ;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_14_d[0] && \q4'aeq_destruct_d [0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_14_d[2:1])
        2'd0: \q4'aeq_destruct_onehotd  = 4'd1;
        2'd1: \q4'aeq_destruct_onehotd  = 4'd2;
        2'd2: \q4'aeq_destruct_onehotd  = 4'd4;
        2'd3: \q4'aeq_destruct_onehotd  = 4'd8;
        default: \q4'aeq_destruct_onehotd  = 4'd0;
      endcase
    else \q4'aeq_destruct_onehotd  = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_d = {\q4'aeq_destruct_d [16:1],
                                                         \q4'aeq_destruct_onehotd [0]};
  assign _88_d = {\q4'aeq_destruct_d [16:1],
                  \q4'aeq_destruct_onehotd [1]};
  assign lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_d = {\q4'aeq_destruct_d [16:1],
                                                         \q4'aeq_destruct_onehotd [2]};
  assign _87_d = {\q4'aeq_destruct_d [16:1],
                  \q4'aeq_destruct_onehotd [3]};
  assign \q4'aeq_destruct_r  = (| (\q4'aeq_destruct_onehotd  & {_87_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_r,
                                                                _88_r,
                                                                lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_14_r = \q4'aeq_destruct_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int,Pointer_QTree_Int) > (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_14QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_14QNone_Int,Pointer_QTree_Int) > (lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int,QTree_Int) > [(t1aes_destruct,Pointer_QTree_Int),
                                                                                     (t2aet_destruct,Pointer_QTree_Int),
                                                                                     (t3aeu_destruct,Pointer_QTree_Int),
                                                                                     (t4aev_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_done;
  assign t1aes_destruct_d = {lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted[0]))};
  assign t2aet_destruct_d = {lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted[1]))};
  assign t3aeu_destruct_d = {lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted[2]))};
  assign t4aev_destruct_d = {lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_done = (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted | ({t4aev_destruct_d[0],
                                                                                                                 t3aeu_destruct_d[0],
                                                                                                                 t2aet_destruct_d[0],
                                                                                                                 t1aes_destruct_d[0]} & {t4aev_destruct_r,
                                                                                                                                         t3aeu_destruct_r,
                                                                                                                                         t2aet_destruct_r,
                                                                                                                                         t1aes_destruct_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_r ? 4'd0 :
                                                            lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_2,QTree_Int) (lizzieLet24_5MQNode_6QNode_Int_1,QTree_Int) > [(_86,QTree_Int),
                                                                                                                    (_85,QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_1QNode_Int,QTree_Int),
                                                                                                                    (_84,QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_6QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_2_d[0] && lizzieLet24_5MQNode_6QNode_Int_1_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_2_d[2:1])
        2'd0: lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_6QNode_Int_1_onehotd = 4'd0;
  assign _86_d = {lizzieLet24_5MQNode_6QNode_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNode_Int_1_onehotd[0]};
  assign _85_d = {lizzieLet24_5MQNode_6QNode_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNode_Int_1_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_d = {lizzieLet24_5MQNode_6QNode_Int_1_d[66:1],
                                                        lizzieLet24_5MQNode_6QNode_Int_1_onehotd[2]};
  assign _84_d = {lizzieLet24_5MQNode_6QNode_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNode_Int_1_onehotd[3]};
  assign lizzieLet24_5MQNode_6QNode_Int_1_r = (| (lizzieLet24_5MQNode_6QNode_Int_1_onehotd & {_84_r,
                                                                                              lizzieLet24_5MQNode_6QNode_Int_1QNode_Int_r,
                                                                                              _85_r,
                                                                                              _86_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_2_r = lizzieLet24_5MQNode_6QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_3,QTree_Int) (lizzieLet24_5MQNode_10QNode_Int,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_6QNode_Int_3QNone_Int,Pointer_MaskQTree),
                                                                                                                                   (_83,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet24_5MQNode_6QNode_Int_3QNode_Int,Pointer_MaskQTree),
                                                                                                                                   (_82,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_10QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_3_d[0] && lizzieLet24_5MQNode_10QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_3_d[2:1])
        2'd0: lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_10QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_d = {lizzieLet24_5MQNode_10QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_10QNode_Int_onehotd[0]};
  assign _83_d = {lizzieLet24_5MQNode_10QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_10QNode_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_d = {lizzieLet24_5MQNode_10QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_10QNode_Int_onehotd[2]};
  assign _82_d = {lizzieLet24_5MQNode_10QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_10QNode_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_10QNode_Int_r = (| (lizzieLet24_5MQNode_10QNode_Int_onehotd & {_82_r,
                                                                                            lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_r,
                                                                                            _83_r,
                                                                                            lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_3_r = lizzieLet24_5MQNode_10QNode_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_3QNone_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_4,QTree_Int) (lizzieLet24_5MQNode_11QNode_Int,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_6QNode_Int_4QNone_Int,Pointer_MaskQTree),
                                                                                                                                   (_81,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int,Pointer_MaskQTree),
                                                                                                                                   (_80,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_11QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_4_d[0] && lizzieLet24_5MQNode_11QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_4_d[2:1])
        2'd0: lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_11QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_d = {lizzieLet24_5MQNode_11QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_11QNode_Int_onehotd[0]};
  assign _81_d = {lizzieLet24_5MQNode_11QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_11QNode_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_d = {lizzieLet24_5MQNode_11QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_11QNode_Int_onehotd[2]};
  assign _80_d = {lizzieLet24_5MQNode_11QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_11QNode_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_11QNode_Int_r = (| (lizzieLet24_5MQNode_11QNode_Int_onehotd & {_80_r,
                                                                                            lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_r,
                                                                                            _81_r,
                                                                                            lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_4_r = lizzieLet24_5MQNode_11QNode_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_4QNone_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNode_Int_5,QTree_Int) (lizzieLet24_5MQNode_3QNode_Int,Pointer_CTf_f_Int) > [(lizzieLet24_5MQNode_6QNode_Int_5QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNode_Int_5QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNode_Int_5QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet24_5MQNode_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_5_d[0] && lizzieLet24_5MQNode_3QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_5_d[2:1])
        2'd0: lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_d = {lizzieLet24_5MQNode_3QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_3QNode_Int_onehotd[0]};
  assign lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_d = {lizzieLet24_5MQNode_3QNode_Int_d[16:1],
                                                       lizzieLet24_5MQNode_3QNode_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_d = {lizzieLet24_5MQNode_3QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_3QNode_Int_onehotd[2]};
  assign lizzieLet24_5MQNode_6QNode_Int_5QError_Int_d = {lizzieLet24_5MQNode_3QNode_Int_d[16:1],
                                                         lizzieLet24_5MQNode_3QNode_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_3QNode_Int_r = (| (lizzieLet24_5MQNode_3QNode_Int_onehotd & {lizzieLet24_5MQNode_6QNode_Int_5QError_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_5_r = lizzieLet24_5MQNode_3QNode_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNode_Int_5QError_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_5QError_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_5QError_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_5QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_5QError_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_5QError_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int3) : [(lizzieLet24_5MQNode_6QNode_Int_5QNode_Int,Pointer_CTf_f_Int),
                              (lizzieLet24_5MQNode_6QNode_Int_9QNode_Int,Pointer_MaskQTree),
                              (lizzieLet24_5MQNode_6QNode_Int_11QNode_Int,Pointer_QTree_Int),
                              (t1aes_destruct,Pointer_QTree_Int),
                              (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1,MyDTInt_Bool),
                              (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1,MyDTInt_Int_Int),
                              (lizzieLet24_5MQNode_6QNode_Int_10QNode_Int,Pointer_MaskQTree),
                              (lizzieLet24_5MQNode_6QNode_Int_12QNode_Int,Pointer_QTree_Int),
                              (t2aet_destruct,Pointer_QTree_Int),
                              (lizzieLet24_5MQNode_6QNode_Int_3QNode_Int,Pointer_MaskQTree),
                              (lizzieLet24_5MQNode_6QNode_Int_13QNode_Int,Pointer_QTree_Int),
                              (t3aeu_destruct,Pointer_QTree_Int)] > (lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3,CTf_f_Int) */
  assign lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_d = Lcall_f_f_Int3_dc((& {lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t1aes_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t2aet_destruct_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_d[0],
                                                                                                                                                                                                                                                                                                                                                                                                                                                                              t3aeu_destruct_d[0]}), lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_d, lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_d, lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_d, t1aes_destruct_d, lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_d, lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_d, lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_d, lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_d, t2aet_destruct_d, lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_d, lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_d, t3aeu_destruct_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_r,
          lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_r,
          lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_r,
          t1aes_destruct_r,
          lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_r,
          lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_r,
          lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_r,
          lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_r,
          t2aet_destruct_r,
          lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_r,
          lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_r,
          t3aeu_destruct_r} = {12 {(lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_r && lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_d[0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3,CTf_f_Int) > (lizzieLet40_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_r = ((! lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_r)
        lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_d;
  CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf[0]);
  assign lizzieLet40_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf :
                                   lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                 1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf <= {163'd0,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                   1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_5QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_11QNode_Int_1t1aes_1lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_10QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_12QNode_Int_1t2aet_1lizzieLet24_5MQNode_6QNode_Int_3QNode_Int_1lizzieLet24_5MQNode_6QNode_Int_13QNode_Int_1t3aeu_1Lcall_f_f_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNode_Int_5QNone_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_5QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6,QTree_Int) (lizzieLet24_5MQNode_4QNode_Int,Go) > [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNode_Int_6QError_Int,Go)] */
  logic [3:0] lizzieLet24_5MQNode_4QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_6_d[0] && lizzieLet24_5MQNode_4QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_6_d[2:1])
        2'd0: lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_4QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d = lizzieLet24_5MQNode_4QNode_Int_onehotd[0];
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_d = lizzieLet24_5MQNode_4QNode_Int_onehotd[1];
  assign lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_d = lizzieLet24_5MQNode_4QNode_Int_onehotd[2];
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_d = lizzieLet24_5MQNode_4QNode_Int_onehotd[3];
  assign lizzieLet24_5MQNode_4QNode_Int_r = (| (lizzieLet24_5MQNode_4QNode_Int_onehotd & {lizzieLet24_5MQNode_6QNode_Int_6QError_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_6_r = lizzieLet24_5MQNode_4QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QError_Int,Go) > [(lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1,Go),
                                                                  (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_6QError_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_d = (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_d = (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_done = (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_d[0],
                                                                                                                   lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_r,
                                                                                                                                                                         lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_6QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_r ? 2'd0 :
                                                             lizzieLet24_5MQNode_6QNode_Int_6QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1,Go)] > (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_r && lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int,QTree_Int) > (lizzieLet41_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet41_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet41_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet41_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_r)
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int,Go) > [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1,Go),
                                                                 (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2,Go),
                                                                 (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3,Go),
                                                                 (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4,Go),
                                                                 (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5,Go)] */
  logic [4:0] lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted;
  logic [4:0] lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted[2]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted[3]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted[4]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_done = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted <= 5'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_r ? 5'd0 :
                                                            lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf,Pointer_MaskQTree),
                                                             (lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_14QNone_Int_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int5_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf,Pointer_MaskQTree),
                                                             (lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_13QNone_Int_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int6_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf,Pointer_MaskQTree),
                                                             (lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_3_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_10QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_12QNone_Int_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int7_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf,Pointer_MaskQTree),
                                                             (lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_4_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNode_Int_11QNone_Int_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int8_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_r)
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QNone_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int,Go) > [(lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1,Go),
                                                                (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_d = (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_d = (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_done = (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_d[0],
                                                                                                               lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_r,
                                                                                                                                                                   lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_r ? 2'd0 :
                                                           lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1,Go)] > (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_d[0]}), lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_d);
  assign {lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_r && lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int,QTree_Int) > (lizzieLet39_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                         1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                           1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2,Go) > (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_r = ((! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_r)
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_6QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_6QNode_Int_7,QTree_Int) (lizzieLet24_5MQNode_5QNode_Int,MyDTInt_Bool) > [(_79,MyDTInt_Bool),
                                                                                                                        (_78,MyDTInt_Bool),
                                                                                                                        (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int,MyDTInt_Bool),
                                                                                                                        (_77,MyDTInt_Bool)] */
  logic [3:0] lizzieLet24_5MQNode_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_7_d[0] && lizzieLet24_5MQNode_5QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_7_d[2:1])
        2'd0: lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_5QNode_Int_onehotd = 4'd0;
  assign _79_d = lizzieLet24_5MQNode_5QNode_Int_onehotd[0];
  assign _78_d = lizzieLet24_5MQNode_5QNode_Int_onehotd[1];
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_d = lizzieLet24_5MQNode_5QNode_Int_onehotd[2];
  assign _77_d = lizzieLet24_5MQNode_5QNode_Int_onehotd[3];
  assign lizzieLet24_5MQNode_5QNode_Int_r = (| (lizzieLet24_5MQNode_5QNode_Int_onehotd & {_77_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_r,
                                                                                          _78_r,
                                                                                          _79_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_7_r = lizzieLet24_5MQNode_5QNode_Int_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int,MyDTInt_Bool) > [(lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1,MyDTInt_Bool),
                                                                                     (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_d = (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_d = (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_done = (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_r ? 2'd0 :
                                                            lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2,MyDTInt_Bool) > (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_r = ((! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_r)
        lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_7QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_6QNode_Int_8,QTree_Int) (lizzieLet24_5MQNode_7QNode_Int,MyDTInt_Int_Int) > [(_76,MyDTInt_Int_Int),
                                                                                                                              (_75,MyDTInt_Int_Int),
                                                                                                                              (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int,MyDTInt_Int_Int),
                                                                                                                              (_74,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet24_5MQNode_7QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_8_d[0] && lizzieLet24_5MQNode_7QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_8_d[2:1])
        2'd0: lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_7QNode_Int_onehotd = 4'd0;
  assign _76_d = lizzieLet24_5MQNode_7QNode_Int_onehotd[0];
  assign _75_d = lizzieLet24_5MQNode_7QNode_Int_onehotd[1];
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_d = lizzieLet24_5MQNode_7QNode_Int_onehotd[2];
  assign _74_d = lizzieLet24_5MQNode_7QNode_Int_onehotd[3];
  assign lizzieLet24_5MQNode_7QNode_Int_r = (| (lizzieLet24_5MQNode_7QNode_Int_onehotd & {_74_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_r,
                                                                                          _75_r,
                                                                                          _76_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_8_r = lizzieLet24_5MQNode_7QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int,MyDTInt_Int_Int) > [(lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1,MyDTInt_Int_Int),
                                                                                           (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_done;
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_d = (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_d = (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_done = (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted | ({lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_r = (& lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_r ? 2'd0 :
                                                            lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_r = ((! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_r)
        lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_8QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_9,QTree_Int) (lizzieLet24_5MQNode_8QNode_Int,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_6QNode_Int_9QNone_Int,Pointer_MaskQTree),
                                                                                                                                  (_73,Pointer_MaskQTree),
                                                                                                                                  (lizzieLet24_5MQNode_6QNode_Int_9QNode_Int,Pointer_MaskQTree),
                                                                                                                                  (_72,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNode_Int_9_d[0] && lizzieLet24_5MQNode_8QNode_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNode_Int_9_d[2:1])
        2'd0: lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_8QNode_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_d = {lizzieLet24_5MQNode_8QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_8QNode_Int_onehotd[0]};
  assign _73_d = {lizzieLet24_5MQNode_8QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_8QNode_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_d = {lizzieLet24_5MQNode_8QNode_Int_d[16:1],
                                                        lizzieLet24_5MQNode_8QNode_Int_onehotd[2]};
  assign _72_d = {lizzieLet24_5MQNode_8QNode_Int_d[16:1],
                  lizzieLet24_5MQNode_8QNode_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_8QNode_Int_r = (| (lizzieLet24_5MQNode_8QNode_Int_onehotd & {_72_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_9QNode_Int_r,
                                                                                          _73_r,
                                                                                          lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNode_Int_9_r = lizzieLet24_5MQNode_8QNode_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNode_Int_9QNone_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_r = ((! lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_r)
        lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNode_Int_9QNone_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNone_Int,QTree_Int) > [(lizzieLet24_5MQNode_6QNone_Int_1,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_2,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_3,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_4,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_5,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_6,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_7,QTree_Int),
                                                                    (lizzieLet24_5MQNode_6QNone_Int_8,QTree_Int)] */
  logic [7:0] lizzieLet24_5MQNode_6QNone_Int_emitted;
  logic [7:0] lizzieLet24_5MQNode_6QNone_Int_done;
  assign lizzieLet24_5MQNode_6QNone_Int_1_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[0]))};
  assign lizzieLet24_5MQNode_6QNone_Int_2_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[1]))};
  assign lizzieLet24_5MQNode_6QNone_Int_3_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[2]))};
  assign lizzieLet24_5MQNode_6QNone_Int_4_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_6QNone_Int_5_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[4]))};
  assign lizzieLet24_5MQNode_6QNone_Int_6_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[5]))};
  assign lizzieLet24_5MQNode_6QNone_Int_7_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[6]))};
  assign lizzieLet24_5MQNode_6QNone_Int_8_d = {lizzieLet24_5MQNode_6QNone_Int_d[66:1],
                                               (lizzieLet24_5MQNode_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_emitted[7]))};
  assign lizzieLet24_5MQNode_6QNone_Int_done = (lizzieLet24_5MQNode_6QNone_Int_emitted | ({lizzieLet24_5MQNode_6QNone_Int_8_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_7_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_6_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_5_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_4_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_3_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_2_d[0],
                                                                                           lizzieLet24_5MQNode_6QNone_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNone_Int_8_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_7_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_6_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_5_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_4_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_3_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_2_r,
                                                                                                                                     lizzieLet24_5MQNode_6QNone_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_emitted <= 8'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_r ? 8'd0 :
                                                 lizzieLet24_5MQNode_6QNone_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int,QTree_Int) > [(t1aed_destruct,Pointer_QTree_Int),
                                                                                     (t2aee_destruct,Pointer_QTree_Int),
                                                                                     (t3aef_destruct,Pointer_QTree_Int),
                                                                                     (t4aeg_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_done;
  assign t1aed_destruct_d = {lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[18:3],
                             (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted[0]))};
  assign t2aee_destruct_d = {lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[34:19],
                             (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted[1]))};
  assign t3aef_destruct_d = {lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[50:35],
                             (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted[2]))};
  assign t4aeg_destruct_d = {lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[66:51],
                             (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_done = (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted | ({t4aeg_destruct_d[0],
                                                                                                                 t3aef_destruct_d[0],
                                                                                                                 t2aee_destruct_d[0],
                                                                                                                 t1aed_destruct_d[0]} & {t4aeg_destruct_r,
                                                                                                                                         t3aef_destruct_r,
                                                                                                                                         t2aee_destruct_r,
                                                                                                                                         t1aed_destruct_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_r ? 4'd0 :
                                                            lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet24_5MQNode_6QNone_Int_2,QTree_Int) (lizzieLet24_5MQNode_6QNone_Int_1,QTree_Int) > [(_71,QTree_Int),
                                                                                                                    (_70,QTree_Int),
                                                                                                                    (lizzieLet24_5MQNode_6QNone_Int_1QNode_Int,QTree_Int),
                                                                                                                    (_69,QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_6QNone_Int_1_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_2_d[0] && lizzieLet24_5MQNode_6QNone_Int_1_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_2_d[2:1])
        2'd0: lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_6QNone_Int_1_onehotd = 4'd0;
  assign _71_d = {lizzieLet24_5MQNode_6QNone_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNone_Int_1_onehotd[0]};
  assign _70_d = {lizzieLet24_5MQNode_6QNone_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNone_Int_1_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_d = {lizzieLet24_5MQNode_6QNone_Int_1_d[66:1],
                                                        lizzieLet24_5MQNode_6QNone_Int_1_onehotd[2]};
  assign _69_d = {lizzieLet24_5MQNode_6QNone_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QNone_Int_1_onehotd[3]};
  assign lizzieLet24_5MQNode_6QNone_Int_1_r = (| (lizzieLet24_5MQNode_6QNone_Int_1_onehotd & {_69_r,
                                                                                              lizzieLet24_5MQNode_6QNone_Int_1QNode_Int_r,
                                                                                              _70_r,
                                                                                              _71_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_2_r = lizzieLet24_5MQNode_6QNone_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_3,QTree_Int) (lizzieLet24_5MQNode_10QNone_Int,Pointer_MaskQTree) > [(_68,Pointer_MaskQTree),
                                                                                                                                   (_67,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int,Pointer_MaskQTree),
                                                                                                                                   (_66,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_10QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_3_d[0] && lizzieLet24_5MQNode_10QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_3_d[2:1])
        2'd0: lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_10QNone_Int_onehotd = 4'd0;
  assign _68_d = {lizzieLet24_5MQNode_10QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_10QNone_Int_onehotd[0]};
  assign _67_d = {lizzieLet24_5MQNode_10QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_10QNone_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_d = {lizzieLet24_5MQNode_10QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_10QNone_Int_onehotd[2]};
  assign _66_d = {lizzieLet24_5MQNode_10QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_10QNone_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_10QNone_Int_r = (| (lizzieLet24_5MQNode_10QNone_Int_onehotd & {_66_r,
                                                                                            lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_r,
                                                                                            _67_r,
                                                                                            _68_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_3_r = lizzieLet24_5MQNode_10QNone_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_4,QTree_Int) (lizzieLet24_5MQNode_11QNone_Int,Pointer_MaskQTree) > [(_65,Pointer_MaskQTree),
                                                                                                                                   (_64,Pointer_MaskQTree),
                                                                                                                                   (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int,Pointer_MaskQTree),
                                                                                                                                   (_63,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_11QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_4_d[0] && lizzieLet24_5MQNode_11QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_4_d[2:1])
        2'd0: lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_11QNone_Int_onehotd = 4'd0;
  assign _65_d = {lizzieLet24_5MQNode_11QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_11QNone_Int_onehotd[0]};
  assign _64_d = {lizzieLet24_5MQNode_11QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_11QNone_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_d = {lizzieLet24_5MQNode_11QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_11QNone_Int_onehotd[2]};
  assign _63_d = {lizzieLet24_5MQNode_11QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_11QNone_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_11QNone_Int_r = (| (lizzieLet24_5MQNode_11QNone_Int_onehotd & {_63_r,
                                                                                            lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_r,
                                                                                            _64_r,
                                                                                            _65_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_4_r = lizzieLet24_5MQNode_11QNone_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNone_Int_5,QTree_Int) (lizzieLet24_5MQNode_3QNone_Int,Pointer_CTf_f_Int) > [(lizzieLet24_5MQNode_6QNone_Int_5QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                  (lizzieLet24_5MQNode_6QNone_Int_5QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet24_5MQNode_3QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_5_d[0] && lizzieLet24_5MQNode_3QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_5_d[2:1])
        2'd0: lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_3QNone_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_d = {lizzieLet24_5MQNode_3QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_3QNone_Int_onehotd[0]};
  assign lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_d = {lizzieLet24_5MQNode_3QNone_Int_d[16:1],
                                                       lizzieLet24_5MQNode_3QNone_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_d = {lizzieLet24_5MQNode_3QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_3QNone_Int_onehotd[2]};
  assign lizzieLet24_5MQNode_6QNone_Int_5QError_Int_d = {lizzieLet24_5MQNode_3QNone_Int_d[16:1],
                                                         lizzieLet24_5MQNode_3QNone_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_3QNone_Int_r = (| (lizzieLet24_5MQNode_3QNone_Int_onehotd & {lizzieLet24_5MQNode_6QNone_Int_5QError_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_5_r = lizzieLet24_5MQNode_3QNone_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNone_Int_5QError_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_5QError_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_5QError_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_5QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_5QError_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_5QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_5QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNone_Int_5QNone_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_5QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6,QTree_Int) (lizzieLet24_5MQNode_4QNone_Int,Go) > [(lizzieLet24_5MQNode_6QNone_Int_6QNone_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int,Go),
                                                                                                    (lizzieLet24_5MQNode_6QNone_Int_6QError_Int,Go)] */
  logic [3:0] lizzieLet24_5MQNode_4QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_6_d[0] && lizzieLet24_5MQNode_4QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_6_d[2:1])
        2'd0: lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_4QNone_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_d = lizzieLet24_5MQNode_4QNone_Int_onehotd[0];
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_d = lizzieLet24_5MQNode_4QNone_Int_onehotd[1];
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d = lizzieLet24_5MQNode_4QNone_Int_onehotd[2];
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_d = lizzieLet24_5MQNode_4QNone_Int_onehotd[3];
  assign lizzieLet24_5MQNode_4QNone_Int_r = (| (lizzieLet24_5MQNode_4QNone_Int_onehotd & {lizzieLet24_5MQNode_6QNone_Int_6QError_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_6_r = lizzieLet24_5MQNode_4QNone_Int_r;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QError_Int,Go) > [(lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1,Go),
                                                                  (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QError_Int_done;
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_d = (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_d = (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_done = (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted | ({lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_d[0],
                                                                                                                   lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_r,
                                                                                                                                                                         lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_6QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_r ? 2'd0 :
                                                             lizzieLet24_5MQNode_6QNone_Int_6QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1,Go)] > (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_r && lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int,QTree_Int) > (lizzieLet31_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                           1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                               1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_r)
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf :
                                                                  lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int,Go) > [(lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1,Go),
                                                                 (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2,Go),
                                                                 (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3,Go),
                                                                 (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4,Go),
                                                                 (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5,Go)] */
  logic [4:0] lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted;
  logic [4:0] lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_done;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted[2]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted[3]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted[4]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_done = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted | ({lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted <= 5'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_r ? 5'd0 :
                                                            lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_done);
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf,Pointer_MaskQTree),
                                                             (t4aeg_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_d[0],
                                                                                                                                             lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_d[0],
                                                                                                                                             t4aeg_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_d, lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_d, t4aeg_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_4QNode_Int_1_argbuf_r,
          t4aeg_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf,Pointer_MaskQTree),
                                                             (t3aef_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_d[0],
                                                                                                                                            t3aef_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_d, lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_d, t3aef_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_2_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_3QNode_Int_1_argbuf_r,
          t3aef_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int2_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf,Pointer_MaskQTree),
                                                             (t2aee_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_d[0],
                                                                                                                                            t2aee_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_d, lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_d, t2aee_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_3_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_r,
          t2aee_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int3_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_MaskQTree___Pointer_QTree_Int,
      Dcon TupGo___Pointer_MaskQTree___Pointer_QTree_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf,Go),
                                                             (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf,Pointer_MaskQTree),
                                                             (t1aed_1_argbuf,Pointer_QTree_Int)] > (f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4,TupGo___Pointer_MaskQTree___Pointer_QTree_Int) */
  assign \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_d  = TupGo___Pointer_MaskQTree___Pointer_QTree_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_d[0],
                                                                                                                                            lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_d[0],
                                                                                                                                            t1aed_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_d, lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_d, t1aed_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_4_argbuf_r,
          lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_r,
          t1aed_1_argbuf_r} = {3 {(\f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_r  && \f'''''''''_f'''''''''_IntTupGo___Pointer_MaskQTree___Pointer_QTree_Int4_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNode_Int_5_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int,Go) > [(lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1,Go),
                                                                 (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_done;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_d = (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_d = (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_done = (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted | ({lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_r ? 2'd0 :
                                                            lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1,Go)] > (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_r && lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet28_2_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d <= {66'd0,
                                                                         1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet28_2_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf :
                                     lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                           1'd0};
    else
      if ((lizzieLet28_2_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
      else if (((! lizzieLet28_2_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_r)
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QNone_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int,Go) > [(lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1,Go),
                                                                (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_done;
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_d = (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_d = (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_done = (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted | ({lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_d[0],
                                                                                                               lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_d[0]} & {lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_r,
                                                                                                                                                                   lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_r = (& lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_emitted <= (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_r ? 2'd0 :
                                                           lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1,Go)] > (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_d[0]}), lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_d);
  assign {lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_r && lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int,QTree_Int) > (lizzieLet29_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                         1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet29_1_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf :
                                     lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                           1'd0};
    else
      if ((lizzieLet29_1_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
      else if (((! lizzieLet29_1_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2,Go) > (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_r = ((! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_r)
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_6QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_7,QTree_Int) (lizzieLet24_5MQNode_8QNone_Int,Pointer_MaskQTree) > [(_62,Pointer_MaskQTree),
                                                                                                                                  (_61,Pointer_MaskQTree),
                                                                                                                                  (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int,Pointer_MaskQTree),
                                                                                                                                  (_60,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_8QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_7_d[0] && lizzieLet24_5MQNode_8QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_7_d[2:1])
        2'd0: lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_8QNone_Int_onehotd = 4'd0;
  assign _62_d = {lizzieLet24_5MQNode_8QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_8QNone_Int_onehotd[0]};
  assign _61_d = {lizzieLet24_5MQNode_8QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_8QNone_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_d = {lizzieLet24_5MQNode_8QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_8QNone_Int_onehotd[2]};
  assign _60_d = {lizzieLet24_5MQNode_8QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_8QNone_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_8QNone_Int_r = (| (lizzieLet24_5MQNode_8QNone_Int_onehotd & {_60_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_r,
                                                                                          _61_r,
                                                                                          _62_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_7_r = lizzieLet24_5MQNode_8QNone_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_7QNode_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_8,QTree_Int) (lizzieLet24_5MQNode_9QNone_Int,Pointer_MaskQTree) > [(_59,Pointer_MaskQTree),
                                                                                                                                  (_58,Pointer_MaskQTree),
                                                                                                                                  (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int,Pointer_MaskQTree),
                                                                                                                                  (_57,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet24_5MQNode_9QNone_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QNone_Int_8_d[0] && lizzieLet24_5MQNode_9QNone_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QNone_Int_8_d[2:1])
        2'd0: lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_9QNone_Int_onehotd = 4'd0;
  assign _59_d = {lizzieLet24_5MQNode_9QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_9QNone_Int_onehotd[0]};
  assign _58_d = {lizzieLet24_5MQNode_9QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_9QNone_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_d = {lizzieLet24_5MQNode_9QNone_Int_d[16:1],
                                                        lizzieLet24_5MQNode_9QNone_Int_onehotd[2]};
  assign _57_d = {lizzieLet24_5MQNode_9QNone_Int_d[16:1],
                  lizzieLet24_5MQNode_9QNone_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_9QNone_Int_r = (| (lizzieLet24_5MQNode_9QNone_Int_onehotd & {_57_r,
                                                                                          lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_r,
                                                                                          _58_r,
                                                                                          _59_r}));
  assign lizzieLet24_5MQNode_6QNone_Int_8_r = lizzieLet24_5MQNode_9QNone_Int_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int,Pointer_MaskQTree) > (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_r = ((! lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_r)
        lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QNone_Int_8QNode_Int_bufchan_d;
  
  /* fork (Ty QTree_Int) : (lizzieLet24_5MQNode_6QVal_Int,QTree_Int) > [(lizzieLet24_5MQNode_6QVal_Int_1,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_2,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_3,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_4,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_5,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_6,QTree_Int),
                                                                   (lizzieLet24_5MQNode_6QVal_Int_7,QTree_Int)] */
  logic [6:0] lizzieLet24_5MQNode_6QVal_Int_emitted;
  logic [6:0] lizzieLet24_5MQNode_6QVal_Int_done;
  assign lizzieLet24_5MQNode_6QVal_Int_1_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[0]))};
  assign lizzieLet24_5MQNode_6QVal_Int_2_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[1]))};
  assign lizzieLet24_5MQNode_6QVal_Int_3_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[2]))};
  assign lizzieLet24_5MQNode_6QVal_Int_4_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[3]))};
  assign lizzieLet24_5MQNode_6QVal_Int_5_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[4]))};
  assign lizzieLet24_5MQNode_6QVal_Int_6_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[5]))};
  assign lizzieLet24_5MQNode_6QVal_Int_7_d = {lizzieLet24_5MQNode_6QVal_Int_d[66:1],
                                              (lizzieLet24_5MQNode_6QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_emitted[6]))};
  assign lizzieLet24_5MQNode_6QVal_Int_done = (lizzieLet24_5MQNode_6QVal_Int_emitted | ({lizzieLet24_5MQNode_6QVal_Int_7_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_6_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_5_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_4_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_3_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_2_d[0],
                                                                                         lizzieLet24_5MQNode_6QVal_Int_1_d[0]} & {lizzieLet24_5MQNode_6QVal_Int_7_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_6_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_5_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_4_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_3_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_2_r,
                                                                                                                                  lizzieLet24_5MQNode_6QVal_Int_1_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_r = (& lizzieLet24_5MQNode_6QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_5MQNode_6QVal_Int_emitted <= 7'd0;
    else
      lizzieLet24_5MQNode_6QVal_Int_emitted <= (lizzieLet24_5MQNode_6QVal_Int_r ? 7'd0 :
                                                lizzieLet24_5MQNode_6QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet24_5MQNode_6QVal_Int_1QVal_Int,QTree_Int) > [(vaei_destruct,Int)] */
  assign vaei_destruct_d = {lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_r = vaei_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet24_5MQNode_6QVal_Int_2,QTree_Int) (lizzieLet24_5MQNode_6QVal_Int_1,QTree_Int) > [(_56,QTree_Int),
                                                                                                                  (lizzieLet24_5MQNode_6QVal_Int_1QVal_Int,QTree_Int),
                                                                                                                  (_55,QTree_Int),
                                                                                                                  (_54,QTree_Int)] */
  logic [3:0] lizzieLet24_5MQNode_6QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_2_d[0] && lizzieLet24_5MQNode_6QVal_Int_1_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_2_d[2:1])
        2'd0: lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_6QVal_Int_1_onehotd = 4'd0;
  assign _56_d = {lizzieLet24_5MQNode_6QVal_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QVal_Int_1_onehotd[0]};
  assign lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_d = {lizzieLet24_5MQNode_6QVal_Int_1_d[66:1],
                                                      lizzieLet24_5MQNode_6QVal_Int_1_onehotd[1]};
  assign _55_d = {lizzieLet24_5MQNode_6QVal_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QVal_Int_1_onehotd[2]};
  assign _54_d = {lizzieLet24_5MQNode_6QVal_Int_1_d[66:1],
                  lizzieLet24_5MQNode_6QVal_Int_1_onehotd[3]};
  assign lizzieLet24_5MQNode_6QVal_Int_1_r = (| (lizzieLet24_5MQNode_6QVal_Int_1_onehotd & {_54_r,
                                                                                            _55_r,
                                                                                            lizzieLet24_5MQNode_6QVal_Int_1QVal_Int_r,
                                                                                            _56_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_2_r = lizzieLet24_5MQNode_6QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QVal_Int_3,QTree_Int) (lizzieLet24_5MQNode_3QVal_Int,Pointer_CTf_f_Int) > [(lizzieLet24_5MQNode_6QVal_Int_3QNone_Int,Pointer_CTf_f_Int),
                                                                                                                                (lizzieLet24_5MQNode_6QVal_Int_3QVal_Int,Pointer_CTf_f_Int),
                                                                                                                                (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int,Pointer_CTf_f_Int),
                                                                                                                                (lizzieLet24_5MQNode_6QVal_Int_3QError_Int,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet24_5MQNode_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_3_d[0] && lizzieLet24_5MQNode_3QVal_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_3_d[2:1])
        2'd0: lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_d = {lizzieLet24_5MQNode_3QVal_Int_d[16:1],
                                                       lizzieLet24_5MQNode_3QVal_Int_onehotd[0]};
  assign lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_d = {lizzieLet24_5MQNode_3QVal_Int_d[16:1],
                                                      lizzieLet24_5MQNode_3QVal_Int_onehotd[1]};
  assign lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_d = {lizzieLet24_5MQNode_3QVal_Int_d[16:1],
                                                       lizzieLet24_5MQNode_3QVal_Int_onehotd[2]};
  assign lizzieLet24_5MQNode_6QVal_Int_3QError_Int_d = {lizzieLet24_5MQNode_3QVal_Int_d[16:1],
                                                        lizzieLet24_5MQNode_3QVal_Int_onehotd[3]};
  assign lizzieLet24_5MQNode_3QVal_Int_r = (| (lizzieLet24_5MQNode_3QVal_Int_onehotd & {lizzieLet24_5MQNode_6QVal_Int_3QError_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_3QVal_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_3_r = lizzieLet24_5MQNode_3QVal_Int_r;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QVal_Int_3QError_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_3QError_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_3QError_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_3QError_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet24_5MQNode_6QVal_Int_3QError_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_3QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_3QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (lizzieLet24_5MQNode_6QVal_Int_3QNone_Int,Pointer_CTf_f_Int) > (lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_d;
  Pointer_CTf_f_Int_t lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_3QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4,QTree_Int) (lizzieLet24_5MQNode_4QVal_Int,Go) > [(lizzieLet24_5MQNode_6QVal_Int_4QNone_Int,Go),
                                                                                                  (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int,Go),
                                                                                                  (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int,Go),
                                                                                                  (lizzieLet24_5MQNode_6QVal_Int_4QError_Int,Go)] */
  logic [3:0] lizzieLet24_5MQNode_4QVal_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_4_d[0] && lizzieLet24_5MQNode_4QVal_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_4_d[2:1])
        2'd0: lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_4QVal_Int_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_d = lizzieLet24_5MQNode_4QVal_Int_onehotd[0];
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_d = lizzieLet24_5MQNode_4QVal_Int_onehotd[1];
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_d = lizzieLet24_5MQNode_4QVal_Int_onehotd[2];
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_d = lizzieLet24_5MQNode_4QVal_Int_onehotd[3];
  assign lizzieLet24_5MQNode_4QVal_Int_r = (| (lizzieLet24_5MQNode_4QVal_Int_onehotd & {lizzieLet24_5MQNode_6QVal_Int_4QError_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_4_r = lizzieLet24_5MQNode_4QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QError_Int,Go) > [(lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1,Go),
                                                                 (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QError_Int_done;
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_d = (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_d = (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_done = (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted | ({lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_d[0],
                                                                                                                 lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_d[0]} & {lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_r,
                                                                                                                                                                      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_r = (& lizzieLet24_5MQNode_6QVal_Int_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_emitted <= (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_r ? 2'd0 :
                                                            lizzieLet24_5MQNode_6QVal_Int_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1,Go)] > (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_d[0]}), lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_d);
  assign {lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_r && lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet33_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                          1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet33_1_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                            1'd0};
    else
      if ((lizzieLet33_1_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                              1'd0};
      else if (((! lizzieLet33_1_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2,Go) > (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_r)
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf :
                                                                 lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int,Go) > [(lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1,Go),
                                                                (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_done;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_d = (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_d = (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_done = (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted | ({lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_d[0],
                                                                                                               lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_d[0]} & {lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_r,
                                                                                                                                                                   lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_r = (& lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_emitted <= (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_r ? 2'd0 :
                                                           lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1,Go)] > (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_d[0]}), lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_d);
  assign {lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_r && lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int,QTree_Int) > (lizzieLet36_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                         1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet36_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                           1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2,Go) > (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_r)
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QNode_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int,Go) > [(lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1,Go),
                                                                (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_done;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_d = (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_d = (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_done = (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted | ({lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_d[0],
                                                                                                               lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_d[0]} & {lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_r,
                                                                                                                                                                   lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_r = (& lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_emitted <= (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_r ? 2'd0 :
                                                           lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1,Go)] > (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int,QTree_Int) */
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_d[0]}), lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_d);
  assign {lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1_r} = {1 {(lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_r && lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int,QTree_Int) > (lizzieLet33_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                         1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_d;
  QTree_Int_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet33_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf :
                                   lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                           1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                             1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2,Go) > (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_r)
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_d;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf :
                                                                lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QNone_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int,Go) > [(lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1,Go),
                                                               (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted;
  logic [1:0] lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_done;
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_d = (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted[0]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_d = (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_d[0] && (! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted[1]));
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_done = (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted | ({lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_d[0],
                                                                                                             lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_d[0]} & {lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_2_r,
                                                                                                                                                                lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_r = (& lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_emitted <= (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_r ? 2'd0 :
                                                          lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1,Go) > (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_r = ((! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_r)
        lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_d;
  Go_t lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf :
                                                               lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf,Go),
                                          (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_5_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_d[0],
                                                                                            lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_d[0],
                                                                                            es_5_1_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_d, lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_d, es_5_1_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QVal_Int_4QVal_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_r,
          es_5_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_6QVal_Int_5,QTree_Int) (lizzieLet24_5MQNode_5QVal_Int,MyDTInt_Bool) > [(_53,MyDTInt_Bool),
                                                                                                                      (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int,MyDTInt_Bool),
                                                                                                                      (_52,MyDTInt_Bool),
                                                                                                                      (_51,MyDTInt_Bool)] */
  logic [3:0] lizzieLet24_5MQNode_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_5_d[0] && lizzieLet24_5MQNode_5QVal_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_5_d[2:1])
        2'd0: lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_5QVal_Int_onehotd = 4'd0;
  assign _53_d = lizzieLet24_5MQNode_5QVal_Int_onehotd[0];
  assign lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_d = lizzieLet24_5MQNode_5QVal_Int_onehotd[1];
  assign _52_d = lizzieLet24_5MQNode_5QVal_Int_onehotd[2];
  assign _51_d = lizzieLet24_5MQNode_5QVal_Int_onehotd[3];
  assign lizzieLet24_5MQNode_5QVal_Int_r = (| (lizzieLet24_5MQNode_5QVal_Int_onehotd & {_51_r,
                                                                                        _52_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_r,
                                                                                        _53_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_5_r = lizzieLet24_5MQNode_5QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int,MyDTInt_Bool) > (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf :
                                                               lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_6QVal_Int_6,QTree_Int) (lizzieLet24_5MQNode_7QVal_Int,MyDTInt_Int_Int) > [(_50,MyDTInt_Int_Int),
                                                                                                                            (lizzieLet24_5MQNode_6QVal_Int_6QVal_Int,MyDTInt_Int_Int),
                                                                                                                            (_49,MyDTInt_Int_Int),
                                                                                                                            (_48,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet24_5MQNode_7QVal_Int_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_6_d[0] && lizzieLet24_5MQNode_7QVal_Int_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_6_d[2:1])
        2'd0: lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd8;
        default: lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet24_5MQNode_7QVal_Int_onehotd = 4'd0;
  assign _50_d = lizzieLet24_5MQNode_7QVal_Int_onehotd[0];
  assign lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_d = lizzieLet24_5MQNode_7QVal_Int_onehotd[1];
  assign _49_d = lizzieLet24_5MQNode_7QVal_Int_onehotd[2];
  assign _48_d = lizzieLet24_5MQNode_7QVal_Int_onehotd[3];
  assign lizzieLet24_5MQNode_7QVal_Int_r = (| (lizzieLet24_5MQNode_7QVal_Int_onehotd & {_48_r,
                                                                                        _49_r,
                                                                                        lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_r,
                                                                                        _50_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_6_r = lizzieLet24_5MQNode_7QVal_Int_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_6QVal_Int_6QVal_Int,MyDTInt_Int_Int) > (lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf :
                                                               lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf,Int),
                                              (vaei_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                                       lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_d[0],
                                                                                                       vaei_1_argbuf_d[0]}), lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_d, lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_d, vaei_1_argbuf_d);
  assign {lizzieLet24_5MQNode_6QVal_Int_6QVal_Int_1_argbuf_r,
          lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_r,
          vaei_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet24_5MQNode_6QVal_Int_7,QTree_Int) (v1aeh_destruct,Int) > [(_47,Int),
                                                                                     (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int,Int),
                                                                                     (_46,Int),
                                                                                     (_45,Int)] */
  logic [3:0] v1aeh_destruct_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_6QVal_Int_7_d[0] && v1aeh_destruct_d[0]))
      unique case (lizzieLet24_5MQNode_6QVal_Int_7_d[2:1])
        2'd0: v1aeh_destruct_onehotd = 4'd1;
        2'd1: v1aeh_destruct_onehotd = 4'd2;
        2'd2: v1aeh_destruct_onehotd = 4'd4;
        2'd3: v1aeh_destruct_onehotd = 4'd8;
        default: v1aeh_destruct_onehotd = 4'd0;
      endcase
    else v1aeh_destruct_onehotd = 4'd0;
  assign _47_d = {v1aeh_destruct_d[32:1], v1aeh_destruct_onehotd[0]};
  assign lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_d = {v1aeh_destruct_d[32:1],
                                                      v1aeh_destruct_onehotd[1]};
  assign _46_d = {v1aeh_destruct_d[32:1], v1aeh_destruct_onehotd[2]};
  assign _45_d = {v1aeh_destruct_d[32:1], v1aeh_destruct_onehotd[3]};
  assign v1aeh_destruct_r = (| (v1aeh_destruct_onehotd & {_45_r,
                                                          _46_r,
                                                          lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_r,
                                                          _47_r}));
  assign lizzieLet24_5MQNode_6QVal_Int_7_r = v1aeh_destruct_r;
  
  /* buf (Ty Int) : (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int,Int) > (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d;
  logic lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_r;
  assign lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_r = ((! lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d[0]) || lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_r)
        lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d <= lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_d;
  Int_t lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_r = (! lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_d = (lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf :
                                                               lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf <= {32'd0,
                                                              1'd0};
    else
      if ((lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_r && lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf <= {32'd0,
                                                                1'd0};
      else if (((! lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_buf <= lizzieLet24_5MQNode_6QVal_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet24_5MQNode_7,QTree_Int) (lizzieLet24_9MQNode,MyDTInt_Int_Int) > [(_44,MyDTInt_Int_Int),
                                                                                                        (lizzieLet24_5MQNode_7QVal_Int,MyDTInt_Int_Int),
                                                                                                        (lizzieLet24_5MQNode_7QNode_Int,MyDTInt_Int_Int),
                                                                                                        (_43,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet24_9MQNode_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_7_d[0] && lizzieLet24_9MQNode_d[0]))
      unique case (lizzieLet24_5MQNode_7_d[2:1])
        2'd0: lizzieLet24_9MQNode_onehotd = 4'd1;
        2'd1: lizzieLet24_9MQNode_onehotd = 4'd2;
        2'd2: lizzieLet24_9MQNode_onehotd = 4'd4;
        2'd3: lizzieLet24_9MQNode_onehotd = 4'd8;
        default: lizzieLet24_9MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet24_9MQNode_onehotd = 4'd0;
  assign _44_d = lizzieLet24_9MQNode_onehotd[0];
  assign lizzieLet24_5MQNode_7QVal_Int_d = lizzieLet24_9MQNode_onehotd[1];
  assign lizzieLet24_5MQNode_7QNode_Int_d = lizzieLet24_9MQNode_onehotd[2];
  assign _43_d = lizzieLet24_9MQNode_onehotd[3];
  assign lizzieLet24_9MQNode_r = (| (lizzieLet24_9MQNode_onehotd & {_43_r,
                                                                    lizzieLet24_5MQNode_7QNode_Int_r,
                                                                    lizzieLet24_5MQNode_7QVal_Int_r,
                                                                    _44_r}));
  assign lizzieLet24_5MQNode_7_r = lizzieLet24_9MQNode_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_8,QTree_Int) (q1ae8_destruct,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_8QNone_Int,Pointer_MaskQTree),
                                                                                                       (_42,Pointer_MaskQTree),
                                                                                                       (lizzieLet24_5MQNode_8QNode_Int,Pointer_MaskQTree),
                                                                                                       (_41,Pointer_MaskQTree)] */
  logic [3:0] q1ae8_destruct_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_8_d[0] && q1ae8_destruct_d[0]))
      unique case (lizzieLet24_5MQNode_8_d[2:1])
        2'd0: q1ae8_destruct_onehotd = 4'd1;
        2'd1: q1ae8_destruct_onehotd = 4'd2;
        2'd2: q1ae8_destruct_onehotd = 4'd4;
        2'd3: q1ae8_destruct_onehotd = 4'd8;
        default: q1ae8_destruct_onehotd = 4'd0;
      endcase
    else q1ae8_destruct_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_8QNone_Int_d = {q1ae8_destruct_d[16:1],
                                             q1ae8_destruct_onehotd[0]};
  assign _42_d = {q1ae8_destruct_d[16:1], q1ae8_destruct_onehotd[1]};
  assign lizzieLet24_5MQNode_8QNode_Int_d = {q1ae8_destruct_d[16:1],
                                             q1ae8_destruct_onehotd[2]};
  assign _41_d = {q1ae8_destruct_d[16:1], q1ae8_destruct_onehotd[3]};
  assign q1ae8_destruct_r = (| (q1ae8_destruct_onehotd & {_41_r,
                                                          lizzieLet24_5MQNode_8QNode_Int_r,
                                                          _42_r,
                                                          lizzieLet24_5MQNode_8QNone_Int_r}));
  assign lizzieLet24_5MQNode_8_r = q1ae8_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet24_5MQNode_9,QTree_Int) (q2ae9_destruct,Pointer_MaskQTree) > [(lizzieLet24_5MQNode_9QNone_Int,Pointer_MaskQTree),
                                                                                                       (_40,Pointer_MaskQTree),
                                                                                                       (lizzieLet24_5MQNode_9QNode_Int,Pointer_MaskQTree),
                                                                                                       (_39,Pointer_MaskQTree)] */
  logic [3:0] q2ae9_destruct_onehotd;
  always_comb
    if ((lizzieLet24_5MQNode_9_d[0] && q2ae9_destruct_d[0]))
      unique case (lizzieLet24_5MQNode_9_d[2:1])
        2'd0: q2ae9_destruct_onehotd = 4'd1;
        2'd1: q2ae9_destruct_onehotd = 4'd2;
        2'd2: q2ae9_destruct_onehotd = 4'd4;
        2'd3: q2ae9_destruct_onehotd = 4'd8;
        default: q2ae9_destruct_onehotd = 4'd0;
      endcase
    else q2ae9_destruct_onehotd = 4'd0;
  assign lizzieLet24_5MQNode_9QNone_Int_d = {q2ae9_destruct_d[16:1],
                                             q2ae9_destruct_onehotd[0]};
  assign _40_d = {q2ae9_destruct_d[16:1], q2ae9_destruct_onehotd[1]};
  assign lizzieLet24_5MQNode_9QNode_Int_d = {q2ae9_destruct_d[16:1],
                                             q2ae9_destruct_onehotd[2]};
  assign _39_d = {q2ae9_destruct_d[16:1], q2ae9_destruct_onehotd[3]};
  assign q2ae9_destruct_r = (| (q2ae9_destruct_onehotd & {_39_r,
                                                          lizzieLet24_5MQNode_9QNode_Int_r,
                                                          _40_r,
                                                          lizzieLet24_5MQNode_9QNone_Int_r}));
  assign lizzieLet24_5MQNode_9_r = q2ae9_destruct_r;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Int) : (lizzieLet24_6,MaskQTree) (readPointer_QTree_Intm3ae5_1_argbuf_rwb,QTree_Int) > [(_38,QTree_Int),
                                                                                                        (_37,QTree_Int),
                                                                                                        (lizzieLet24_6MQNode,QTree_Int)] */
  logic [2:0] readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet24_6_d[0] && readPointer_QTree_Intm3ae5_1_argbuf_rwb_d[0]))
      unique case (lizzieLet24_6_d[2:1])
        2'd0: readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd = 3'd0;
  assign _38_d = {readPointer_QTree_Intm3ae5_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd[0]};
  assign _37_d = {readPointer_QTree_Intm3ae5_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet24_6MQNode_d = {readPointer_QTree_Intm3ae5_1_argbuf_rwb_d[66:1],
                                  readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Intm3ae5_1_argbuf_rwb_r = (| (readPointer_QTree_Intm3ae5_1_argbuf_rwb_onehotd & {lizzieLet24_6MQNode_r,
                                                                                                            _37_r,
                                                                                                            _38_r}));
  assign lizzieLet24_6_r = readPointer_QTree_Intm3ae5_1_argbuf_rwb_r;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Int) : (lizzieLet24_7,MaskQTree) (m2ae4_2,Pointer_QTree_Int) > [(_36,Pointer_QTree_Int),
                                                                                        (lizzieLet24_7MQVal,Pointer_QTree_Int),
                                                                                        (_35,Pointer_QTree_Int)] */
  logic [2:0] m2ae4_2_onehotd;
  always_comb
    if ((lizzieLet24_7_d[0] && m2ae4_2_d[0]))
      unique case (lizzieLet24_7_d[2:1])
        2'd0: m2ae4_2_onehotd = 3'd1;
        2'd1: m2ae4_2_onehotd = 3'd2;
        2'd2: m2ae4_2_onehotd = 3'd4;
        default: m2ae4_2_onehotd = 3'd0;
      endcase
    else m2ae4_2_onehotd = 3'd0;
  assign _36_d = {m2ae4_2_d[16:1], m2ae4_2_onehotd[0]};
  assign lizzieLet24_7MQVal_d = {m2ae4_2_d[16:1],
                                 m2ae4_2_onehotd[1]};
  assign _35_d = {m2ae4_2_d[16:1], m2ae4_2_onehotd[2]};
  assign m2ae4_2_r = (| (m2ae4_2_onehotd & {_35_r,
                                            lizzieLet24_7MQVal_r,
                                            _36_r}));
  assign lizzieLet24_7_r = m2ae4_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_7MQVal,Pointer_QTree_Int) > (lizzieLet24_7MQVal_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_7MQVal_bufchan_d;
  logic lizzieLet24_7MQVal_bufchan_r;
  assign lizzieLet24_7MQVal_r = ((! lizzieLet24_7MQVal_bufchan_d[0]) || lizzieLet24_7MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_7MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet24_7MQVal_r)
        lizzieLet24_7MQVal_bufchan_d <= lizzieLet24_7MQVal_d;
  Pointer_QTree_Int_t lizzieLet24_7MQVal_bufchan_buf;
  assign lizzieLet24_7MQVal_bufchan_r = (! lizzieLet24_7MQVal_bufchan_buf[0]);
  assign lizzieLet24_7MQVal_1_argbuf_d = (lizzieLet24_7MQVal_bufchan_buf[0] ? lizzieLet24_7MQVal_bufchan_buf :
                                          lizzieLet24_7MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_7MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_7MQVal_1_argbuf_r && lizzieLet24_7MQVal_bufchan_buf[0]))
        lizzieLet24_7MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet24_7MQVal_1_argbuf_r) && (! lizzieLet24_7MQVal_bufchan_buf[0])))
        lizzieLet24_7MQVal_bufchan_buf <= lizzieLet24_7MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Int) : (lizzieLet24_8,MaskQTree) (m3ae5_2,Pointer_QTree_Int) > [(_34,Pointer_QTree_Int),
                                                                                        (lizzieLet24_8MQVal,Pointer_QTree_Int),
                                                                                        (_33,Pointer_QTree_Int)] */
  logic [2:0] m3ae5_2_onehotd;
  always_comb
    if ((lizzieLet24_8_d[0] && m3ae5_2_d[0]))
      unique case (lizzieLet24_8_d[2:1])
        2'd0: m3ae5_2_onehotd = 3'd1;
        2'd1: m3ae5_2_onehotd = 3'd2;
        2'd2: m3ae5_2_onehotd = 3'd4;
        default: m3ae5_2_onehotd = 3'd0;
      endcase
    else m3ae5_2_onehotd = 3'd0;
  assign _34_d = {m3ae5_2_d[16:1], m3ae5_2_onehotd[0]};
  assign lizzieLet24_8MQVal_d = {m3ae5_2_d[16:1],
                                 m3ae5_2_onehotd[1]};
  assign _33_d = {m3ae5_2_d[16:1], m3ae5_2_onehotd[2]};
  assign m3ae5_2_r = (| (m3ae5_2_onehotd & {_33_r,
                                            lizzieLet24_8MQVal_r,
                                            _34_r}));
  assign lizzieLet24_8_r = m3ae5_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_8MQVal,Pointer_QTree_Int) > (lizzieLet24_8MQVal_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_8MQVal_bufchan_d;
  logic lizzieLet24_8MQVal_bufchan_r;
  assign lizzieLet24_8MQVal_r = ((! lizzieLet24_8MQVal_bufchan_d[0]) || lizzieLet24_8MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_8MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet24_8MQVal_r)
        lizzieLet24_8MQVal_bufchan_d <= lizzieLet24_8MQVal_d;
  Pointer_QTree_Int_t lizzieLet24_8MQVal_bufchan_buf;
  assign lizzieLet24_8MQVal_bufchan_r = (! lizzieLet24_8MQVal_bufchan_buf[0]);
  assign lizzieLet24_8MQVal_1_argbuf_d = (lizzieLet24_8MQVal_bufchan_buf[0] ? lizzieLet24_8MQVal_bufchan_buf :
                                          lizzieLet24_8MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_8MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet24_8MQVal_1_argbuf_r && lizzieLet24_8MQVal_bufchan_buf[0]))
        lizzieLet24_8MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet24_8MQVal_1_argbuf_r) && (! lizzieLet24_8MQVal_bufchan_buf[0])))
        lizzieLet24_8MQVal_bufchan_buf <= lizzieLet24_8MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty MyDTInt_Int_Int) : (lizzieLet24_9,MaskQTree) (op_addae7_goMux_mux,MyDTInt_Int_Int) > [(_32,MyDTInt_Int_Int),
                                                                                                (lizzieLet24_9MQVal,MyDTInt_Int_Int),
                                                                                                (lizzieLet24_9MQNode,MyDTInt_Int_Int)] */
  logic [2:0] op_addae7_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_9_d[0] && op_addae7_goMux_mux_d[0]))
      unique case (lizzieLet24_9_d[2:1])
        2'd0: op_addae7_goMux_mux_onehotd = 3'd1;
        2'd1: op_addae7_goMux_mux_onehotd = 3'd2;
        2'd2: op_addae7_goMux_mux_onehotd = 3'd4;
        default: op_addae7_goMux_mux_onehotd = 3'd0;
      endcase
    else op_addae7_goMux_mux_onehotd = 3'd0;
  assign _32_d = op_addae7_goMux_mux_onehotd[0];
  assign lizzieLet24_9MQVal_d = op_addae7_goMux_mux_onehotd[1];
  assign lizzieLet24_9MQNode_d = op_addae7_goMux_mux_onehotd[2];
  assign op_addae7_goMux_mux_r = (| (op_addae7_goMux_mux_onehotd & {lizzieLet24_9MQNode_r,
                                                                    lizzieLet24_9MQVal_r,
                                                                    _32_r}));
  assign lizzieLet24_9_r = op_addae7_goMux_mux_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet24_9MQVal,MyDTInt_Int_Int) > (lizzieLet24_9MQVal_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet24_9MQVal_bufchan_d;
  logic lizzieLet24_9MQVal_bufchan_r;
  assign lizzieLet24_9MQVal_r = ((! lizzieLet24_9MQVal_bufchan_d[0]) || lizzieLet24_9MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_9MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_9MQVal_r)
        lizzieLet24_9MQVal_bufchan_d <= lizzieLet24_9MQVal_d;
  MyDTInt_Int_Int_t lizzieLet24_9MQVal_bufchan_buf;
  assign lizzieLet24_9MQVal_bufchan_r = (! lizzieLet24_9MQVal_bufchan_buf[0]);
  assign lizzieLet24_9MQVal_1_argbuf_d = (lizzieLet24_9MQVal_bufchan_buf[0] ? lizzieLet24_9MQVal_bufchan_buf :
                                          lizzieLet24_9MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_9MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_9MQVal_1_argbuf_r && lizzieLet24_9MQVal_bufchan_buf[0]))
        lizzieLet24_9MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_9MQVal_1_argbuf_r) && (! lizzieLet24_9MQVal_bufchan_buf[0])))
        lizzieLet24_9MQVal_bufchan_buf <= lizzieLet24_9MQVal_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_main1_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                     (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_main1_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_main1_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_main1_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_main1_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_main1_3I#_3_onehotd [1];
  assign \arg0_1Dcon_main1_3I#_3_r  = (| (\arg0_1Dcon_main1_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                              lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_main1_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int0) : (lizzieLet46_1Lcall_$wnnz_Int0,CT$wnnz_Int) > [(wwsjT_4_destruct,Int#),
                                                                                  (ww1Xkr_2_destruct,Int#),
                                                                                  (ww2Xku_1_destruct,Int#),
                                                                                  (sc_0_7_destruct,Pointer_CT$wnnz_Int)] */
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int0_emitted;
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int0_done;
  assign wwsjT_4_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int0_d[35:4],
                               (lizzieLet46_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int0_emitted[0]))};
  assign ww1Xkr_2_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int0_d[67:36],
                                (lizzieLet46_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int0_emitted[1]))};
  assign ww2Xku_1_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int0_d[99:68],
                                (lizzieLet46_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int0_emitted[2]))};
  assign sc_0_7_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int0_d[115:100],
                              (lizzieLet46_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int0_emitted[3]))};
  assign lizzieLet46_1Lcall_$wnnz_Int0_done = (lizzieLet46_1Lcall_$wnnz_Int0_emitted | ({sc_0_7_destruct_d[0],
                                                                                         ww2Xku_1_destruct_d[0],
                                                                                         ww1Xkr_2_destruct_d[0],
                                                                                         wwsjT_4_destruct_d[0]} & {sc_0_7_destruct_r,
                                                                                                                   ww2Xku_1_destruct_r,
                                                                                                                   ww1Xkr_2_destruct_r,
                                                                                                                   wwsjT_4_destruct_r}));
  assign lizzieLet46_1Lcall_$wnnz_Int0_r = (& lizzieLet46_1Lcall_$wnnz_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet46_1Lcall_$wnnz_Int0_emitted <= 4'd0;
    else
      lizzieLet46_1Lcall_$wnnz_Int0_emitted <= (lizzieLet46_1Lcall_$wnnz_Int0_r ? 4'd0 :
                                                lizzieLet46_1Lcall_$wnnz_Int0_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int1) : (lizzieLet46_1Lcall_$wnnz_Int1,CT$wnnz_Int) > [(wwsjT_3_destruct,Int#),
                                                                                  (ww1Xkr_1_destruct,Int#),
                                                                                  (sc_0_6_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a88_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int1_emitted;
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int1_done;
  assign wwsjT_3_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int1_d[35:4],
                               (lizzieLet46_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int1_emitted[0]))};
  assign ww1Xkr_1_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int1_d[67:36],
                                (lizzieLet46_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int1_emitted[1]))};
  assign sc_0_6_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int1_d[83:68],
                              (lizzieLet46_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int1_emitted[2]))};
  assign q4a88_3_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int1_d[99:84],
                               (lizzieLet46_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int1_emitted[3]))};
  assign lizzieLet46_1Lcall_$wnnz_Int1_done = (lizzieLet46_1Lcall_$wnnz_Int1_emitted | ({q4a88_3_destruct_d[0],
                                                                                         sc_0_6_destruct_d[0],
                                                                                         ww1Xkr_1_destruct_d[0],
                                                                                         wwsjT_3_destruct_d[0]} & {q4a88_3_destruct_r,
                                                                                                                   sc_0_6_destruct_r,
                                                                                                                   ww1Xkr_1_destruct_r,
                                                                                                                   wwsjT_3_destruct_r}));
  assign lizzieLet46_1Lcall_$wnnz_Int1_r = (& lizzieLet46_1Lcall_$wnnz_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet46_1Lcall_$wnnz_Int1_emitted <= 4'd0;
    else
      lizzieLet46_1Lcall_$wnnz_Int1_emitted <= (lizzieLet46_1Lcall_$wnnz_Int1_r ? 4'd0 :
                                                lizzieLet46_1Lcall_$wnnz_Int1_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int2) : (lizzieLet46_1Lcall_$wnnz_Int2,CT$wnnz_Int) > [(wwsjT_2_destruct,Int#),
                                                                                  (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a88_2_destruct,Pointer_QTree_Int),
                                                                                  (q3a87_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int2_emitted;
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int2_done;
  assign wwsjT_2_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int2_d[35:4],
                               (lizzieLet46_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int2_emitted[0]))};
  assign sc_0_5_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int2_d[51:36],
                              (lizzieLet46_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int2_emitted[1]))};
  assign q4a88_2_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int2_d[67:52],
                               (lizzieLet46_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int2_emitted[2]))};
  assign q3a87_2_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int2_d[83:68],
                               (lizzieLet46_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int2_emitted[3]))};
  assign lizzieLet46_1Lcall_$wnnz_Int2_done = (lizzieLet46_1Lcall_$wnnz_Int2_emitted | ({q3a87_2_destruct_d[0],
                                                                                         q4a88_2_destruct_d[0],
                                                                                         sc_0_5_destruct_d[0],
                                                                                         wwsjT_2_destruct_d[0]} & {q3a87_2_destruct_r,
                                                                                                                   q4a88_2_destruct_r,
                                                                                                                   sc_0_5_destruct_r,
                                                                                                                   wwsjT_2_destruct_r}));
  assign lizzieLet46_1Lcall_$wnnz_Int2_r = (& lizzieLet46_1Lcall_$wnnz_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet46_1Lcall_$wnnz_Int2_emitted <= 4'd0;
    else
      lizzieLet46_1Lcall_$wnnz_Int2_emitted <= (lizzieLet46_1Lcall_$wnnz_Int2_r ? 4'd0 :
                                                lizzieLet46_1Lcall_$wnnz_Int2_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int3) : (lizzieLet46_1Lcall_$wnnz_Int3,CT$wnnz_Int) > [(sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4a88_1_destruct,Pointer_QTree_Int),
                                                                                  (q3a87_1_destruct,Pointer_QTree_Int),
                                                                                  (q2a86_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int3_emitted;
  logic [3:0] lizzieLet46_1Lcall_$wnnz_Int3_done;
  assign sc_0_4_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int3_d[19:4],
                              (lizzieLet46_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int3_emitted[0]))};
  assign q4a88_1_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int3_d[35:20],
                               (lizzieLet46_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int3_emitted[1]))};
  assign q3a87_1_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int3_d[51:36],
                               (lizzieLet46_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int3_emitted[2]))};
  assign q2a86_1_destruct_d = {lizzieLet46_1Lcall_$wnnz_Int3_d[67:52],
                               (lizzieLet46_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet46_1Lcall_$wnnz_Int3_emitted[3]))};
  assign lizzieLet46_1Lcall_$wnnz_Int3_done = (lizzieLet46_1Lcall_$wnnz_Int3_emitted | ({q2a86_1_destruct_d[0],
                                                                                         q3a87_1_destruct_d[0],
                                                                                         q4a88_1_destruct_d[0],
                                                                                         sc_0_4_destruct_d[0]} & {q2a86_1_destruct_r,
                                                                                                                  q3a87_1_destruct_r,
                                                                                                                  q4a88_1_destruct_r,
                                                                                                                  sc_0_4_destruct_r}));
  assign lizzieLet46_1Lcall_$wnnz_Int3_r = (& lizzieLet46_1Lcall_$wnnz_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet46_1Lcall_$wnnz_Int3_emitted <= 4'd0;
    else
      lizzieLet46_1Lcall_$wnnz_Int3_emitted <= (lizzieLet46_1Lcall_$wnnz_Int3_r ? 4'd0 :
                                                lizzieLet46_1Lcall_$wnnz_Int3_done);
  
  /* demux (Ty CT$wnnz_Int,
       Ty CT$wnnz_Int) : (lizzieLet46_2,CT$wnnz_Int) (lizzieLet46_1,CT$wnnz_Int) > [(_31,CT$wnnz_Int),
                                                                                    (lizzieLet46_1Lcall_$wnnz_Int3,CT$wnnz_Int),
                                                                                    (lizzieLet46_1Lcall_$wnnz_Int2,CT$wnnz_Int),
                                                                                    (lizzieLet46_1Lcall_$wnnz_Int1,CT$wnnz_Int),
                                                                                    (lizzieLet46_1Lcall_$wnnz_Int0,CT$wnnz_Int)] */
  logic [4:0] lizzieLet46_1_onehotd;
  always_comb
    if ((lizzieLet46_2_d[0] && lizzieLet46_1_d[0]))
      unique case (lizzieLet46_2_d[3:1])
        3'd0: lizzieLet46_1_onehotd = 5'd1;
        3'd1: lizzieLet46_1_onehotd = 5'd2;
        3'd2: lizzieLet46_1_onehotd = 5'd4;
        3'd3: lizzieLet46_1_onehotd = 5'd8;
        3'd4: lizzieLet46_1_onehotd = 5'd16;
        default: lizzieLet46_1_onehotd = 5'd0;
      endcase
    else lizzieLet46_1_onehotd = 5'd0;
  assign _31_d = {lizzieLet46_1_d[115:1], lizzieLet46_1_onehotd[0]};
  assign lizzieLet46_1Lcall_$wnnz_Int3_d = {lizzieLet46_1_d[115:1],
                                            lizzieLet46_1_onehotd[1]};
  assign lizzieLet46_1Lcall_$wnnz_Int2_d = {lizzieLet46_1_d[115:1],
                                            lizzieLet46_1_onehotd[2]};
  assign lizzieLet46_1Lcall_$wnnz_Int1_d = {lizzieLet46_1_d[115:1],
                                            lizzieLet46_1_onehotd[3]};
  assign lizzieLet46_1Lcall_$wnnz_Int0_d = {lizzieLet46_1_d[115:1],
                                            lizzieLet46_1_onehotd[4]};
  assign lizzieLet46_1_r = (| (lizzieLet46_1_onehotd & {lizzieLet46_1Lcall_$wnnz_Int0_r,
                                                        lizzieLet46_1Lcall_$wnnz_Int1_r,
                                                        lizzieLet46_1Lcall_$wnnz_Int2_r,
                                                        lizzieLet46_1Lcall_$wnnz_Int3_r,
                                                        _31_r}));
  assign lizzieLet46_2_r = lizzieLet46_1_r;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Go) : (lizzieLet46_3,CT$wnnz_Int) (go_15_goMux_data,Go) > [(_30,Go),
                                                                     (lizzieLet46_3Lcall_$wnnz_Int3,Go),
                                                                     (lizzieLet46_3Lcall_$wnnz_Int2,Go),
                                                                     (lizzieLet46_3Lcall_$wnnz_Int1,Go),
                                                                     (lizzieLet46_3Lcall_$wnnz_Int0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet46_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet46_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _30_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet46_3Lcall_$wnnz_Int3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet46_3Lcall_$wnnz_Int2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet46_3Lcall_$wnnz_Int1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet46_3Lcall_$wnnz_Int0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet46_3Lcall_$wnnz_Int0_r,
                                                              lizzieLet46_3Lcall_$wnnz_Int1_r,
                                                              lizzieLet46_3Lcall_$wnnz_Int2_r,
                                                              lizzieLet46_3Lcall_$wnnz_Int3_r,
                                                              _30_r}));
  assign lizzieLet46_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet46_3Lcall_$wnnz_Int0,Go) > (lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf,Go) */
  Go_t lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d;
  logic lizzieLet46_3Lcall_$wnnz_Int0_bufchan_r;
  assign lizzieLet46_3Lcall_$wnnz_Int0_r = ((! lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d[0]) || lizzieLet46_3Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet46_3Lcall_$wnnz_Int0_r)
        lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d <= lizzieLet46_3Lcall_$wnnz_Int0_d;
  Go_t lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf;
  assign lizzieLet46_3Lcall_$wnnz_Int0_bufchan_r = (! lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_d = (lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf[0] ? lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf :
                                                     lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_r && lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf[0]))
        lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_r) && (! lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf[0])))
        lizzieLet46_3Lcall_$wnnz_Int0_bufchan_buf <= lizzieLet46_3Lcall_$wnnz_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet46_3Lcall_$wnnz_Int1,Go) > (lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf,Go) */
  Go_t lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d;
  logic lizzieLet46_3Lcall_$wnnz_Int1_bufchan_r;
  assign lizzieLet46_3Lcall_$wnnz_Int1_r = ((! lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d[0]) || lizzieLet46_3Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet46_3Lcall_$wnnz_Int1_r)
        lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d <= lizzieLet46_3Lcall_$wnnz_Int1_d;
  Go_t lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf;
  assign lizzieLet46_3Lcall_$wnnz_Int1_bufchan_r = (! lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_d = (lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf[0] ? lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf :
                                                     lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_r && lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf[0]))
        lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet46_3Lcall_$wnnz_Int1_1_argbuf_r) && (! lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf[0])))
        lizzieLet46_3Lcall_$wnnz_Int1_bufchan_buf <= lizzieLet46_3Lcall_$wnnz_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet46_3Lcall_$wnnz_Int2,Go) > (lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf,Go) */
  Go_t lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet46_3Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet46_3Lcall_$wnnz_Int2_r = ((! lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet46_3Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet46_3Lcall_$wnnz_Int2_r)
        lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d <= lizzieLet46_3Lcall_$wnnz_Int2_d;
  Go_t lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet46_3Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_d = (lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf :
                                                     lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_r && lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet46_3Lcall_$wnnz_Int2_1_argbuf_r) && (! lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet46_3Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet46_3Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet46_3Lcall_$wnnz_Int3,Go) > (lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf,Go) */
  Go_t lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet46_3Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet46_3Lcall_$wnnz_Int3_r = ((! lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet46_3Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet46_3Lcall_$wnnz_Int3_r)
        lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d <= lizzieLet46_3Lcall_$wnnz_Int3_d;
  Go_t lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet46_3Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_d = (lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf :
                                                     lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_r && lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet46_3Lcall_$wnnz_Int3_1_argbuf_r) && (! lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet46_3Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet46_3Lcall_$wnnz_Int3_bufchan_d;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Int#) : (lizzieLet46_4,CT$wnnz_Int) (srtarg_0_goMux_mux,Int#) > [(lizzieLet46_4L$wnnz_Intsbos,Int#),
                                                                           (lizzieLet46_4Lcall_$wnnz_Int3,Int#),
                                                                           (lizzieLet46_4Lcall_$wnnz_Int2,Int#),
                                                                           (lizzieLet46_4Lcall_$wnnz_Int1,Int#),
                                                                           (lizzieLet46_4Lcall_$wnnz_Int0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet46_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet46_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet46_4L$wnnz_Intsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                          srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet46_4Lcall_$wnnz_Int3_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet46_4Lcall_$wnnz_Int2_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet46_4Lcall_$wnnz_Int1_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet46_4Lcall_$wnnz_Int0_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet46_4Lcall_$wnnz_Int0_r,
                                                                  lizzieLet46_4Lcall_$wnnz_Int1_r,
                                                                  lizzieLet46_4Lcall_$wnnz_Int2_r,
                                                                  lizzieLet46_4Lcall_$wnnz_Int3_r,
                                                                  lizzieLet46_4L$wnnz_Intsbos_r}));
  assign lizzieLet46_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet46_4L$wnnz_Intsbos,Int#) > [(lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#),
                                                       (lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet46_4L$wnnz_Intsbos_emitted;
  logic [1:0] lizzieLet46_4L$wnnz_Intsbos_done;
  assign lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_d = {lizzieLet46_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet46_4L$wnnz_Intsbos_d[0] && (! lizzieLet46_4L$wnnz_Intsbos_emitted[0]))};
  assign lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_d = {lizzieLet46_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet46_4L$wnnz_Intsbos_d[0] && (! lizzieLet46_4L$wnnz_Intsbos_emitted[1]))};
  assign lizzieLet46_4L$wnnz_Intsbos_done = (lizzieLet46_4L$wnnz_Intsbos_emitted | ({lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                     lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet46_4L$wnnz_Intsbos_r = (& lizzieLet46_4L$wnnz_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet46_4L$wnnz_Intsbos_emitted <= 2'd0;
    else
      lizzieLet46_4L$wnnz_Intsbos_emitted <= (lizzieLet46_4L$wnnz_Intsbos_r ? 2'd0 :
                                              lizzieLet46_4L$wnnz_Intsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_Int_goConst,Go) */
  assign call_$wnnz_Int_goConst_d = lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_1_r = call_$wnnz_Int_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#) > ($wnnz_Int_resbuf,Int#) */
  \Int#_t  lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                     1'd0};
    else
      if (lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_Int_resbuf_d  = (lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                       1'd0};
    else
      if ((\$wnnz_Int_resbuf_r  && lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                         1'd0};
      else if (((! \$wnnz_Int_resbuf_r ) && (! lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet46_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int2) : [(lizzieLet46_4Lcall_$wnnz_Int3,Int#),
                                (sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                (q4a88_1_destruct,Pointer_QTree_Int),
                                (q3a87_1_destruct,Pointer_QTree_Int)] > (lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) */
  assign lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_d = Lcall_$wnnz_Int2_dc((& {lizzieLet46_4Lcall_$wnnz_Int3_d[0],
                                                                                                               sc_0_4_destruct_d[0],
                                                                                                               q4a88_1_destruct_d[0],
                                                                                                               q3a87_1_destruct_d[0]}), lizzieLet46_4Lcall_$wnnz_Int3_d, sc_0_4_destruct_d, q4a88_1_destruct_d, q3a87_1_destruct_d);
  assign {lizzieLet46_4Lcall_$wnnz_Int3_r,
          sc_0_4_destruct_r,
          q4a88_1_destruct_r,
          q3a87_1_destruct_r} = {4 {(lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_r && lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) > (lizzieLet47_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_r = ((! lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_r)
        lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d <= lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_d;
  CT$wnnz_Int_t lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet47_1_argbuf_d = (lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf :
                                   lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet47_1_argbuf_r && lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet47_1_argbuf_r) && (! lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet46_4Lcall_$wnnz_Int3_1sc_0_4_1q4a88_1_1q3a87_1_1Lcall_$wnnz_Int2_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1a85_destruct,Pointer_QTree_Int),
                                                                 (q2a86_destruct,Pointer_QTree_Int),
                                                                 (q3a87_destruct,Pointer_QTree_Int),
                                                                 (q4a88_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1a85_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2a86_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3a87_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4a88_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4a88_destruct_d[0],
                                                                         q3a87_destruct_d[0],
                                                                         q2a86_destruct_d[0],
                                                                         q1a85_destruct_d[0]} & {q4a88_destruct_r,
                                                                                                 q3a87_destruct_r,
                                                                                                 q2a86_destruct_r,
                                                                                                 q1a85_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_29,QTree_Int),
                                                                            (_28,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_27,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _29_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _28_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _27_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_27_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _28_r,
                                                      _29_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_8_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                 (lizzieLet4_3QVal_Int,Go),
                                                                 (lizzieLet4_3QNode_Int,Go),
                                                                 (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_8_goMux_data_onehotd = 4'd1;
        2'd1: go_8_goMux_data_onehotd = 4'd2;
        2'd2: go_8_goMux_data_onehotd = 4'd4;
        2'd3: go_8_goMux_data_onehotd = 4'd8;
        default: go_8_goMux_data_onehotd = 4'd0;
      endcase
    else go_8_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_8_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_8_goMux_data_onehotd[3];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                            lizzieLet4_3QNode_Int_r,
                                                            lizzieLet4_3QVal_Int_r,
                                                            lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_8_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet28_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet28_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet28_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet28_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet28_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C4) (go_15_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                            go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                      go_15_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_15_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet46_3Lcall_$wnnz_Int0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_15_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet29_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz_Int) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                (q4a88_destruct,Pointer_QTree_Int),
                                (q3a87_destruct,Pointer_QTree_Int),
                                (q2a86_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3,CT$wnnz_Int) */
  assign lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_d = Lcall_$wnnz_Int3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                                  q4a88_destruct_d[0],
                                                                                                  q3a87_destruct_d[0],
                                                                                                  q2a86_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4a88_destruct_d, q3a87_destruct_d, q2a86_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4a88_destruct_r,
          q3a87_destruct_r,
          q2a86_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_r && lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3,CT$wnnz_Int) > (lizzieLet5_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_r = ((! lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d <= {115'd0,
                                                                                 1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_r)
        lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d <= lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_d;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                     1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4a88_1q3a87_1q2a86_1Lcall_$wnnz_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Int,
          Dcon Lcall_f'''''''''_f'''''''''_Int0) : (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0,CTf'''''''''_f'''''''''_Int) > [(es_1_2_destruct,Pointer_QTree_Int),
                                                                                                                                  (es_2_3_destruct,Pointer_QTree_Int),
                                                                                                                                  (es_3_4_destruct,Pointer_QTree_Int),
                                                                                                                                  (sc_0_11_destruct,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [3:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted ;
  logic [3:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_done ;
  assign es_1_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [19:4],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted [0]))};
  assign es_2_3_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [35:20],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted [1]))};
  assign es_3_4_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [51:36],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted [2]))};
  assign sc_0_11_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [67:52],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted [3]))};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_done  = (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted  | ({sc_0_11_destruct_d[0],
                                                                                                                             es_3_4_destruct_d[0],
                                                                                                                             es_2_3_destruct_d[0],
                                                                                                                             es_1_2_destruct_d[0]} & {sc_0_11_destruct_r,
                                                                                                                                                      es_3_4_destruct_r,
                                                                                                                                                      es_2_3_destruct_r,
                                                                                                                                                      es_1_2_destruct_r}));
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_r  = (& \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted  <= 4'd0;
    else
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_emitted  <= (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_r  ? 4'd0 :
                                                                  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Int,
          Dcon Lcall_f'''''''''_f'''''''''_Int1) : (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1,CTf'''''''''_f'''''''''_Int) > [(es_2_2_destruct,Pointer_QTree_Int),
                                                                                                                                  (es_3_3_destruct,Pointer_QTree_Int),
                                                                                                                                  (sc_0_10_destruct,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                  (q1aey_3_destruct,Pointer_MaskQTree),
                                                                                                                                  (t1aeD_3_destruct,Pointer_QTree_Int)] */
  logic [4:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted ;
  logic [4:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_done ;
  assign es_2_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [19:4],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted [0]))};
  assign es_3_3_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [35:20],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted [1]))};
  assign sc_0_10_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [51:36],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted [2]))};
  assign q1aey_3_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [67:52],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted [3]))};
  assign t1aeD_3_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [83:68],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted [4]))};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_done  = (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted  | ({t1aeD_3_destruct_d[0],
                                                                                                                             q1aey_3_destruct_d[0],
                                                                                                                             sc_0_10_destruct_d[0],
                                                                                                                             es_3_3_destruct_d[0],
                                                                                                                             es_2_2_destruct_d[0]} & {t1aeD_3_destruct_r,
                                                                                                                                                      q1aey_3_destruct_r,
                                                                                                                                                      sc_0_10_destruct_r,
                                                                                                                                                      es_3_3_destruct_r,
                                                                                                                                                      es_2_2_destruct_r}));
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_r  = (& \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted  <= 5'd0;
    else
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_emitted  <= (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_r  ? 5'd0 :
                                                                  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Int,
          Dcon Lcall_f'''''''''_f'''''''''_Int2) : (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2,CTf'''''''''_f'''''''''_Int) > [(es_3_2_destruct,Pointer_QTree_Int),
                                                                                                                                  (sc_0_9_destruct,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                  (q1aey_2_destruct,Pointer_MaskQTree),
                                                                                                                                  (t1aeD_2_destruct,Pointer_QTree_Int),
                                                                                                                                  (q2aez_2_destruct,Pointer_MaskQTree),
                                                                                                                                  (t2aeE_2_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted ;
  logic [5:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_done ;
  assign es_3_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [19:4],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [0]))};
  assign sc_0_9_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [35:20],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [1]))};
  assign q1aey_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [51:36],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [2]))};
  assign t1aeD_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [67:52],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [3]))};
  assign q2aez_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [83:68],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [4]))};
  assign t2aeE_2_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [99:84],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted [5]))};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_done  = (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted  | ({t2aeE_2_destruct_d[0],
                                                                                                                             q2aez_2_destruct_d[0],
                                                                                                                             t1aeD_2_destruct_d[0],
                                                                                                                             q1aey_2_destruct_d[0],
                                                                                                                             sc_0_9_destruct_d[0],
                                                                                                                             es_3_2_destruct_d[0]} & {t2aeE_2_destruct_r,
                                                                                                                                                      q2aez_2_destruct_r,
                                                                                                                                                      t1aeD_2_destruct_r,
                                                                                                                                                      q1aey_2_destruct_r,
                                                                                                                                                      sc_0_9_destruct_r,
                                                                                                                                                      es_3_2_destruct_r}));
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_r  = (& \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted  <= 6'd0;
    else
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_emitted  <= (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_r  ? 6'd0 :
                                                                  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_done );
  
  /* destruct (Ty CTf'''''''''_f'''''''''_Int,
          Dcon Lcall_f'''''''''_f'''''''''_Int3) : (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3,CTf'''''''''_f'''''''''_Int) > [(sc_0_8_destruct,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                  (q1aey_1_destruct,Pointer_MaskQTree),
                                                                                                                                  (t1aeD_1_destruct,Pointer_QTree_Int),
                                                                                                                                  (q2aez_1_destruct,Pointer_MaskQTree),
                                                                                                                                  (t2aeE_1_destruct,Pointer_QTree_Int),
                                                                                                                                  (q3aeA_1_destruct,Pointer_MaskQTree),
                                                                                                                                  (t3aeF_1_destruct,Pointer_QTree_Int)] */
  logic [6:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted ;
  logic [6:0] \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_done ;
  assign sc_0_8_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [19:4],
                              (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [0]))};
  assign q1aey_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [35:20],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [1]))};
  assign t1aeD_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [51:36],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [2]))};
  assign q2aez_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [67:52],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [3]))};
  assign t2aeE_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [83:68],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [4]))};
  assign q3aeA_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [99:84],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [5]))};
  assign t3aeF_1_destruct_d = {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [115:100],
                               (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d [0] && (! \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted [6]))};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_done  = (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted  | ({t3aeF_1_destruct_d[0],
                                                                                                                             q3aeA_1_destruct_d[0],
                                                                                                                             t2aeE_1_destruct_d[0],
                                                                                                                             q2aez_1_destruct_d[0],
                                                                                                                             t1aeD_1_destruct_d[0],
                                                                                                                             q1aey_1_destruct_d[0],
                                                                                                                             sc_0_8_destruct_d[0]} & {t3aeF_1_destruct_r,
                                                                                                                                                      q3aeA_1_destruct_r,
                                                                                                                                                      t2aeE_1_destruct_r,
                                                                                                                                                      q2aez_1_destruct_r,
                                                                                                                                                      t1aeD_1_destruct_r,
                                                                                                                                                      q1aey_1_destruct_r,
                                                                                                                                                      sc_0_8_destruct_r}));
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_r  = (& \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted  <= 7'd0;
    else
      \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_emitted  <= (\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_r  ? 7'd0 :
                                                                  \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_done );
  
  /* demux (Ty CTf'''''''''_f'''''''''_Int,
       Ty CTf'''''''''_f'''''''''_Int) : (lizzieLet50_2,CTf'''''''''_f'''''''''_Int) (lizzieLet50_1,CTf'''''''''_f'''''''''_Int) > [(_26,CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3,CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2,CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1,CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0,CTf'''''''''_f'''''''''_Int)] */
  logic [4:0] lizzieLet50_1_onehotd;
  always_comb
    if ((lizzieLet50_2_d[0] && lizzieLet50_1_d[0]))
      unique case (lizzieLet50_2_d[3:1])
        3'd0: lizzieLet50_1_onehotd = 5'd1;
        3'd1: lizzieLet50_1_onehotd = 5'd2;
        3'd2: lizzieLet50_1_onehotd = 5'd4;
        3'd3: lizzieLet50_1_onehotd = 5'd8;
        3'd4: lizzieLet50_1_onehotd = 5'd16;
        default: lizzieLet50_1_onehotd = 5'd0;
      endcase
    else lizzieLet50_1_onehotd = 5'd0;
  assign _26_d = {lizzieLet50_1_d[115:1], lizzieLet50_1_onehotd[0]};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_d  = {lizzieLet50_1_d[115:1],
                                                              lizzieLet50_1_onehotd[1]};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_d  = {lizzieLet50_1_d[115:1],
                                                              lizzieLet50_1_onehotd[2]};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_d  = {lizzieLet50_1_d[115:1],
                                                              lizzieLet50_1_onehotd[3]};
  assign \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_d  = {lizzieLet50_1_d[115:1],
                                                              lizzieLet50_1_onehotd[4]};
  assign lizzieLet50_1_r = (| (lizzieLet50_1_onehotd & {\lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int0_r ,
                                                        \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int1_r ,
                                                        \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int2_r ,
                                                        \lizzieLet50_1Lcall_f'''''''''_f'''''''''_Int3_r ,
                                                        _26_r}));
  assign lizzieLet50_2_r = lizzieLet50_1_r;
  
  /* demux (Ty CTf'''''''''_f'''''''''_Int,
       Ty Go) : (lizzieLet50_3,CTf'''''''''_f'''''''''_Int) (go_16_goMux_data,Go) > [(_25,Go),
                                                                                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3,Go),
                                                                                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2,Go),
                                                                                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1,Go),
                                                                                     (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0,Go)] */
  logic [4:0] go_16_goMux_data_onehotd;
  always_comb
    if ((lizzieLet50_3_d[0] && go_16_goMux_data_d[0]))
      unique case (lizzieLet50_3_d[3:1])
        3'd0: go_16_goMux_data_onehotd = 5'd1;
        3'd1: go_16_goMux_data_onehotd = 5'd2;
        3'd2: go_16_goMux_data_onehotd = 5'd4;
        3'd3: go_16_goMux_data_onehotd = 5'd8;
        3'd4: go_16_goMux_data_onehotd = 5'd16;
        default: go_16_goMux_data_onehotd = 5'd0;
      endcase
    else go_16_goMux_data_onehotd = 5'd0;
  assign _25_d = go_16_goMux_data_onehotd[0];
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_d  = go_16_goMux_data_onehotd[1];
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_d  = go_16_goMux_data_onehotd[2];
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_d  = go_16_goMux_data_onehotd[3];
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_d  = go_16_goMux_data_onehotd[4];
  assign go_16_goMux_data_r = (| (go_16_goMux_data_onehotd & {\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_r ,
                                                              \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_r ,
                                                              \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_r ,
                                                              \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_r ,
                                                              _25_r}));
  assign lizzieLet50_3_r = go_16_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0,Go) > (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf,Go) */
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_r ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_r  = ((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d [0]) || \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_r )
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_d ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_r  = (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0]);
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_d  = (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0] ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  :
                                                                       \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_r  && \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0]))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_r ) && (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0])))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1,Go) > (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf,Go) */
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_r ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_r  = ((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d [0]) || \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_r )
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_d ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_r  = (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0]);
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_d  = (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0] ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  :
                                                                       \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_r  && \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0]))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_1_argbuf_r ) && (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0])))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2,Go) > (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf,Go) */
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_r ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_r  = ((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d [0]) || \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_r )
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_d ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_r  = (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0]);
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_d  = (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0] ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  :
                                                                       \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_r  && \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0]))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_1_argbuf_r ) && (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0])))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3,Go) > (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf,Go) */
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d ;
  logic \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_r ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_r  = ((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d [0]) || \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_r )
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_d ;
  Go_t \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf ;
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_r  = (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0]);
  assign \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_d  = (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0] ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  :
                                                                       \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_r  && \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0]))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_1_argbuf_r ) && (! \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0])))
        \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int3_bufchan_d ;
  
  /* demux (Ty CTf'''''''''_f'''''''''_Int,
       Ty Pointer_QTree_Int) : (lizzieLet50_4,CTf'''''''''_f'''''''''_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos,Pointer_QTree_Int),
                                                                                                                       (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3,Pointer_QTree_Int),
                                                                                                                       (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2,Pointer_QTree_Int),
                                                                                                                       (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1,Pointer_QTree_Int),
                                                                                                                       (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet50_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet50_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                            srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                              srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                              srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                              srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                              srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_r ,
                                                                      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_r ,
                                                                      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_r ,
                                                                      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_r ,
                                                                      \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_r }));
  assign lizzieLet50_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0,Pointer_QTree_Int),
                         (es_1_2_destruct,Pointer_QTree_Int),
                         (es_2_3_destruct,Pointer_QTree_Int),
                         (es_3_4_destruct,Pointer_QTree_Int)] > (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int,QTree_Int) */
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_d [0],
                                                                                                                 es_1_2_destruct_d[0],
                                                                                                                 es_2_3_destruct_d[0],
                                                                                                                 es_3_4_destruct_d[0]}), \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_d , es_1_2_destruct_d, es_2_3_destruct_d, es_3_4_destruct_d);
  assign {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_r ,
          es_1_2_destruct_r,
          es_2_3_destruct_r,
          es_3_4_destruct_r} = {4 {(\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_r  && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int,QTree_Int) > (lizzieLet54_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_r ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_r  = ((! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d [0]) || \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                       1'd0};
    else
      if (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_r )
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_d ;
  QTree_Int_t \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_r  = (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet54_1_argbuf_d = (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf [0] ? \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf  :
                                   \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                         1'd0};
    else
      if ((lizzieLet54_1_argbuf_r && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf [0]))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                           1'd0};
      else if (((! lizzieLet54_1_argbuf_r) && (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf [0])))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_buf  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int0_1es_1_2_1es_2_3_1es_3_4_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Int,
      Dcon Lcall_f'''''''''_f'''''''''_Int0) : [(lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1,Pointer_QTree_Int),
                                                (es_2_2_destruct,Pointer_QTree_Int),
                                                (es_3_3_destruct,Pointer_QTree_Int),
                                                (sc_0_10_destruct,Pointer_CTf'''''''''_f'''''''''_Int)] > (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0,CTf'''''''''_f'''''''''_Int) */
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_d  = \Lcall_f'''''''''_f'''''''''_Int0_dc ((& {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_d [0],
                                                                                                                                                                  es_2_2_destruct_d[0],
                                                                                                                                                                  es_3_3_destruct_d[0],
                                                                                                                                                                  sc_0_10_destruct_d[0]}), \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_d , es_2_2_destruct_d, es_3_3_destruct_d, sc_0_10_destruct_d);
  assign {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_r ,
          es_2_2_destruct_r,
          es_3_3_destruct_r,
          sc_0_10_destruct_r} = {4 {(\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_r  && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0,CTf'''''''''_f'''''''''_Int) > (lizzieLet53_1_argbuf,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_r ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_r  = ((! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d [0]) || \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d  <= {115'd0,
                                                                                                                               1'd0};
    else
      if (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_r )
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_d ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_r  = (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0]);
  assign lizzieLet53_1_argbuf_d = (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0] ? \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  :
                                   \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= {115'd0,
                                                                                                                                 1'd0};
    else
      if ((lizzieLet53_1_argbuf_r && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0]))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= {115'd0,
                                                                                                                                   1'd0};
      else if (((! lizzieLet53_1_argbuf_r) && (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf [0])))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_buf  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int1_1es_2_2_1es_3_3_1sc_0_10_1Lcall_f'''''''''_f'''''''''_Int0_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Int,
      Dcon Lcall_f'''''''''_f'''''''''_Int1) : [(lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2,Pointer_QTree_Int),
                                                (es_3_2_destruct,Pointer_QTree_Int),
                                                (sc_0_9_destruct,Pointer_CTf'''''''''_f'''''''''_Int),
                                                (q1aey_2_destruct,Pointer_MaskQTree),
                                                (t1aeD_2_destruct,Pointer_QTree_Int)] > (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1,CTf'''''''''_f'''''''''_Int) */
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_d  = \Lcall_f'''''''''_f'''''''''_Int1_dc ((& {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_d [0],
                                                                                                                                                                           es_3_2_destruct_d[0],
                                                                                                                                                                           sc_0_9_destruct_d[0],
                                                                                                                                                                           q1aey_2_destruct_d[0],
                                                                                                                                                                           t1aeD_2_destruct_d[0]}), \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_d , es_3_2_destruct_d, sc_0_9_destruct_d, q1aey_2_destruct_d, t1aeD_2_destruct_d);
  assign {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_r ,
          es_3_2_destruct_r,
          sc_0_9_destruct_r,
          q1aey_2_destruct_r,
          t1aeD_2_destruct_r} = {5 {(\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_r  && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1,CTf'''''''''_f'''''''''_Int) > (lizzieLet52_1_argbuf,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_r ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_r  = ((! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d [0]) || \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d  <= {115'd0,
                                                                                                                                        1'd0};
    else
      if (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_r )
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_d ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_r  = (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0]);
  assign lizzieLet52_1_argbuf_d = (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0] ? \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  :
                                   \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                          1'd0};
    else
      if ((lizzieLet52_1_argbuf_r && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0]))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                            1'd0};
      else if (((! lizzieLet52_1_argbuf_r) && (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf [0])))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_buf  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int2_1es_3_2_1sc_0_9_1q1aey_2_1t1aeD_2_1Lcall_f'''''''''_f'''''''''_Int1_bufchan_d ;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Int,
      Dcon Lcall_f'''''''''_f'''''''''_Int2) : [(lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3,Pointer_QTree_Int),
                                                (sc_0_8_destruct,Pointer_CTf'''''''''_f'''''''''_Int),
                                                (q1aey_1_destruct,Pointer_MaskQTree),
                                                (t1aeD_1_destruct,Pointer_QTree_Int),
                                                (q2aez_1_destruct,Pointer_MaskQTree),
                                                (t2aeE_1_destruct,Pointer_QTree_Int)] > (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2,CTf'''''''''_f'''''''''_Int) */
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_d  = \Lcall_f'''''''''_f'''''''''_Int2_dc ((& {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_d [0],
                                                                                                                                                                                     sc_0_8_destruct_d[0],
                                                                                                                                                                                     q1aey_1_destruct_d[0],
                                                                                                                                                                                     t1aeD_1_destruct_d[0],
                                                                                                                                                                                     q2aez_1_destruct_d[0],
                                                                                                                                                                                     t2aeE_1_destruct_d[0]}), \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_d , sc_0_8_destruct_d, q1aey_1_destruct_d, t1aeD_1_destruct_d, q2aez_1_destruct_d, t2aeE_1_destruct_d);
  assign {\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_r ,
          sc_0_8_destruct_r,
          q1aey_1_destruct_r,
          t1aeD_1_destruct_r,
          q2aez_1_destruct_r,
          t2aeE_1_destruct_r} = {6 {(\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_r  && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2,CTf'''''''''_f'''''''''_Int) > (lizzieLet51_1_argbuf,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d ;
  logic \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_r ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_r  = ((! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d [0]) || \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d  <= {115'd0,
                                                                                                                                                  1'd0};
    else
      if (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_r )
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_d ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf ;
  assign \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_r  = (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0]);
  assign lizzieLet51_1_argbuf_d = (\lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0] ? \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  :
                                   \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                                    1'd0};
    else
      if ((lizzieLet51_1_argbuf_r && \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0]))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                                      1'd0};
      else if (((! lizzieLet51_1_argbuf_r) && (! \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf [0])))
        \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_buf  <= \lizzieLet50_4Lcall_f'''''''''_f'''''''''_Int3_1sc_0_8_1q1aey_1_1t1aeD_1_1q2aez_1_1t2aeE_1_1Lcall_f'''''''''_f'''''''''_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos,Pointer_QTree_Int) > [(lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                                 (lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted ;
  logic [1:0] \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_done ;
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d [16:1],
                                                                                 (\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d [0] && (! \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted [0]))};
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d [16:1],
                                                                                 (\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_d [0] && (! \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted [1]))};
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_done  = (\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted  | ({\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                         \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                     \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_r  = (& \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_emitted  <= (\lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_r  ? 2'd0 :
                                                                \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f'''''''''_f'''''''''_Int_goConst,Go) */
  assign \call_f'''''''''_f'''''''''_Int_goConst_d  = \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet50_4Lf'''''''''_f'''''''''_Intsbos_1_merge_merge_fork_1_r  = \call_f'''''''''_f'''''''''_Int_goConst_r ;
  
  /* destruct (Ty CTf'_f'_Int,
          Dcon Lcall_f'_f'_Int0) : (lizzieLet55_1Lcall_f'_f'_Int0,CTf'_f'_Int) > [(es_5_2_destruct,Pointer_QTree_Int),
                                                                                  (es_6_4_destruct,Pointer_QTree_Int),
                                                                                  (es_7_3_destruct,Pointer_QTree_Int),
                                                                                  (sc_0_15_destruct,Pointer_CTf'_f'_Int)] */
  logic [3:0] \lizzieLet55_1Lcall_f'_f'_Int0_emitted ;
  logic [3:0] \lizzieLet55_1Lcall_f'_f'_Int0_done ;
  assign es_5_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int0_d [19:4],
                              (\lizzieLet55_1Lcall_f'_f'_Int0_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int0_emitted [0]))};
  assign es_6_4_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int0_d [35:20],
                              (\lizzieLet55_1Lcall_f'_f'_Int0_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int0_emitted [1]))};
  assign es_7_3_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int0_d [51:36],
                              (\lizzieLet55_1Lcall_f'_f'_Int0_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int0_emitted [2]))};
  assign sc_0_15_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int0_d [67:52],
                               (\lizzieLet55_1Lcall_f'_f'_Int0_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int0_emitted [3]))};
  assign \lizzieLet55_1Lcall_f'_f'_Int0_done  = (\lizzieLet55_1Lcall_f'_f'_Int0_emitted  | ({sc_0_15_destruct_d[0],
                                                                                             es_7_3_destruct_d[0],
                                                                                             es_6_4_destruct_d[0],
                                                                                             es_5_2_destruct_d[0]} & {sc_0_15_destruct_r,
                                                                                                                      es_7_3_destruct_r,
                                                                                                                      es_6_4_destruct_r,
                                                                                                                      es_5_2_destruct_r}));
  assign \lizzieLet55_1Lcall_f'_f'_Int0_r  = (& \lizzieLet55_1Lcall_f'_f'_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_1Lcall_f'_f'_Int0_emitted  <= 4'd0;
    else
      \lizzieLet55_1Lcall_f'_f'_Int0_emitted  <= (\lizzieLet55_1Lcall_f'_f'_Int0_r  ? 4'd0 :
                                                  \lizzieLet55_1Lcall_f'_f'_Int0_done );
  
  /* destruct (Ty CTf'_f'_Int,
          Dcon Lcall_f'_f'_Int1) : (lizzieLet55_1Lcall_f'_f'_Int1,CTf'_f'_Int) > [(es_6_3_destruct,Pointer_QTree_Int),
                                                                                  (es_7_2_destruct,Pointer_QTree_Int),
                                                                                  (sc_0_14_destruct,Pointer_CTf'_f'_Int),
                                                                                  (q1aeR_3_destruct,Pointer_QTree_Int),
                                                                                  (t1aeW_3_destruct,Pointer_QTree_Int),
                                                                                  (is_zaeJ_4_destruct,MyDTInt_Bool),
                                                                                  (op_addaeK_4_destruct,MyDTInt_Int_Int)] */
  logic [6:0] \lizzieLet55_1Lcall_f'_f'_Int1_emitted ;
  logic [6:0] \lizzieLet55_1Lcall_f'_f'_Int1_done ;
  assign es_6_3_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int1_d [19:4],
                              (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [0]))};
  assign es_7_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int1_d [35:20],
                              (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [1]))};
  assign sc_0_14_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int1_d [51:36],
                               (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [2]))};
  assign q1aeR_3_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int1_d [67:52],
                               (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [3]))};
  assign t1aeW_3_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int1_d [83:68],
                               (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [4]))};
  assign is_zaeJ_4_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [5]));
  assign op_addaeK_4_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int1_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int1_emitted [6]));
  assign \lizzieLet55_1Lcall_f'_f'_Int1_done  = (\lizzieLet55_1Lcall_f'_f'_Int1_emitted  | ({op_addaeK_4_destruct_d[0],
                                                                                             is_zaeJ_4_destruct_d[0],
                                                                                             t1aeW_3_destruct_d[0],
                                                                                             q1aeR_3_destruct_d[0],
                                                                                             sc_0_14_destruct_d[0],
                                                                                             es_7_2_destruct_d[0],
                                                                                             es_6_3_destruct_d[0]} & {op_addaeK_4_destruct_r,
                                                                                                                      is_zaeJ_4_destruct_r,
                                                                                                                      t1aeW_3_destruct_r,
                                                                                                                      q1aeR_3_destruct_r,
                                                                                                                      sc_0_14_destruct_r,
                                                                                                                      es_7_2_destruct_r,
                                                                                                                      es_6_3_destruct_r}));
  assign \lizzieLet55_1Lcall_f'_f'_Int1_r  = (& \lizzieLet55_1Lcall_f'_f'_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_1Lcall_f'_f'_Int1_emitted  <= 7'd0;
    else
      \lizzieLet55_1Lcall_f'_f'_Int1_emitted  <= (\lizzieLet55_1Lcall_f'_f'_Int1_r  ? 7'd0 :
                                                  \lizzieLet55_1Lcall_f'_f'_Int1_done );
  
  /* destruct (Ty CTf'_f'_Int,
          Dcon Lcall_f'_f'_Int2) : (lizzieLet55_1Lcall_f'_f'_Int2,CTf'_f'_Int) > [(es_7_1_destruct,Pointer_QTree_Int),
                                                                                  (sc_0_13_destruct,Pointer_CTf'_f'_Int),
                                                                                  (q1aeR_2_destruct,Pointer_QTree_Int),
                                                                                  (t1aeW_2_destruct,Pointer_QTree_Int),
                                                                                  (is_zaeJ_3_destruct,MyDTInt_Bool),
                                                                                  (op_addaeK_3_destruct,MyDTInt_Int_Int),
                                                                                  (q2aeS_2_destruct,Pointer_QTree_Int),
                                                                                  (t2aeX_2_destruct,Pointer_QTree_Int)] */
  logic [7:0] \lizzieLet55_1Lcall_f'_f'_Int2_emitted ;
  logic [7:0] \lizzieLet55_1Lcall_f'_f'_Int2_done ;
  assign es_7_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [19:4],
                              (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [0]))};
  assign sc_0_13_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [35:20],
                               (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [1]))};
  assign q1aeR_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [51:36],
                               (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [2]))};
  assign t1aeW_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [67:52],
                               (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [3]))};
  assign is_zaeJ_3_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [4]));
  assign op_addaeK_3_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [5]));
  assign q2aeS_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [83:68],
                               (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [6]))};
  assign t2aeX_2_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int2_d [99:84],
                               (\lizzieLet55_1Lcall_f'_f'_Int2_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int2_emitted [7]))};
  assign \lizzieLet55_1Lcall_f'_f'_Int2_done  = (\lizzieLet55_1Lcall_f'_f'_Int2_emitted  | ({t2aeX_2_destruct_d[0],
                                                                                             q2aeS_2_destruct_d[0],
                                                                                             op_addaeK_3_destruct_d[0],
                                                                                             is_zaeJ_3_destruct_d[0],
                                                                                             t1aeW_2_destruct_d[0],
                                                                                             q1aeR_2_destruct_d[0],
                                                                                             sc_0_13_destruct_d[0],
                                                                                             es_7_1_destruct_d[0]} & {t2aeX_2_destruct_r,
                                                                                                                      q2aeS_2_destruct_r,
                                                                                                                      op_addaeK_3_destruct_r,
                                                                                                                      is_zaeJ_3_destruct_r,
                                                                                                                      t1aeW_2_destruct_r,
                                                                                                                      q1aeR_2_destruct_r,
                                                                                                                      sc_0_13_destruct_r,
                                                                                                                      es_7_1_destruct_r}));
  assign \lizzieLet55_1Lcall_f'_f'_Int2_r  = (& \lizzieLet55_1Lcall_f'_f'_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_1Lcall_f'_f'_Int2_emitted  <= 8'd0;
    else
      \lizzieLet55_1Lcall_f'_f'_Int2_emitted  <= (\lizzieLet55_1Lcall_f'_f'_Int2_r  ? 8'd0 :
                                                  \lizzieLet55_1Lcall_f'_f'_Int2_done );
  
  /* destruct (Ty CTf'_f'_Int,
          Dcon Lcall_f'_f'_Int3) : (lizzieLet55_1Lcall_f'_f'_Int3,CTf'_f'_Int) > [(sc_0_12_destruct,Pointer_CTf'_f'_Int),
                                                                                  (q1aeR_1_destruct,Pointer_QTree_Int),
                                                                                  (t1aeW_1_destruct,Pointer_QTree_Int),
                                                                                  (is_zaeJ_2_destruct,MyDTInt_Bool),
                                                                                  (op_addaeK_2_destruct,MyDTInt_Int_Int),
                                                                                  (q2aeS_1_destruct,Pointer_QTree_Int),
                                                                                  (t2aeX_1_destruct,Pointer_QTree_Int),
                                                                                  (q3aeT_1_destruct,Pointer_QTree_Int),
                                                                                  (t3aeY_1_destruct,Pointer_QTree_Int)] */
  logic [8:0] \lizzieLet55_1Lcall_f'_f'_Int3_emitted ;
  logic [8:0] \lizzieLet55_1Lcall_f'_f'_Int3_done ;
  assign sc_0_12_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [19:4],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [0]))};
  assign q1aeR_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [35:20],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [1]))};
  assign t1aeW_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [51:36],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [2]))};
  assign is_zaeJ_2_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [3]));
  assign op_addaeK_2_destruct_d = (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [4]));
  assign q2aeS_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [67:52],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [5]))};
  assign t2aeX_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [83:68],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [6]))};
  assign q3aeT_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [99:84],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [7]))};
  assign t3aeY_1_destruct_d = {\lizzieLet55_1Lcall_f'_f'_Int3_d [115:100],
                               (\lizzieLet55_1Lcall_f'_f'_Int3_d [0] && (! \lizzieLet55_1Lcall_f'_f'_Int3_emitted [8]))};
  assign \lizzieLet55_1Lcall_f'_f'_Int3_done  = (\lizzieLet55_1Lcall_f'_f'_Int3_emitted  | ({t3aeY_1_destruct_d[0],
                                                                                             q3aeT_1_destruct_d[0],
                                                                                             t2aeX_1_destruct_d[0],
                                                                                             q2aeS_1_destruct_d[0],
                                                                                             op_addaeK_2_destruct_d[0],
                                                                                             is_zaeJ_2_destruct_d[0],
                                                                                             t1aeW_1_destruct_d[0],
                                                                                             q1aeR_1_destruct_d[0],
                                                                                             sc_0_12_destruct_d[0]} & {t3aeY_1_destruct_r,
                                                                                                                       q3aeT_1_destruct_r,
                                                                                                                       t2aeX_1_destruct_r,
                                                                                                                       q2aeS_1_destruct_r,
                                                                                                                       op_addaeK_2_destruct_r,
                                                                                                                       is_zaeJ_2_destruct_r,
                                                                                                                       t1aeW_1_destruct_r,
                                                                                                                       q1aeR_1_destruct_r,
                                                                                                                       sc_0_12_destruct_r}));
  assign \lizzieLet55_1Lcall_f'_f'_Int3_r  = (& \lizzieLet55_1Lcall_f'_f'_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_1Lcall_f'_f'_Int3_emitted  <= 9'd0;
    else
      \lizzieLet55_1Lcall_f'_f'_Int3_emitted  <= (\lizzieLet55_1Lcall_f'_f'_Int3_r  ? 9'd0 :
                                                  \lizzieLet55_1Lcall_f'_f'_Int3_done );
  
  /* demux (Ty CTf'_f'_Int,
       Ty CTf'_f'_Int) : (lizzieLet55_2,CTf'_f'_Int) (lizzieLet55_1,CTf'_f'_Int) > [(_24,CTf'_f'_Int),
                                                                                    (lizzieLet55_1Lcall_f'_f'_Int3,CTf'_f'_Int),
                                                                                    (lizzieLet55_1Lcall_f'_f'_Int2,CTf'_f'_Int),
                                                                                    (lizzieLet55_1Lcall_f'_f'_Int1,CTf'_f'_Int),
                                                                                    (lizzieLet55_1Lcall_f'_f'_Int0,CTf'_f'_Int)] */
  logic [4:0] lizzieLet55_1_onehotd;
  always_comb
    if ((lizzieLet55_2_d[0] && lizzieLet55_1_d[0]))
      unique case (lizzieLet55_2_d[3:1])
        3'd0: lizzieLet55_1_onehotd = 5'd1;
        3'd1: lizzieLet55_1_onehotd = 5'd2;
        3'd2: lizzieLet55_1_onehotd = 5'd4;
        3'd3: lizzieLet55_1_onehotd = 5'd8;
        3'd4: lizzieLet55_1_onehotd = 5'd16;
        default: lizzieLet55_1_onehotd = 5'd0;
      endcase
    else lizzieLet55_1_onehotd = 5'd0;
  assign _24_d = {lizzieLet55_1_d[115:1], lizzieLet55_1_onehotd[0]};
  assign \lizzieLet55_1Lcall_f'_f'_Int3_d  = {lizzieLet55_1_d[115:1],
                                              lizzieLet55_1_onehotd[1]};
  assign \lizzieLet55_1Lcall_f'_f'_Int2_d  = {lizzieLet55_1_d[115:1],
                                              lizzieLet55_1_onehotd[2]};
  assign \lizzieLet55_1Lcall_f'_f'_Int1_d  = {lizzieLet55_1_d[115:1],
                                              lizzieLet55_1_onehotd[3]};
  assign \lizzieLet55_1Lcall_f'_f'_Int0_d  = {lizzieLet55_1_d[115:1],
                                              lizzieLet55_1_onehotd[4]};
  assign lizzieLet55_1_r = (| (lizzieLet55_1_onehotd & {\lizzieLet55_1Lcall_f'_f'_Int0_r ,
                                                        \lizzieLet55_1Lcall_f'_f'_Int1_r ,
                                                        \lizzieLet55_1Lcall_f'_f'_Int2_r ,
                                                        \lizzieLet55_1Lcall_f'_f'_Int3_r ,
                                                        _24_r}));
  assign lizzieLet55_2_r = lizzieLet55_1_r;
  
  /* demux (Ty CTf'_f'_Int,
       Ty Go) : (lizzieLet55_3,CTf'_f'_Int) (go_17_goMux_data,Go) > [(_23,Go),
                                                                     (lizzieLet55_3Lcall_f'_f'_Int3,Go),
                                                                     (lizzieLet55_3Lcall_f'_f'_Int2,Go),
                                                                     (lizzieLet55_3Lcall_f'_f'_Int1,Go),
                                                                     (lizzieLet55_3Lcall_f'_f'_Int0,Go)] */
  logic [4:0] go_17_goMux_data_onehotd;
  always_comb
    if ((lizzieLet55_3_d[0] && go_17_goMux_data_d[0]))
      unique case (lizzieLet55_3_d[3:1])
        3'd0: go_17_goMux_data_onehotd = 5'd1;
        3'd1: go_17_goMux_data_onehotd = 5'd2;
        3'd2: go_17_goMux_data_onehotd = 5'd4;
        3'd3: go_17_goMux_data_onehotd = 5'd8;
        3'd4: go_17_goMux_data_onehotd = 5'd16;
        default: go_17_goMux_data_onehotd = 5'd0;
      endcase
    else go_17_goMux_data_onehotd = 5'd0;
  assign _23_d = go_17_goMux_data_onehotd[0];
  assign \lizzieLet55_3Lcall_f'_f'_Int3_d  = go_17_goMux_data_onehotd[1];
  assign \lizzieLet55_3Lcall_f'_f'_Int2_d  = go_17_goMux_data_onehotd[2];
  assign \lizzieLet55_3Lcall_f'_f'_Int1_d  = go_17_goMux_data_onehotd[3];
  assign \lizzieLet55_3Lcall_f'_f'_Int0_d  = go_17_goMux_data_onehotd[4];
  assign go_17_goMux_data_r = (| (go_17_goMux_data_onehotd & {\lizzieLet55_3Lcall_f'_f'_Int0_r ,
                                                              \lizzieLet55_3Lcall_f'_f'_Int1_r ,
                                                              \lizzieLet55_3Lcall_f'_f'_Int2_r ,
                                                              \lizzieLet55_3Lcall_f'_f'_Int3_r ,
                                                              _23_r}));
  assign lizzieLet55_3_r = go_17_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet55_3Lcall_f'_f'_Int0,Go) > (lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf,Go) */
  Go_t \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_r ;
  assign \lizzieLet55_3Lcall_f'_f'_Int0_r  = ((! \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d [0]) || \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet55_3Lcall_f'_f'_Int0_r )
        \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d  <= \lizzieLet55_3Lcall_f'_f'_Int0_d ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf ;
  assign \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_r  = (! \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf [0]);
  assign \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_d  = (\lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf [0] ? \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf  :
                                                       \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_r  && \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf [0]))
        \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet55_3Lcall_f'_f'_Int0_1_argbuf_r ) && (! \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf [0])))
        \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_buf  <= \lizzieLet55_3Lcall_f'_f'_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet55_3Lcall_f'_f'_Int1,Go) > (lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf,Go) */
  Go_t \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_r ;
  assign \lizzieLet55_3Lcall_f'_f'_Int1_r  = ((! \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d [0]) || \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet55_3Lcall_f'_f'_Int1_r )
        \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d  <= \lizzieLet55_3Lcall_f'_f'_Int1_d ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf ;
  assign \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_r  = (! \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf [0]);
  assign \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_d  = (\lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf [0] ? \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf  :
                                                       \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_r  && \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf [0]))
        \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet55_3Lcall_f'_f'_Int1_1_argbuf_r ) && (! \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf [0])))
        \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_buf  <= \lizzieLet55_3Lcall_f'_f'_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet55_3Lcall_f'_f'_Int2,Go) > (lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf,Go) */
  Go_t \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_r ;
  assign \lizzieLet55_3Lcall_f'_f'_Int2_r  = ((! \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d [0]) || \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet55_3Lcall_f'_f'_Int2_r )
        \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d  <= \lizzieLet55_3Lcall_f'_f'_Int2_d ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf ;
  assign \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_r  = (! \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf [0]);
  assign \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_d  = (\lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf [0] ? \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf  :
                                                       \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_r  && \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf [0]))
        \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet55_3Lcall_f'_f'_Int2_1_argbuf_r ) && (! \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf [0])))
        \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_buf  <= \lizzieLet55_3Lcall_f'_f'_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet55_3Lcall_f'_f'_Int3,Go) > (lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf,Go) */
  Go_t \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d ;
  logic \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_r ;
  assign \lizzieLet55_3Lcall_f'_f'_Int3_r  = ((! \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d [0]) || \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet55_3Lcall_f'_f'_Int3_r )
        \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d  <= \lizzieLet55_3Lcall_f'_f'_Int3_d ;
  Go_t \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf ;
  assign \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_r  = (! \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf [0]);
  assign \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_d  = (\lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf [0] ? \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf  :
                                                       \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_r  && \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf [0]))
        \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet55_3Lcall_f'_f'_Int3_1_argbuf_r ) && (! \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf [0])))
        \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_buf  <= \lizzieLet55_3Lcall_f'_f'_Int3_bufchan_d ;
  
  /* demux (Ty CTf'_f'_Int,
       Ty Pointer_QTree_Int) : (lizzieLet55_4,CTf'_f'_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet55_4Lf'_f'_Intsbos,Pointer_QTree_Int),
                                                                                                       (lizzieLet55_4Lcall_f'_f'_Int3,Pointer_QTree_Int),
                                                                                                       (lizzieLet55_4Lcall_f'_f'_Int2,Pointer_QTree_Int),
                                                                                                       (lizzieLet55_4Lcall_f'_f'_Int1,Pointer_QTree_Int),
                                                                                                       (lizzieLet55_4Lcall_f'_f'_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet55_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet55_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet55_4Lf'_f'_Intsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                            srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet55_4Lcall_f'_f'_Int3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet55_4Lcall_f'_f'_Int2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet55_4Lcall_f'_f'_Int1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet55_4Lcall_f'_f'_Int0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                              srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet55_4Lcall_f'_f'_Int0_r ,
                                                                      \lizzieLet55_4Lcall_f'_f'_Int1_r ,
                                                                      \lizzieLet55_4Lcall_f'_f'_Int2_r ,
                                                                      \lizzieLet55_4Lcall_f'_f'_Int3_r ,
                                                                      \lizzieLet55_4Lf'_f'_Intsbos_r }));
  assign lizzieLet55_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet55_4Lcall_f'_f'_Int0,Pointer_QTree_Int),
                         (es_5_2_destruct,Pointer_QTree_Int),
                         (es_6_4_destruct,Pointer_QTree_Int),
                         (es_7_3_destruct,Pointer_QTree_Int)] > (lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int,QTree_Int) */
  assign \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet55_4Lcall_f'_f'_Int0_d [0],
                                                                                                 es_5_2_destruct_d[0],
                                                                                                 es_6_4_destruct_d[0],
                                                                                                 es_7_3_destruct_d[0]}), \lizzieLet55_4Lcall_f'_f'_Int0_d , es_5_2_destruct_d, es_6_4_destruct_d, es_7_3_destruct_d);
  assign {\lizzieLet55_4Lcall_f'_f'_Int0_r ,
          es_5_2_destruct_r,
          es_6_4_destruct_r,
          es_7_3_destruct_r} = {4 {(\lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r  && \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int,QTree_Int) > (lizzieLet59_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r ;
  assign \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r  = ((! \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d [0]) || \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                       1'd0};
    else
      if (\lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_r )
        \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d  <= \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_d ;
  QTree_Int_t \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf ;
  assign \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_r  = (! \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet59_1_argbuf_d = (\lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0] ? \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  :
                                   \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet59_1_argbuf_r && \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0]))
        \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                           1'd0};
      else if (((! lizzieLet59_1_argbuf_r) && (! \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf [0])))
        \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_buf  <= \lizzieLet55_4Lcall_f'_f'_Int0_1es_5_2_1es_6_4_1es_7_3_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int,
      Dcon Lcall_f'_f'_Int0) : [(lizzieLet55_4Lcall_f'_f'_Int1,Pointer_QTree_Int),
                                (es_6_3_destruct,Pointer_QTree_Int),
                                (es_7_2_destruct,Pointer_QTree_Int),
                                (sc_0_14_destruct,Pointer_CTf'_f'_Int)] > (lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0,CTf'_f'_Int) */
  assign \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_d  = \Lcall_f'_f'_Int0_dc ((& {\lizzieLet55_4Lcall_f'_f'_Int1_d [0],
                                                                                                                  es_6_3_destruct_d[0],
                                                                                                                  es_7_2_destruct_d[0],
                                                                                                                  sc_0_14_destruct_d[0]}), \lizzieLet55_4Lcall_f'_f'_Int1_d , es_6_3_destruct_d, es_7_2_destruct_d, sc_0_14_destruct_d);
  assign {\lizzieLet55_4Lcall_f'_f'_Int1_r ,
          es_6_3_destruct_r,
          es_7_2_destruct_r,
          sc_0_14_destruct_r} = {4 {(\lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_r  && \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_d [0])}};
  
  /* buf (Ty CTf'_f'_Int) : (lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0,CTf'_f'_Int) > (lizzieLet58_1_argbuf,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_r ;
  assign \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_r  = ((! \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d [0]) || \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d  <= {115'd0,
                                                                                               1'd0};
    else
      if (\lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_r )
        \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d  <= \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_d ;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf ;
  assign \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_r  = (! \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf [0]);
  assign lizzieLet58_1_argbuf_d = (\lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf [0] ? \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf  :
                                   \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf  <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet58_1_argbuf_r && \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf [0]))
        \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf  <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet58_1_argbuf_r) && (! \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf [0])))
        \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_buf  <= \lizzieLet55_4Lcall_f'_f'_Int1_1es_6_3_1es_7_2_1sc_0_14_1Lcall_f'_f'_Int0_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int,
      Dcon Lcall_f'_f'_Int1) : [(lizzieLet55_4Lcall_f'_f'_Int2,Pointer_QTree_Int),
                                (es_7_1_destruct,Pointer_QTree_Int),
                                (sc_0_13_destruct,Pointer_CTf'_f'_Int),
                                (q1aeR_2_destruct,Pointer_QTree_Int),
                                (t1aeW_2_destruct,Pointer_QTree_Int),
                                (is_zaeJ_3_1,MyDTInt_Bool),
                                (op_addaeK_3_1,MyDTInt_Int_Int)] > (lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1,CTf'_f'_Int) */
  assign \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_d  = \Lcall_f'_f'_Int1_dc ((& {\lizzieLet55_4Lcall_f'_f'_Int2_d [0],
                                                                                                                                                    es_7_1_destruct_d[0],
                                                                                                                                                    sc_0_13_destruct_d[0],
                                                                                                                                                    q1aeR_2_destruct_d[0],
                                                                                                                                                    t1aeW_2_destruct_d[0],
                                                                                                                                                    is_zaeJ_3_1_d[0],
                                                                                                                                                    op_addaeK_3_1_d[0]}), \lizzieLet55_4Lcall_f'_f'_Int2_d , es_7_1_destruct_d, sc_0_13_destruct_d, q1aeR_2_destruct_d, t1aeW_2_destruct_d, is_zaeJ_3_1_d, op_addaeK_3_1_d);
  assign {\lizzieLet55_4Lcall_f'_f'_Int2_r ,
          es_7_1_destruct_r,
          sc_0_13_destruct_r,
          q1aeR_2_destruct_r,
          t1aeW_2_destruct_r,
          is_zaeJ_3_1_r,
          op_addaeK_3_1_r} = {7 {(\lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_r  && \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_d [0])}};
  
  /* buf (Ty CTf'_f'_Int) : (lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1,CTf'_f'_Int) > (lizzieLet57_1_argbuf,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_r ;
  assign \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_r  = ((! \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d [0]) || \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d  <= {115'd0,
                                                                                                                                 1'd0};
    else
      if (\lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_r )
        \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d  <= \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_d ;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf ;
  assign \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_r  = (! \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf [0]);
  assign lizzieLet57_1_argbuf_d = (\lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf [0] ? \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf  :
                                   \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                   1'd0};
    else
      if ((lizzieLet57_1_argbuf_r && \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf [0]))
        \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf  <= {115'd0,
                                                                                                                                     1'd0};
      else if (((! lizzieLet57_1_argbuf_r) && (! \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf [0])))
        \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_buf  <= \lizzieLet55_4Lcall_f'_f'_Int2_1es_7_1_1sc_0_13_1q1aeR_2_1t1aeW_2_1is_zaeJ_3_1op_addaeK_3_1Lcall_f'_f'_Int1_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int,
      Dcon Lcall_f'_f'_Int2) : [(lizzieLet55_4Lcall_f'_f'_Int3,Pointer_QTree_Int),
                                (sc_0_12_destruct,Pointer_CTf'_f'_Int),
                                (q1aeR_1_destruct,Pointer_QTree_Int),
                                (t1aeW_1_destruct,Pointer_QTree_Int),
                                (is_zaeJ_2_1,MyDTInt_Bool),
                                (op_addaeK_2_1,MyDTInt_Int_Int),
                                (q2aeS_1_destruct,Pointer_QTree_Int),
                                (t2aeX_1_destruct,Pointer_QTree_Int)] > (lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2,CTf'_f'_Int) */
  assign \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_d  = \Lcall_f'_f'_Int2_dc ((& {\lizzieLet55_4Lcall_f'_f'_Int3_d [0],
                                                                                                                                                              sc_0_12_destruct_d[0],
                                                                                                                                                              q1aeR_1_destruct_d[0],
                                                                                                                                                              t1aeW_1_destruct_d[0],
                                                                                                                                                              is_zaeJ_2_1_d[0],
                                                                                                                                                              op_addaeK_2_1_d[0],
                                                                                                                                                              q2aeS_1_destruct_d[0],
                                                                                                                                                              t2aeX_1_destruct_d[0]}), \lizzieLet55_4Lcall_f'_f'_Int3_d , sc_0_12_destruct_d, q1aeR_1_destruct_d, t1aeW_1_destruct_d, is_zaeJ_2_1_d, op_addaeK_2_1_d, q2aeS_1_destruct_d, t2aeX_1_destruct_d);
  assign {\lizzieLet55_4Lcall_f'_f'_Int3_r ,
          sc_0_12_destruct_r,
          q1aeR_1_destruct_r,
          t1aeW_1_destruct_r,
          is_zaeJ_2_1_r,
          op_addaeK_2_1_r,
          q2aeS_1_destruct_r,
          t2aeX_1_destruct_r} = {8 {(\lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_r  && \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_d [0])}};
  
  /* buf (Ty CTf'_f'_Int) : (lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2,CTf'_f'_Int) > (lizzieLet56_1_argbuf,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d ;
  logic \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_r ;
  assign \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_r  = ((! \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d [0]) || \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d  <= {115'd0,
                                                                                                                                           1'd0};
    else
      if (\lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_r )
        \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d  <= \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_d ;
  \CTf'_f'_Int_t  \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf ;
  assign \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_r  = (! \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf [0]);
  assign lizzieLet56_1_argbuf_d = (\lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf [0] ? \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf  :
                                   \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                             1'd0};
    else
      if ((lizzieLet56_1_argbuf_r && \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf [0]))
        \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf  <= {115'd0,
                                                                                                                                               1'd0};
      else if (((! lizzieLet56_1_argbuf_r) && (! \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf [0])))
        \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_buf  <= \lizzieLet55_4Lcall_f'_f'_Int3_1sc_0_12_1q1aeR_1_1t1aeW_1_1is_zaeJ_2_1op_addaeK_2_1q2aeS_1_1t2aeX_1_1Lcall_f'_f'_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet55_4Lf'_f'_Intsbos,Pointer_QTree_Int) > [(lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                 (lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet55_4Lf'_f'_Intsbos_emitted ;
  logic [1:0] \lizzieLet55_4Lf'_f'_Intsbos_done ;
  assign \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet55_4Lf'_f'_Intsbos_d [16:1],
                                                                 (\lizzieLet55_4Lf'_f'_Intsbos_d [0] && (! \lizzieLet55_4Lf'_f'_Intsbos_emitted [0]))};
  assign \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet55_4Lf'_f'_Intsbos_d [16:1],
                                                                 (\lizzieLet55_4Lf'_f'_Intsbos_d [0] && (! \lizzieLet55_4Lf'_f'_Intsbos_emitted [1]))};
  assign \lizzieLet55_4Lf'_f'_Intsbos_done  = (\lizzieLet55_4Lf'_f'_Intsbos_emitted  | ({\lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                         \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                     \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet55_4Lf'_f'_Intsbos_r  = (& \lizzieLet55_4Lf'_f'_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \lizzieLet55_4Lf'_f'_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet55_4Lf'_f'_Intsbos_emitted  <= (\lizzieLet55_4Lf'_f'_Intsbos_r  ? 2'd0 :
                                                \lizzieLet55_4Lf'_f'_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f'_f'_Int_goConst,Go) */
  assign \call_f'_f'_Int_goConst_d  = \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_1_r  = \call_f'_f'_Int_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (f'_f'_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_r )
        \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Int_t \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \f'_f'_Int_resbuf_d  = (\lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf  :
                                 \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((\f'_f'_Int_resbuf_r  && \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! \f'_f'_Int_resbuf_r ) && (! \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet55_4Lf'_f'_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int0) : (lizzieLet60_1Lcall_f_f_Int0,CTf_f_Int) > [(es_12_destruct,Pointer_QTree_Int),
                                                                            (es_13_1_destruct,Pointer_QTree_Int),
                                                                            (es_14_2_destruct,Pointer_QTree_Int),
                                                                            (sc_0_19_destruct,Pointer_CTf_f_Int)] */
  logic [3:0] lizzieLet60_1Lcall_f_f_Int0_emitted;
  logic [3:0] lizzieLet60_1Lcall_f_f_Int0_done;
  assign es_12_destruct_d = {lizzieLet60_1Lcall_f_f_Int0_d[19:4],
                             (lizzieLet60_1Lcall_f_f_Int0_d[0] && (! lizzieLet60_1Lcall_f_f_Int0_emitted[0]))};
  assign es_13_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int0_d[35:20],
                               (lizzieLet60_1Lcall_f_f_Int0_d[0] && (! lizzieLet60_1Lcall_f_f_Int0_emitted[1]))};
  assign es_14_2_destruct_d = {lizzieLet60_1Lcall_f_f_Int0_d[51:36],
                               (lizzieLet60_1Lcall_f_f_Int0_d[0] && (! lizzieLet60_1Lcall_f_f_Int0_emitted[2]))};
  assign sc_0_19_destruct_d = {lizzieLet60_1Lcall_f_f_Int0_d[67:52],
                               (lizzieLet60_1Lcall_f_f_Int0_d[0] && (! lizzieLet60_1Lcall_f_f_Int0_emitted[3]))};
  assign lizzieLet60_1Lcall_f_f_Int0_done = (lizzieLet60_1Lcall_f_f_Int0_emitted | ({sc_0_19_destruct_d[0],
                                                                                     es_14_2_destruct_d[0],
                                                                                     es_13_1_destruct_d[0],
                                                                                     es_12_destruct_d[0]} & {sc_0_19_destruct_r,
                                                                                                             es_14_2_destruct_r,
                                                                                                             es_13_1_destruct_r,
                                                                                                             es_12_destruct_r}));
  assign lizzieLet60_1Lcall_f_f_Int0_r = (& lizzieLet60_1Lcall_f_f_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f_f_Int0_emitted <= 4'd0;
    else
      lizzieLet60_1Lcall_f_f_Int0_emitted <= (lizzieLet60_1Lcall_f_f_Int0_r ? 4'd0 :
                                              lizzieLet60_1Lcall_f_f_Int0_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int1) : (lizzieLet60_1Lcall_f_f_Int1,CTf_f_Int) > [(es_13_destruct,Pointer_QTree_Int),
                                                                            (es_14_1_destruct,Pointer_QTree_Int),
                                                                            (sc_0_18_destruct,Pointer_CTf_f_Int),
                                                                            (q1ae8_3_destruct,Pointer_MaskQTree),
                                                                            (q1'aen_3_destruct,Pointer_QTree_Int),
                                                                            (t1aes_3_destruct,Pointer_QTree_Int),
                                                                            (is_zae6_4_destruct,MyDTInt_Bool),
                                                                            (op_addae7_4_destruct,MyDTInt_Int_Int)] */
  logic [7:0] lizzieLet60_1Lcall_f_f_Int1_emitted;
  logic [7:0] lizzieLet60_1Lcall_f_f_Int1_done;
  assign es_13_destruct_d = {lizzieLet60_1Lcall_f_f_Int1_d[19:4],
                             (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[0]))};
  assign es_14_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int1_d[35:20],
                               (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[1]))};
  assign sc_0_18_destruct_d = {lizzieLet60_1Lcall_f_f_Int1_d[51:36],
                               (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[2]))};
  assign q1ae8_3_destruct_d = {lizzieLet60_1Lcall_f_f_Int1_d[67:52],
                               (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[3]))};
  assign \q1'aen_3_destruct_d  = {lizzieLet60_1Lcall_f_f_Int1_d[83:68],
                                  (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[4]))};
  assign t1aes_3_destruct_d = {lizzieLet60_1Lcall_f_f_Int1_d[99:84],
                               (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[5]))};
  assign is_zae6_4_destruct_d = (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[6]));
  assign op_addae7_4_destruct_d = (lizzieLet60_1Lcall_f_f_Int1_d[0] && (! lizzieLet60_1Lcall_f_f_Int1_emitted[7]));
  assign lizzieLet60_1Lcall_f_f_Int1_done = (lizzieLet60_1Lcall_f_f_Int1_emitted | ({op_addae7_4_destruct_d[0],
                                                                                     is_zae6_4_destruct_d[0],
                                                                                     t1aes_3_destruct_d[0],
                                                                                     \q1'aen_3_destruct_d [0],
                                                                                     q1ae8_3_destruct_d[0],
                                                                                     sc_0_18_destruct_d[0],
                                                                                     es_14_1_destruct_d[0],
                                                                                     es_13_destruct_d[0]} & {op_addae7_4_destruct_r,
                                                                                                             is_zae6_4_destruct_r,
                                                                                                             t1aes_3_destruct_r,
                                                                                                             \q1'aen_3_destruct_r ,
                                                                                                             q1ae8_3_destruct_r,
                                                                                                             sc_0_18_destruct_r,
                                                                                                             es_14_1_destruct_r,
                                                                                                             es_13_destruct_r}));
  assign lizzieLet60_1Lcall_f_f_Int1_r = (& lizzieLet60_1Lcall_f_f_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f_f_Int1_emitted <= 8'd0;
    else
      lizzieLet60_1Lcall_f_f_Int1_emitted <= (lizzieLet60_1Lcall_f_f_Int1_r ? 8'd0 :
                                              lizzieLet60_1Lcall_f_f_Int1_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int2) : (lizzieLet60_1Lcall_f_f_Int2,CTf_f_Int) > [(es_14_destruct,Pointer_QTree_Int),
                                                                            (sc_0_17_destruct,Pointer_CTf_f_Int),
                                                                            (q1ae8_2_destruct,Pointer_MaskQTree),
                                                                            (q1'aen_2_destruct,Pointer_QTree_Int),
                                                                            (t1aes_2_destruct,Pointer_QTree_Int),
                                                                            (is_zae6_3_destruct,MyDTInt_Bool),
                                                                            (op_addae7_3_destruct,MyDTInt_Int_Int),
                                                                            (q2ae9_2_destruct,Pointer_MaskQTree),
                                                                            (q2'aeo_2_destruct,Pointer_QTree_Int),
                                                                            (t2aet_2_destruct,Pointer_QTree_Int)] */
  logic [9:0] lizzieLet60_1Lcall_f_f_Int2_emitted;
  logic [9:0] lizzieLet60_1Lcall_f_f_Int2_done;
  assign es_14_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[19:4],
                             (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[0]))};
  assign sc_0_17_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[35:20],
                               (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[1]))};
  assign q1ae8_2_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[51:36],
                               (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[2]))};
  assign \q1'aen_2_destruct_d  = {lizzieLet60_1Lcall_f_f_Int2_d[67:52],
                                  (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[3]))};
  assign t1aes_2_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[83:68],
                               (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[4]))};
  assign is_zae6_3_destruct_d = (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[5]));
  assign op_addae7_3_destruct_d = (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[6]));
  assign q2ae9_2_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[99:84],
                               (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[7]))};
  assign \q2'aeo_2_destruct_d  = {lizzieLet60_1Lcall_f_f_Int2_d[115:100],
                                  (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[8]))};
  assign t2aet_2_destruct_d = {lizzieLet60_1Lcall_f_f_Int2_d[131:116],
                               (lizzieLet60_1Lcall_f_f_Int2_d[0] && (! lizzieLet60_1Lcall_f_f_Int2_emitted[9]))};
  assign lizzieLet60_1Lcall_f_f_Int2_done = (lizzieLet60_1Lcall_f_f_Int2_emitted | ({t2aet_2_destruct_d[0],
                                                                                     \q2'aeo_2_destruct_d [0],
                                                                                     q2ae9_2_destruct_d[0],
                                                                                     op_addae7_3_destruct_d[0],
                                                                                     is_zae6_3_destruct_d[0],
                                                                                     t1aes_2_destruct_d[0],
                                                                                     \q1'aen_2_destruct_d [0],
                                                                                     q1ae8_2_destruct_d[0],
                                                                                     sc_0_17_destruct_d[0],
                                                                                     es_14_destruct_d[0]} & {t2aet_2_destruct_r,
                                                                                                             \q2'aeo_2_destruct_r ,
                                                                                                             q2ae9_2_destruct_r,
                                                                                                             op_addae7_3_destruct_r,
                                                                                                             is_zae6_3_destruct_r,
                                                                                                             t1aes_2_destruct_r,
                                                                                                             \q1'aen_2_destruct_r ,
                                                                                                             q1ae8_2_destruct_r,
                                                                                                             sc_0_17_destruct_r,
                                                                                                             es_14_destruct_r}));
  assign lizzieLet60_1Lcall_f_f_Int2_r = (& lizzieLet60_1Lcall_f_f_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f_f_Int2_emitted <= 10'd0;
    else
      lizzieLet60_1Lcall_f_f_Int2_emitted <= (lizzieLet60_1Lcall_f_f_Int2_r ? 10'd0 :
                                              lizzieLet60_1Lcall_f_f_Int2_done);
  
  /* destruct (Ty CTf_f_Int,
          Dcon Lcall_f_f_Int3) : (lizzieLet60_1Lcall_f_f_Int3,CTf_f_Int) > [(sc_0_16_destruct,Pointer_CTf_f_Int),
                                                                            (q1ae8_1_destruct,Pointer_MaskQTree),
                                                                            (q1'aen_1_destruct,Pointer_QTree_Int),
                                                                            (t1aes_1_destruct,Pointer_QTree_Int),
                                                                            (is_zae6_2_destruct,MyDTInt_Bool),
                                                                            (op_addae7_2_destruct,MyDTInt_Int_Int),
                                                                            (q2ae9_1_destruct,Pointer_MaskQTree),
                                                                            (q2'aeo_1_destruct,Pointer_QTree_Int),
                                                                            (t2aet_1_destruct,Pointer_QTree_Int),
                                                                            (q3aea_1_destruct,Pointer_MaskQTree),
                                                                            (q3'aep_1_destruct,Pointer_QTree_Int),
                                                                            (t3aeu_1_destruct,Pointer_QTree_Int)] */
  logic [11:0] lizzieLet60_1Lcall_f_f_Int3_emitted;
  logic [11:0] lizzieLet60_1Lcall_f_f_Int3_done;
  assign sc_0_16_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[19:4],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[0]))};
  assign q1ae8_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[35:20],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[1]))};
  assign \q1'aen_1_destruct_d  = {lizzieLet60_1Lcall_f_f_Int3_d[51:36],
                                  (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[2]))};
  assign t1aes_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[67:52],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[3]))};
  assign is_zae6_2_destruct_d = (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[4]));
  assign op_addae7_2_destruct_d = (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[5]));
  assign q2ae9_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[83:68],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[6]))};
  assign \q2'aeo_1_destruct_d  = {lizzieLet60_1Lcall_f_f_Int3_d[99:84],
                                  (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[7]))};
  assign t2aet_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[115:100],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[8]))};
  assign q3aea_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[131:116],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[9]))};
  assign \q3'aep_1_destruct_d  = {lizzieLet60_1Lcall_f_f_Int3_d[147:132],
                                  (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[10]))};
  assign t3aeu_1_destruct_d = {lizzieLet60_1Lcall_f_f_Int3_d[163:148],
                               (lizzieLet60_1Lcall_f_f_Int3_d[0] && (! lizzieLet60_1Lcall_f_f_Int3_emitted[11]))};
  assign lizzieLet60_1Lcall_f_f_Int3_done = (lizzieLet60_1Lcall_f_f_Int3_emitted | ({t3aeu_1_destruct_d[0],
                                                                                     \q3'aep_1_destruct_d [0],
                                                                                     q3aea_1_destruct_d[0],
                                                                                     t2aet_1_destruct_d[0],
                                                                                     \q2'aeo_1_destruct_d [0],
                                                                                     q2ae9_1_destruct_d[0],
                                                                                     op_addae7_2_destruct_d[0],
                                                                                     is_zae6_2_destruct_d[0],
                                                                                     t1aes_1_destruct_d[0],
                                                                                     \q1'aen_1_destruct_d [0],
                                                                                     q1ae8_1_destruct_d[0],
                                                                                     sc_0_16_destruct_d[0]} & {t3aeu_1_destruct_r,
                                                                                                               \q3'aep_1_destruct_r ,
                                                                                                               q3aea_1_destruct_r,
                                                                                                               t2aet_1_destruct_r,
                                                                                                               \q2'aeo_1_destruct_r ,
                                                                                                               q2ae9_1_destruct_r,
                                                                                                               op_addae7_2_destruct_r,
                                                                                                               is_zae6_2_destruct_r,
                                                                                                               t1aes_1_destruct_r,
                                                                                                               \q1'aen_1_destruct_r ,
                                                                                                               q1ae8_1_destruct_r,
                                                                                                               sc_0_16_destruct_r}));
  assign lizzieLet60_1Lcall_f_f_Int3_r = (& lizzieLet60_1Lcall_f_f_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_1Lcall_f_f_Int3_emitted <= 12'd0;
    else
      lizzieLet60_1Lcall_f_f_Int3_emitted <= (lizzieLet60_1Lcall_f_f_Int3_r ? 12'd0 :
                                              lizzieLet60_1Lcall_f_f_Int3_done);
  
  /* demux (Ty CTf_f_Int,
       Ty CTf_f_Int) : (lizzieLet60_2,CTf_f_Int) (lizzieLet60_1,CTf_f_Int) > [(_22,CTf_f_Int),
                                                                              (lizzieLet60_1Lcall_f_f_Int3,CTf_f_Int),
                                                                              (lizzieLet60_1Lcall_f_f_Int2,CTf_f_Int),
                                                                              (lizzieLet60_1Lcall_f_f_Int1,CTf_f_Int),
                                                                              (lizzieLet60_1Lcall_f_f_Int0,CTf_f_Int)] */
  logic [4:0] lizzieLet60_1_onehotd;
  always_comb
    if ((lizzieLet60_2_d[0] && lizzieLet60_1_d[0]))
      unique case (lizzieLet60_2_d[3:1])
        3'd0: lizzieLet60_1_onehotd = 5'd1;
        3'd1: lizzieLet60_1_onehotd = 5'd2;
        3'd2: lizzieLet60_1_onehotd = 5'd4;
        3'd3: lizzieLet60_1_onehotd = 5'd8;
        3'd4: lizzieLet60_1_onehotd = 5'd16;
        default: lizzieLet60_1_onehotd = 5'd0;
      endcase
    else lizzieLet60_1_onehotd = 5'd0;
  assign _22_d = {lizzieLet60_1_d[163:1], lizzieLet60_1_onehotd[0]};
  assign lizzieLet60_1Lcall_f_f_Int3_d = {lizzieLet60_1_d[163:1],
                                          lizzieLet60_1_onehotd[1]};
  assign lizzieLet60_1Lcall_f_f_Int2_d = {lizzieLet60_1_d[163:1],
                                          lizzieLet60_1_onehotd[2]};
  assign lizzieLet60_1Lcall_f_f_Int1_d = {lizzieLet60_1_d[163:1],
                                          lizzieLet60_1_onehotd[3]};
  assign lizzieLet60_1Lcall_f_f_Int0_d = {lizzieLet60_1_d[163:1],
                                          lizzieLet60_1_onehotd[4]};
  assign lizzieLet60_1_r = (| (lizzieLet60_1_onehotd & {lizzieLet60_1Lcall_f_f_Int0_r,
                                                        lizzieLet60_1Lcall_f_f_Int1_r,
                                                        lizzieLet60_1Lcall_f_f_Int2_r,
                                                        lizzieLet60_1Lcall_f_f_Int3_r,
                                                        _22_r}));
  assign lizzieLet60_2_r = lizzieLet60_1_r;
  
  /* demux (Ty CTf_f_Int,
       Ty Go) : (lizzieLet60_3,CTf_f_Int) (go_18_goMux_data,Go) > [(_21,Go),
                                                                   (lizzieLet60_3Lcall_f_f_Int3,Go),
                                                                   (lizzieLet60_3Lcall_f_f_Int2,Go),
                                                                   (lizzieLet60_3Lcall_f_f_Int1,Go),
                                                                   (lizzieLet60_3Lcall_f_f_Int0,Go)] */
  logic [4:0] go_18_goMux_data_onehotd;
  always_comb
    if ((lizzieLet60_3_d[0] && go_18_goMux_data_d[0]))
      unique case (lizzieLet60_3_d[3:1])
        3'd0: go_18_goMux_data_onehotd = 5'd1;
        3'd1: go_18_goMux_data_onehotd = 5'd2;
        3'd2: go_18_goMux_data_onehotd = 5'd4;
        3'd3: go_18_goMux_data_onehotd = 5'd8;
        3'd4: go_18_goMux_data_onehotd = 5'd16;
        default: go_18_goMux_data_onehotd = 5'd0;
      endcase
    else go_18_goMux_data_onehotd = 5'd0;
  assign _21_d = go_18_goMux_data_onehotd[0];
  assign lizzieLet60_3Lcall_f_f_Int3_d = go_18_goMux_data_onehotd[1];
  assign lizzieLet60_3Lcall_f_f_Int2_d = go_18_goMux_data_onehotd[2];
  assign lizzieLet60_3Lcall_f_f_Int1_d = go_18_goMux_data_onehotd[3];
  assign lizzieLet60_3Lcall_f_f_Int0_d = go_18_goMux_data_onehotd[4];
  assign go_18_goMux_data_r = (| (go_18_goMux_data_onehotd & {lizzieLet60_3Lcall_f_f_Int0_r,
                                                              lizzieLet60_3Lcall_f_f_Int1_r,
                                                              lizzieLet60_3Lcall_f_f_Int2_r,
                                                              lizzieLet60_3Lcall_f_f_Int3_r,
                                                              _21_r}));
  assign lizzieLet60_3_r = go_18_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f_f_Int0,Go) > (lizzieLet60_3Lcall_f_f_Int0_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f_f_Int0_bufchan_d;
  logic lizzieLet60_3Lcall_f_f_Int0_bufchan_r;
  assign lizzieLet60_3Lcall_f_f_Int0_r = ((! lizzieLet60_3Lcall_f_f_Int0_bufchan_d[0]) || lizzieLet60_3Lcall_f_f_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f_f_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f_f_Int0_r)
        lizzieLet60_3Lcall_f_f_Int0_bufchan_d <= lizzieLet60_3Lcall_f_f_Int0_d;
  Go_t lizzieLet60_3Lcall_f_f_Int0_bufchan_buf;
  assign lizzieLet60_3Lcall_f_f_Int0_bufchan_r = (! lizzieLet60_3Lcall_f_f_Int0_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f_f_Int0_1_argbuf_d = (lizzieLet60_3Lcall_f_f_Int0_bufchan_buf[0] ? lizzieLet60_3Lcall_f_f_Int0_bufchan_buf :
                                                   lizzieLet60_3Lcall_f_f_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_3Lcall_f_f_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f_f_Int0_1_argbuf_r && lizzieLet60_3Lcall_f_f_Int0_bufchan_buf[0]))
        lizzieLet60_3Lcall_f_f_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f_f_Int0_1_argbuf_r) && (! lizzieLet60_3Lcall_f_f_Int0_bufchan_buf[0])))
        lizzieLet60_3Lcall_f_f_Int0_bufchan_buf <= lizzieLet60_3Lcall_f_f_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f_f_Int1,Go) > (lizzieLet60_3Lcall_f_f_Int1_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f_f_Int1_bufchan_d;
  logic lizzieLet60_3Lcall_f_f_Int1_bufchan_r;
  assign lizzieLet60_3Lcall_f_f_Int1_r = ((! lizzieLet60_3Lcall_f_f_Int1_bufchan_d[0]) || lizzieLet60_3Lcall_f_f_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f_f_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f_f_Int1_r)
        lizzieLet60_3Lcall_f_f_Int1_bufchan_d <= lizzieLet60_3Lcall_f_f_Int1_d;
  Go_t lizzieLet60_3Lcall_f_f_Int1_bufchan_buf;
  assign lizzieLet60_3Lcall_f_f_Int1_bufchan_r = (! lizzieLet60_3Lcall_f_f_Int1_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f_f_Int1_1_argbuf_d = (lizzieLet60_3Lcall_f_f_Int1_bufchan_buf[0] ? lizzieLet60_3Lcall_f_f_Int1_bufchan_buf :
                                                   lizzieLet60_3Lcall_f_f_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_3Lcall_f_f_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f_f_Int1_1_argbuf_r && lizzieLet60_3Lcall_f_f_Int1_bufchan_buf[0]))
        lizzieLet60_3Lcall_f_f_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f_f_Int1_1_argbuf_r) && (! lizzieLet60_3Lcall_f_f_Int1_bufchan_buf[0])))
        lizzieLet60_3Lcall_f_f_Int1_bufchan_buf <= lizzieLet60_3Lcall_f_f_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f_f_Int2,Go) > (lizzieLet60_3Lcall_f_f_Int2_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f_f_Int2_bufchan_d;
  logic lizzieLet60_3Lcall_f_f_Int2_bufchan_r;
  assign lizzieLet60_3Lcall_f_f_Int2_r = ((! lizzieLet60_3Lcall_f_f_Int2_bufchan_d[0]) || lizzieLet60_3Lcall_f_f_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f_f_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f_f_Int2_r)
        lizzieLet60_3Lcall_f_f_Int2_bufchan_d <= lizzieLet60_3Lcall_f_f_Int2_d;
  Go_t lizzieLet60_3Lcall_f_f_Int2_bufchan_buf;
  assign lizzieLet60_3Lcall_f_f_Int2_bufchan_r = (! lizzieLet60_3Lcall_f_f_Int2_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f_f_Int2_1_argbuf_d = (lizzieLet60_3Lcall_f_f_Int2_bufchan_buf[0] ? lizzieLet60_3Lcall_f_f_Int2_bufchan_buf :
                                                   lizzieLet60_3Lcall_f_f_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_3Lcall_f_f_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f_f_Int2_1_argbuf_r && lizzieLet60_3Lcall_f_f_Int2_bufchan_buf[0]))
        lizzieLet60_3Lcall_f_f_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f_f_Int2_1_argbuf_r) && (! lizzieLet60_3Lcall_f_f_Int2_bufchan_buf[0])))
        lizzieLet60_3Lcall_f_f_Int2_bufchan_buf <= lizzieLet60_3Lcall_f_f_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet60_3Lcall_f_f_Int3,Go) > (lizzieLet60_3Lcall_f_f_Int3_1_argbuf,Go) */
  Go_t lizzieLet60_3Lcall_f_f_Int3_bufchan_d;
  logic lizzieLet60_3Lcall_f_f_Int3_bufchan_r;
  assign lizzieLet60_3Lcall_f_f_Int3_r = ((! lizzieLet60_3Lcall_f_f_Int3_bufchan_d[0]) || lizzieLet60_3Lcall_f_f_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_3Lcall_f_f_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet60_3Lcall_f_f_Int3_r)
        lizzieLet60_3Lcall_f_f_Int3_bufchan_d <= lizzieLet60_3Lcall_f_f_Int3_d;
  Go_t lizzieLet60_3Lcall_f_f_Int3_bufchan_buf;
  assign lizzieLet60_3Lcall_f_f_Int3_bufchan_r = (! lizzieLet60_3Lcall_f_f_Int3_bufchan_buf[0]);
  assign lizzieLet60_3Lcall_f_f_Int3_1_argbuf_d = (lizzieLet60_3Lcall_f_f_Int3_bufchan_buf[0] ? lizzieLet60_3Lcall_f_f_Int3_bufchan_buf :
                                                   lizzieLet60_3Lcall_f_f_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_3Lcall_f_f_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet60_3Lcall_f_f_Int3_1_argbuf_r && lizzieLet60_3Lcall_f_f_Int3_bufchan_buf[0]))
        lizzieLet60_3Lcall_f_f_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet60_3Lcall_f_f_Int3_1_argbuf_r) && (! lizzieLet60_3Lcall_f_f_Int3_bufchan_buf[0])))
        lizzieLet60_3Lcall_f_f_Int3_bufchan_buf <= lizzieLet60_3Lcall_f_f_Int3_bufchan_d;
  
  /* demux (Ty CTf_f_Int,
       Ty Pointer_QTree_Int) : (lizzieLet60_4,CTf_f_Int) (srtarg_0_3_goMux_mux,Pointer_QTree_Int) > [(lizzieLet60_4Lf_f_Intsbos,Pointer_QTree_Int),
                                                                                                     (lizzieLet60_4Lcall_f_f_Int3,Pointer_QTree_Int),
                                                                                                     (lizzieLet60_4Lcall_f_f_Int2,Pointer_QTree_Int),
                                                                                                     (lizzieLet60_4Lcall_f_f_Int1,Pointer_QTree_Int),
                                                                                                     (lizzieLet60_4Lcall_f_f_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_3_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet60_4_d[0] && srtarg_0_3_goMux_mux_d[0]))
      unique case (lizzieLet60_4_d[3:1])
        3'd0: srtarg_0_3_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_3_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_3_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_3_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_3_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_3_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_3_goMux_mux_onehotd = 5'd0;
  assign lizzieLet60_4Lf_f_Intsbos_d = {srtarg_0_3_goMux_mux_d[16:1],
                                        srtarg_0_3_goMux_mux_onehotd[0]};
  assign lizzieLet60_4Lcall_f_f_Int3_d = {srtarg_0_3_goMux_mux_d[16:1],
                                          srtarg_0_3_goMux_mux_onehotd[1]};
  assign lizzieLet60_4Lcall_f_f_Int2_d = {srtarg_0_3_goMux_mux_d[16:1],
                                          srtarg_0_3_goMux_mux_onehotd[2]};
  assign lizzieLet60_4Lcall_f_f_Int1_d = {srtarg_0_3_goMux_mux_d[16:1],
                                          srtarg_0_3_goMux_mux_onehotd[3]};
  assign lizzieLet60_4Lcall_f_f_Int0_d = {srtarg_0_3_goMux_mux_d[16:1],
                                          srtarg_0_3_goMux_mux_onehotd[4]};
  assign srtarg_0_3_goMux_mux_r = (| (srtarg_0_3_goMux_mux_onehotd & {lizzieLet60_4Lcall_f_f_Int0_r,
                                                                      lizzieLet60_4Lcall_f_f_Int1_r,
                                                                      lizzieLet60_4Lcall_f_f_Int2_r,
                                                                      lizzieLet60_4Lcall_f_f_Int3_r,
                                                                      lizzieLet60_4Lf_f_Intsbos_r}));
  assign lizzieLet60_4_r = srtarg_0_3_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet60_4Lcall_f_f_Int0,Pointer_QTree_Int),
                         (es_12_destruct,Pointer_QTree_Int),
                         (es_13_1_destruct,Pointer_QTree_Int),
                         (es_14_2_destruct,Pointer_QTree_Int)] > (lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int,QTree_Int) */
  assign lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d = QNode_Int_dc((& {lizzieLet60_4Lcall_f_f_Int0_d[0],
                                                                                              es_12_destruct_d[0],
                                                                                              es_13_1_destruct_d[0],
                                                                                              es_14_2_destruct_d[0]}), lizzieLet60_4Lcall_f_f_Int0_d, es_12_destruct_d, es_13_1_destruct_d, es_14_2_destruct_d);
  assign {lizzieLet60_4Lcall_f_f_Int0_r,
          es_12_destruct_r,
          es_13_1_destruct_r,
          es_14_2_destruct_r} = {4 {(lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r && lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int,QTree_Int) > (lizzieLet64_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d;
  logic lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r;
  assign lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r = ((! lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d[0]) || lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d <= {66'd0,
                                                                                    1'd0};
    else
      if (lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r)
        lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d <= lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d;
  QTree_Int_t lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf;
  assign lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r = (! lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet64_1_argbuf_d = (lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf[0] ? lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf :
                                   lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                      1'd0};
    else
      if ((lizzieLet64_1_argbuf_r && lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf[0]))
        lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                        1'd0};
      else if (((! lizzieLet64_1_argbuf_r) && (! lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf[0])))
        lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf <= lizzieLet60_4Lcall_f_f_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int0) : [(lizzieLet60_4Lcall_f_f_Int1,Pointer_QTree_Int),
                              (es_13_destruct,Pointer_QTree_Int),
                              (es_14_1_destruct,Pointer_QTree_Int),
                              (sc_0_18_destruct,Pointer_CTf_f_Int)] > (lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0,CTf_f_Int) */
  assign lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_d = Lcall_f_f_Int0_dc((& {lizzieLet60_4Lcall_f_f_Int1_d[0],
                                                                                                        es_13_destruct_d[0],
                                                                                                        es_14_1_destruct_d[0],
                                                                                                        sc_0_18_destruct_d[0]}), lizzieLet60_4Lcall_f_f_Int1_d, es_13_destruct_d, es_14_1_destruct_d, sc_0_18_destruct_d);
  assign {lizzieLet60_4Lcall_f_f_Int1_r,
          es_13_destruct_r,
          es_14_1_destruct_r,
          sc_0_18_destruct_r} = {4 {(lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_r && lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_d[0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0,CTf_f_Int) > (lizzieLet63_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d;
  logic lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_r;
  assign lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_r = ((! lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d[0]) || lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d <= {163'd0,
                                                                                         1'd0};
    else
      if (lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_r)
        lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d <= lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_d;
  CTf_f_Int_t lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf;
  assign lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_r = (! lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf[0]);
  assign lizzieLet63_1_argbuf_d = (lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf[0] ? lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf :
                                   lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf <= {163'd0,
                                                                                           1'd0};
    else
      if ((lizzieLet63_1_argbuf_r && lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf[0]))
        lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf <= {163'd0,
                                                                                             1'd0};
      else if (((! lizzieLet63_1_argbuf_r) && (! lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf[0])))
        lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_buf <= lizzieLet60_4Lcall_f_f_Int1_1es_13_1es_14_1_1sc_0_18_1Lcall_f_f_Int0_bufchan_d;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int1) : [(lizzieLet60_4Lcall_f_f_Int2,Pointer_QTree_Int),
                              (es_14_destruct,Pointer_QTree_Int),
                              (sc_0_17_destruct,Pointer_CTf_f_Int),
                              (q1ae8_2_destruct,Pointer_MaskQTree),
                              (q1'aen_2_destruct,Pointer_QTree_Int),
                              (t1aes_2_destruct,Pointer_QTree_Int),
                              (is_zae6_3_1,MyDTInt_Bool),
                              (op_addae7_3_1,MyDTInt_Int_Int)] > (lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1,CTf_f_Int) */
  assign \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_d  = Lcall_f_f_Int1_dc((& {lizzieLet60_4Lcall_f_f_Int2_d[0],
                                                                                                                                                     es_14_destruct_d[0],
                                                                                                                                                     sc_0_17_destruct_d[0],
                                                                                                                                                     q1ae8_2_destruct_d[0],
                                                                                                                                                     \q1'aen_2_destruct_d [0],
                                                                                                                                                     t1aes_2_destruct_d[0],
                                                                                                                                                     is_zae6_3_1_d[0],
                                                                                                                                                     op_addae7_3_1_d[0]}), lizzieLet60_4Lcall_f_f_Int2_d, es_14_destruct_d, sc_0_17_destruct_d, q1ae8_2_destruct_d, \q1'aen_2_destruct_d , t1aes_2_destruct_d, is_zae6_3_1_d, op_addae7_3_1_d);
  assign {lizzieLet60_4Lcall_f_f_Int2_r,
          es_14_destruct_r,
          sc_0_17_destruct_r,
          q1ae8_2_destruct_r,
          \q1'aen_2_destruct_r ,
          t1aes_2_destruct_r,
          is_zae6_3_1_r,
          op_addae7_3_1_r} = {8 {(\lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_r  && \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_d [0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1,CTf_f_Int) > (lizzieLet62_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d ;
  logic \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_r ;
  assign \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_r  = ((! \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d [0]) || \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d  <= {163'd0,
                                                                                                                                      1'd0};
    else
      if (\lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_r )
        \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d  <= \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_d ;
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf ;
  assign \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_r  = (! \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf [0]);
  assign lizzieLet62_1_argbuf_d = (\lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf [0] ? \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf  :
                                   \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf  <= {163'd0,
                                                                                                                                        1'd0};
    else
      if ((lizzieLet62_1_argbuf_r && \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf [0]))
        \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf  <= {163'd0,
                                                                                                                                          1'd0};
      else if (((! lizzieLet62_1_argbuf_r) && (! \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf [0])))
        \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_buf  <= \lizzieLet60_4Lcall_f_f_Int2_1es_14_1sc_0_17_1q1ae8_2_1q1'aen_2_1t1aes_2_1is_zae6_3_1op_addae7_3_1Lcall_f_f_Int1_bufchan_d ;
  
  /* dcon (Ty CTf_f_Int,
      Dcon Lcall_f_f_Int2) : [(lizzieLet60_4Lcall_f_f_Int3,Pointer_QTree_Int),
                              (sc_0_16_destruct,Pointer_CTf_f_Int),
                              (q1ae8_1_destruct,Pointer_MaskQTree),
                              (q1'aen_1_destruct,Pointer_QTree_Int),
                              (t1aes_1_destruct,Pointer_QTree_Int),
                              (is_zae6_2_1,MyDTInt_Bool),
                              (op_addae7_2_1,MyDTInt_Int_Int),
                              (q2ae9_1_destruct,Pointer_MaskQTree),
                              (q2'aeo_1_destruct,Pointer_QTree_Int),
                              (t2aet_1_destruct,Pointer_QTree_Int)] > (lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2,CTf_f_Int) */
  assign \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_d  = Lcall_f_f_Int2_dc((& {lizzieLet60_4Lcall_f_f_Int3_d[0],
                                                                                                                                                                          sc_0_16_destruct_d[0],
                                                                                                                                                                          q1ae8_1_destruct_d[0],
                                                                                                                                                                          \q1'aen_1_destruct_d [0],
                                                                                                                                                                          t1aes_1_destruct_d[0],
                                                                                                                                                                          is_zae6_2_1_d[0],
                                                                                                                                                                          op_addae7_2_1_d[0],
                                                                                                                                                                          q2ae9_1_destruct_d[0],
                                                                                                                                                                          \q2'aeo_1_destruct_d [0],
                                                                                                                                                                          t2aet_1_destruct_d[0]}), lizzieLet60_4Lcall_f_f_Int3_d, sc_0_16_destruct_d, q1ae8_1_destruct_d, \q1'aen_1_destruct_d , t1aes_1_destruct_d, is_zae6_2_1_d, op_addae7_2_1_d, q2ae9_1_destruct_d, \q2'aeo_1_destruct_d , t2aet_1_destruct_d);
  assign {lizzieLet60_4Lcall_f_f_Int3_r,
          sc_0_16_destruct_r,
          q1ae8_1_destruct_r,
          \q1'aen_1_destruct_r ,
          t1aes_1_destruct_r,
          is_zae6_2_1_r,
          op_addae7_2_1_r,
          q2ae9_1_destruct_r,
          \q2'aeo_1_destruct_r ,
          t2aet_1_destruct_r} = {10 {(\lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_r  && \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_d [0])}};
  
  /* buf (Ty CTf_f_Int) : (lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2,CTf_f_Int) > (lizzieLet61_1_argbuf,CTf_f_Int) */
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d ;
  logic \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_r ;
  assign \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_r  = ((! \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d [0]) || \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d  <= {163'd0,
                                                                                                                                                           1'd0};
    else
      if (\lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_r )
        \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d  <= \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_d ;
  CTf_f_Int_t \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf ;
  assign \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_r  = (! \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf [0]);
  assign lizzieLet61_1_argbuf_d = (\lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf [0] ? \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf  :
                                   \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf  <= {163'd0,
                                                                                                                                                             1'd0};
    else
      if ((lizzieLet61_1_argbuf_r && \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf [0]))
        \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf  <= {163'd0,
                                                                                                                                                               1'd0};
      else if (((! lizzieLet61_1_argbuf_r) && (! \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf [0])))
        \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_buf  <= \lizzieLet60_4Lcall_f_f_Int3_1sc_0_16_1q1ae8_1_1q1'aen_1_1t1aes_1_1is_zae6_2_1op_addae7_2_1q2ae9_1_1q2'aeo_1_1t2aet_1_1Lcall_f_f_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet60_4Lf_f_Intsbos,Pointer_QTree_Int) > [(lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                               (lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet60_4Lf_f_Intsbos_emitted;
  logic [1:0] lizzieLet60_4Lf_f_Intsbos_done;
  assign lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_d = {lizzieLet60_4Lf_f_Intsbos_d[16:1],
                                                             (lizzieLet60_4Lf_f_Intsbos_d[0] && (! lizzieLet60_4Lf_f_Intsbos_emitted[0]))};
  assign lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_d = {lizzieLet60_4Lf_f_Intsbos_d[16:1],
                                                             (lizzieLet60_4Lf_f_Intsbos_d[0] && (! lizzieLet60_4Lf_f_Intsbos_emitted[1]))};
  assign lizzieLet60_4Lf_f_Intsbos_done = (lizzieLet60_4Lf_f_Intsbos_emitted | ({lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                 lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                         lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet60_4Lf_f_Intsbos_r = (& lizzieLet60_4Lf_f_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet60_4Lf_f_Intsbos_emitted <= 2'd0;
    else
      lizzieLet60_4Lf_f_Intsbos_emitted <= (lizzieLet60_4Lf_f_Intsbos_r ? 2'd0 :
                                            lizzieLet60_4Lf_f_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f_f_Int_goConst,Go) */
  assign call_f_f_Int_goConst_d = lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_1_r = call_f_f_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (f_f_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign f_f_Int_resbuf_d = (lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                             lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((f_f_Int_resbuf_r && lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! f_f_Int_resbuf_r) && (! lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet60_4Lf_f_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet6_1MQNode,MaskQTree) > [(q1aey_destruct,Pointer_MaskQTree),
                                                           (q2aez_destruct,Pointer_MaskQTree),
                                                           (q3aeA_destruct,Pointer_MaskQTree),
                                                           (q5aeB_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet6_1MQNode_emitted;
  logic [3:0] lizzieLet6_1MQNode_done;
  assign q1aey_destruct_d = {lizzieLet6_1MQNode_d[18:3],
                             (lizzieLet6_1MQNode_d[0] && (! lizzieLet6_1MQNode_emitted[0]))};
  assign q2aez_destruct_d = {lizzieLet6_1MQNode_d[34:19],
                             (lizzieLet6_1MQNode_d[0] && (! lizzieLet6_1MQNode_emitted[1]))};
  assign q3aeA_destruct_d = {lizzieLet6_1MQNode_d[50:35],
                             (lizzieLet6_1MQNode_d[0] && (! lizzieLet6_1MQNode_emitted[2]))};
  assign q5aeB_destruct_d = {lizzieLet6_1MQNode_d[66:51],
                             (lizzieLet6_1MQNode_d[0] && (! lizzieLet6_1MQNode_emitted[3]))};
  assign lizzieLet6_1MQNode_done = (lizzieLet6_1MQNode_emitted | ({q5aeB_destruct_d[0],
                                                                   q3aeA_destruct_d[0],
                                                                   q2aez_destruct_d[0],
                                                                   q1aey_destruct_d[0]} & {q5aeB_destruct_r,
                                                                                           q3aeA_destruct_r,
                                                                                           q2aez_destruct_r,
                                                                                           q1aey_destruct_r}));
  assign lizzieLet6_1MQNode_r = (& lizzieLet6_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1MQNode_emitted <= 4'd0;
    else
      lizzieLet6_1MQNode_emitted <= (lizzieLet6_1MQNode_r ? 4'd0 :
                                     lizzieLet6_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet6_2,MaskQTree) (lizzieLet6_1,MaskQTree) > [(_20,MaskQTree),
                                                                            (_19,MaskQTree),
                                                                            (lizzieLet6_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 3'd1;
        2'd1: lizzieLet6_1_onehotd = 3'd2;
        2'd2: lizzieLet6_1_onehotd = 3'd4;
        default: lizzieLet6_1_onehotd = 3'd0;
      endcase
    else lizzieLet6_1_onehotd = 3'd0;
  assign _20_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign _19_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1MQNode_d = {lizzieLet6_1_d[66:1],
                                 lizzieLet6_1_onehotd[2]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {lizzieLet6_1MQNode_r,
                                                      _19_r,
                                                      _20_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet6_3,MaskQTree) (go_9_goMux_data,Go) > [(lizzieLet6_3MQNone,Go),
                                                                 (lizzieLet6_3MQVal,Go),
                                                                 (lizzieLet6_3MQNode,Go)] */
  logic [2:0] go_9_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && go_9_goMux_data_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: go_9_goMux_data_onehotd = 3'd1;
        2'd1: go_9_goMux_data_onehotd = 3'd2;
        2'd2: go_9_goMux_data_onehotd = 3'd4;
        default: go_9_goMux_data_onehotd = 3'd0;
      endcase
    else go_9_goMux_data_onehotd = 3'd0;
  assign lizzieLet6_3MQNone_d = go_9_goMux_data_onehotd[0];
  assign lizzieLet6_3MQVal_d = go_9_goMux_data_onehotd[1];
  assign lizzieLet6_3MQNode_d = go_9_goMux_data_onehotd[2];
  assign go_9_goMux_data_r = (| (go_9_goMux_data_onehotd & {lizzieLet6_3MQNode_r,
                                                            lizzieLet6_3MQVal_r,
                                                            lizzieLet6_3MQNone_r}));
  assign lizzieLet6_3_r = go_9_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_3MQNone,Go) > [(lizzieLet6_3MQNone_1,Go),
                                          (lizzieLet6_3MQNone_2,Go)] */
  logic [1:0] lizzieLet6_3MQNone_emitted;
  logic [1:0] lizzieLet6_3MQNone_done;
  assign lizzieLet6_3MQNone_1_d = (lizzieLet6_3MQNone_d[0] && (! lizzieLet6_3MQNone_emitted[0]));
  assign lizzieLet6_3MQNone_2_d = (lizzieLet6_3MQNone_d[0] && (! lizzieLet6_3MQNone_emitted[1]));
  assign lizzieLet6_3MQNone_done = (lizzieLet6_3MQNone_emitted | ({lizzieLet6_3MQNone_2_d[0],
                                                                   lizzieLet6_3MQNone_1_d[0]} & {lizzieLet6_3MQNone_2_r,
                                                                                                 lizzieLet6_3MQNone_1_r}));
  assign lizzieLet6_3MQNone_r = (& lizzieLet6_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQNone_emitted <= 2'd0;
    else
      lizzieLet6_3MQNone_emitted <= (lizzieLet6_3MQNone_r ? 2'd0 :
                                     lizzieLet6_3MQNone_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_3MQNone_1,Go)] > (lizzieLet6_3MQNone_1QNone_Int,QTree_Int) */
  assign lizzieLet6_3MQNone_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_3MQNone_1_d[0]}), lizzieLet6_3MQNone_1_d);
  assign {lizzieLet6_3MQNone_1_r} = {1 {(lizzieLet6_3MQNone_1QNone_Int_r && lizzieLet6_3MQNone_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_3MQNone_1QNone_Int,QTree_Int) > (lizzieLet7_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_3MQNone_1QNone_Int_bufchan_d;
  logic lizzieLet6_3MQNone_1QNone_Int_bufchan_r;
  assign lizzieLet6_3MQNone_1QNone_Int_r = ((! lizzieLet6_3MQNone_1QNone_Int_bufchan_d[0]) || lizzieLet6_3MQNone_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3MQNone_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_3MQNone_1QNone_Int_r)
        lizzieLet6_3MQNone_1QNone_Int_bufchan_d <= lizzieLet6_3MQNone_1QNone_Int_d;
  QTree_Int_t lizzieLet6_3MQNone_1QNone_Int_bufchan_buf;
  assign lizzieLet6_3MQNone_1QNone_Int_bufchan_r = (! lizzieLet6_3MQNone_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_3MQNone_1QNone_Int_bufchan_buf[0] ? lizzieLet6_3MQNone_1QNone_Int_bufchan_buf :
                                  lizzieLet6_3MQNone_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_3MQNone_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_3MQNone_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_3MQNone_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_3MQNone_1QNone_Int_bufchan_buf <= lizzieLet6_3MQNone_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_3MQNone_2,Go) > (lizzieLet6_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet6_3MQNone_2_bufchan_d;
  logic lizzieLet6_3MQNone_2_bufchan_r;
  assign lizzieLet6_3MQNone_2_r = ((! lizzieLet6_3MQNone_2_bufchan_d[0]) || lizzieLet6_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3MQNone_2_r)
        lizzieLet6_3MQNone_2_bufchan_d <= lizzieLet6_3MQNone_2_d;
  Go_t lizzieLet6_3MQNone_2_bufchan_buf;
  assign lizzieLet6_3MQNone_2_bufchan_r = (! lizzieLet6_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet6_3MQNone_2_argbuf_d = (lizzieLet6_3MQNone_2_bufchan_buf[0] ? lizzieLet6_3MQNone_2_bufchan_buf :
                                          lizzieLet6_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3MQNone_2_argbuf_r && lizzieLet6_3MQNone_2_bufchan_buf[0]))
        lizzieLet6_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3MQNone_2_argbuf_r) && (! lizzieLet6_3MQNone_2_bufchan_buf[0])))
        lizzieLet6_3MQNone_2_bufchan_buf <= lizzieLet6_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet6_3MQNone_2_argbuf,Go),
                           (lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf,Go),
                           (lizzieLet6_3MQVal_1_argbuf,Go),
                           (lizzieLet6_4MQNode_3QNone_Int_2_argbuf,Go),
                           (lizzieLet6_4MQNode_3QVal_Int_2_argbuf,Go),
                           (lizzieLet6_4MQNode_3QError_Int_2_argbuf,Go)] > (go_16_goMux_choice,C6) (go_16_goMux_data,Go) */
  logic [5:0] lizzieLet6_3MQNone_2_argbuf_select_d;
  assign lizzieLet6_3MQNone_2_argbuf_select_d = ((| lizzieLet6_3MQNone_2_argbuf_select_q) ? lizzieLet6_3MQNone_2_argbuf_select_q :
                                                 (lizzieLet6_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                  (\lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_d [0] ? 6'd2 :
                                                   (lizzieLet6_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                    (lizzieLet6_4MQNode_3QNone_Int_2_argbuf_d[0] ? 6'd8 :
                                                     (lizzieLet6_4MQNode_3QVal_Int_2_argbuf_d[0] ? 6'd16 :
                                                      (lizzieLet6_4MQNode_3QError_Int_2_argbuf_d[0] ? 6'd32 :
                                                       6'd0)))))));
  logic [5:0] lizzieLet6_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet6_3MQNone_2_argbuf_select_q <= (lizzieLet6_3MQNone_2_argbuf_done ? 6'd0 :
                                               lizzieLet6_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet6_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_3MQNone_2_argbuf_emit_q <= (lizzieLet6_3MQNone_2_argbuf_done ? 2'd0 :
                                             lizzieLet6_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_3MQNone_2_argbuf_emit_d;
  assign lizzieLet6_3MQNone_2_argbuf_emit_d = (lizzieLet6_3MQNone_2_argbuf_emit_q | ({go_16_goMux_choice_d[0],
                                                                                      go_16_goMux_data_d[0]} & {go_16_goMux_choice_r,
                                                                                                                go_16_goMux_data_r}));
  logic lizzieLet6_3MQNone_2_argbuf_done;
  assign lizzieLet6_3MQNone_2_argbuf_done = (& lizzieLet6_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet6_4MQNode_3QError_Int_2_argbuf_r,
          lizzieLet6_4MQNode_3QVal_Int_2_argbuf_r,
          lizzieLet6_4MQNode_3QNone_Int_2_argbuf_r,
          lizzieLet6_3MQVal_1_argbuf_r,
          \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_r ,
          lizzieLet6_3MQNone_2_argbuf_r} = (lizzieLet6_3MQNone_2_argbuf_done ? lizzieLet6_3MQNone_2_argbuf_select_d :
                                            6'd0);
  assign go_16_goMux_data_d = ((lizzieLet6_3MQNone_2_argbuf_select_d[0] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet6_3MQNone_2_argbuf_d :
                               ((lizzieLet6_3MQNone_2_argbuf_select_d[1] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? \lizzieLet50_3Lcall_f'''''''''_f'''''''''_Int0_1_argbuf_d  :
                                ((lizzieLet6_3MQNone_2_argbuf_select_d[2] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet6_3MQVal_1_argbuf_d :
                                 ((lizzieLet6_3MQNone_2_argbuf_select_d[3] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet6_4MQNode_3QNone_Int_2_argbuf_d :
                                  ((lizzieLet6_3MQNone_2_argbuf_select_d[4] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet6_4MQNode_3QVal_Int_2_argbuf_d :
                                   ((lizzieLet6_3MQNone_2_argbuf_select_d[5] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet6_4MQNode_3QError_Int_2_argbuf_d :
                                    1'd0))))));
  assign go_16_goMux_choice_d = ((lizzieLet6_3MQNone_2_argbuf_select_d[0] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet6_3MQNone_2_argbuf_select_d[1] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet6_3MQNone_2_argbuf_select_d[2] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet6_3MQNone_2_argbuf_select_d[3] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet6_3MQNone_2_argbuf_select_d[4] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet6_3MQNone_2_argbuf_select_d[5] && (! lizzieLet6_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet6_3MQVal,Go) > (lizzieLet6_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet6_3MQVal_bufchan_d;
  logic lizzieLet6_3MQVal_bufchan_r;
  assign lizzieLet6_3MQVal_r = ((! lizzieLet6_3MQVal_bufchan_d[0]) || lizzieLet6_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3MQVal_r)
        lizzieLet6_3MQVal_bufchan_d <= lizzieLet6_3MQVal_d;
  Go_t lizzieLet6_3MQVal_bufchan_buf;
  assign lizzieLet6_3MQVal_bufchan_r = (! lizzieLet6_3MQVal_bufchan_buf[0]);
  assign lizzieLet6_3MQVal_1_argbuf_d = (lizzieLet6_3MQVal_bufchan_buf[0] ? lizzieLet6_3MQVal_bufchan_buf :
                                         lizzieLet6_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3MQVal_1_argbuf_r && lizzieLet6_3MQVal_bufchan_buf[0]))
        lizzieLet6_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3MQVal_1_argbuf_r) && (! lizzieLet6_3MQVal_bufchan_buf[0])))
        lizzieLet6_3MQVal_bufchan_buf <= lizzieLet6_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Int) : (lizzieLet6_4,MaskQTree) (readPointer_QTree_Intq4'aex_1_argbuf_rwb,QTree_Int) > [(_18,QTree_Int),
                                                                                                        (_17,QTree_Int),
                                                                                                        (lizzieLet6_4MQNode,QTree_Int)] */
  logic [2:0] \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd ;
  always_comb
    if ((lizzieLet6_4_d[0] && \readPointer_QTree_Intq4'aex_1_argbuf_rwb_d [0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  = 3'd1;
        2'd1: \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  = 3'd2;
        2'd2: \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  = 3'd4;
        default: \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  = 3'd0;
      endcase
    else \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  = 3'd0;
  assign _18_d = {\readPointer_QTree_Intq4'aex_1_argbuf_rwb_d [66:1],
                  \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd [0]};
  assign _17_d = {\readPointer_QTree_Intq4'aex_1_argbuf_rwb_d [66:1],
                  \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd [1]};
  assign lizzieLet6_4MQNode_d = {\readPointer_QTree_Intq4'aex_1_argbuf_rwb_d [66:1],
                                 \readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd [2]};
  assign \readPointer_QTree_Intq4'aex_1_argbuf_rwb_r  = (| (\readPointer_QTree_Intq4'aex_1_argbuf_rwb_onehotd  & {lizzieLet6_4MQNode_r,
                                                                                                                  _17_r,
                                                                                                                  _18_r}));
  assign lizzieLet6_4_r = \readPointer_QTree_Intq4'aex_1_argbuf_rwb_r ;
  
  /* fork (Ty QTree_Int) : (lizzieLet6_4MQNode,QTree_Int) > [(lizzieLet6_4MQNode_1,QTree_Int),
                                                        (lizzieLet6_4MQNode_2,QTree_Int),
                                                        (lizzieLet6_4MQNode_3,QTree_Int),
                                                        (lizzieLet6_4MQNode_4,QTree_Int),
                                                        (lizzieLet6_4MQNode_5,QTree_Int),
                                                        (lizzieLet6_4MQNode_6,QTree_Int),
                                                        (lizzieLet6_4MQNode_7,QTree_Int),
                                                        (lizzieLet6_4MQNode_8,QTree_Int)] */
  logic [7:0] lizzieLet6_4MQNode_emitted;
  logic [7:0] lizzieLet6_4MQNode_done;
  assign lizzieLet6_4MQNode_1_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[0]))};
  assign lizzieLet6_4MQNode_2_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[1]))};
  assign lizzieLet6_4MQNode_3_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[2]))};
  assign lizzieLet6_4MQNode_4_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[3]))};
  assign lizzieLet6_4MQNode_5_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[4]))};
  assign lizzieLet6_4MQNode_6_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[5]))};
  assign lizzieLet6_4MQNode_7_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[6]))};
  assign lizzieLet6_4MQNode_8_d = {lizzieLet6_4MQNode_d[66:1],
                                   (lizzieLet6_4MQNode_d[0] && (! lizzieLet6_4MQNode_emitted[7]))};
  assign lizzieLet6_4MQNode_done = (lizzieLet6_4MQNode_emitted | ({lizzieLet6_4MQNode_8_d[0],
                                                                   lizzieLet6_4MQNode_7_d[0],
                                                                   lizzieLet6_4MQNode_6_d[0],
                                                                   lizzieLet6_4MQNode_5_d[0],
                                                                   lizzieLet6_4MQNode_4_d[0],
                                                                   lizzieLet6_4MQNode_3_d[0],
                                                                   lizzieLet6_4MQNode_2_d[0],
                                                                   lizzieLet6_4MQNode_1_d[0]} & {lizzieLet6_4MQNode_8_r,
                                                                                                 lizzieLet6_4MQNode_7_r,
                                                                                                 lizzieLet6_4MQNode_6_r,
                                                                                                 lizzieLet6_4MQNode_5_r,
                                                                                                 lizzieLet6_4MQNode_4_r,
                                                                                                 lizzieLet6_4MQNode_3_r,
                                                                                                 lizzieLet6_4MQNode_2_r,
                                                                                                 lizzieLet6_4MQNode_1_r}));
  assign lizzieLet6_4MQNode_r = (& lizzieLet6_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4MQNode_emitted <= 8'd0;
    else
      lizzieLet6_4MQNode_emitted <= (lizzieLet6_4MQNode_r ? 8'd0 :
                                     lizzieLet6_4MQNode_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_4MQNode_1QNode_Int,QTree_Int) > [(t1aeD_destruct,Pointer_QTree_Int),
                                                                         (t2aeE_destruct,Pointer_QTree_Int),
                                                                         (t3aeF_destruct,Pointer_QTree_Int),
                                                                         (t4aeG_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_4MQNode_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_4MQNode_1QNode_Int_done;
  assign t1aeD_destruct_d = {lizzieLet6_4MQNode_1QNode_Int_d[18:3],
                             (lizzieLet6_4MQNode_1QNode_Int_d[0] && (! lizzieLet6_4MQNode_1QNode_Int_emitted[0]))};
  assign t2aeE_destruct_d = {lizzieLet6_4MQNode_1QNode_Int_d[34:19],
                             (lizzieLet6_4MQNode_1QNode_Int_d[0] && (! lizzieLet6_4MQNode_1QNode_Int_emitted[1]))};
  assign t3aeF_destruct_d = {lizzieLet6_4MQNode_1QNode_Int_d[50:35],
                             (lizzieLet6_4MQNode_1QNode_Int_d[0] && (! lizzieLet6_4MQNode_1QNode_Int_emitted[2]))};
  assign t4aeG_destruct_d = {lizzieLet6_4MQNode_1QNode_Int_d[66:51],
                             (lizzieLet6_4MQNode_1QNode_Int_d[0] && (! lizzieLet6_4MQNode_1QNode_Int_emitted[3]))};
  assign lizzieLet6_4MQNode_1QNode_Int_done = (lizzieLet6_4MQNode_1QNode_Int_emitted | ({t4aeG_destruct_d[0],
                                                                                         t3aeF_destruct_d[0],
                                                                                         t2aeE_destruct_d[0],
                                                                                         t1aeD_destruct_d[0]} & {t4aeG_destruct_r,
                                                                                                                 t3aeF_destruct_r,
                                                                                                                 t2aeE_destruct_r,
                                                                                                                 t1aeD_destruct_r}));
  assign lizzieLet6_4MQNode_1QNode_Int_r = (& lizzieLet6_4MQNode_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4MQNode_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_4MQNode_1QNode_Int_emitted <= (lizzieLet6_4MQNode_1QNode_Int_r ? 4'd0 :
                                                lizzieLet6_4MQNode_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_4MQNode_2,QTree_Int) (lizzieLet6_4MQNode_1,QTree_Int) > [(_16,QTree_Int),
                                                                                            (_15,QTree_Int),
                                                                                            (lizzieLet6_4MQNode_1QNode_Int,QTree_Int),
                                                                                            (_14,QTree_Int)] */
  logic [3:0] lizzieLet6_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_2_d[0] && lizzieLet6_4MQNode_1_d[0]))
      unique case (lizzieLet6_4MQNode_2_d[2:1])
        2'd0: lizzieLet6_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet6_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet6_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet6_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet6_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_4MQNode_1_onehotd = 4'd0;
  assign _16_d = {lizzieLet6_4MQNode_1_d[66:1],
                  lizzieLet6_4MQNode_1_onehotd[0]};
  assign _15_d = {lizzieLet6_4MQNode_1_d[66:1],
                  lizzieLet6_4MQNode_1_onehotd[1]};
  assign lizzieLet6_4MQNode_1QNode_Int_d = {lizzieLet6_4MQNode_1_d[66:1],
                                            lizzieLet6_4MQNode_1_onehotd[2]};
  assign _14_d = {lizzieLet6_4MQNode_1_d[66:1],
                  lizzieLet6_4MQNode_1_onehotd[3]};
  assign lizzieLet6_4MQNode_1_r = (| (lizzieLet6_4MQNode_1_onehotd & {_14_r,
                                                                      lizzieLet6_4MQNode_1QNode_Int_r,
                                                                      _15_r,
                                                                      _16_r}));
  assign lizzieLet6_4MQNode_2_r = lizzieLet6_4MQNode_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_4MQNode_3,QTree_Int) (lizzieLet6_3MQNode,Go) > [(lizzieLet6_4MQNode_3QNone_Int,Go),
                                                                            (lizzieLet6_4MQNode_3QVal_Int,Go),
                                                                            (lizzieLet6_4MQNode_3QNode_Int,Go),
                                                                            (lizzieLet6_4MQNode_3QError_Int,Go)] */
  logic [3:0] lizzieLet6_3MQNode_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_3_d[0] && lizzieLet6_3MQNode_d[0]))
      unique case (lizzieLet6_4MQNode_3_d[2:1])
        2'd0: lizzieLet6_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet6_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet6_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet6_3MQNode_onehotd = 4'd8;
        default: lizzieLet6_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet6_3MQNode_onehotd = 4'd0;
  assign lizzieLet6_4MQNode_3QNone_Int_d = lizzieLet6_3MQNode_onehotd[0];
  assign lizzieLet6_4MQNode_3QVal_Int_d = lizzieLet6_3MQNode_onehotd[1];
  assign lizzieLet6_4MQNode_3QNode_Int_d = lizzieLet6_3MQNode_onehotd[2];
  assign lizzieLet6_4MQNode_3QError_Int_d = lizzieLet6_3MQNode_onehotd[3];
  assign lizzieLet6_3MQNode_r = (| (lizzieLet6_3MQNode_onehotd & {lizzieLet6_4MQNode_3QError_Int_r,
                                                                  lizzieLet6_4MQNode_3QNode_Int_r,
                                                                  lizzieLet6_4MQNode_3QVal_Int_r,
                                                                  lizzieLet6_4MQNode_3QNone_Int_r}));
  assign lizzieLet6_4MQNode_3_r = lizzieLet6_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet6_4MQNode_3QError_Int,Go) > [(lizzieLet6_4MQNode_3QError_Int_1,Go),
                                                      (lizzieLet6_4MQNode_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_4MQNode_3QError_Int_emitted;
  logic [1:0] lizzieLet6_4MQNode_3QError_Int_done;
  assign lizzieLet6_4MQNode_3QError_Int_1_d = (lizzieLet6_4MQNode_3QError_Int_d[0] && (! lizzieLet6_4MQNode_3QError_Int_emitted[0]));
  assign lizzieLet6_4MQNode_3QError_Int_2_d = (lizzieLet6_4MQNode_3QError_Int_d[0] && (! lizzieLet6_4MQNode_3QError_Int_emitted[1]));
  assign lizzieLet6_4MQNode_3QError_Int_done = (lizzieLet6_4MQNode_3QError_Int_emitted | ({lizzieLet6_4MQNode_3QError_Int_2_d[0],
                                                                                           lizzieLet6_4MQNode_3QError_Int_1_d[0]} & {lizzieLet6_4MQNode_3QError_Int_2_r,
                                                                                                                                     lizzieLet6_4MQNode_3QError_Int_1_r}));
  assign lizzieLet6_4MQNode_3QError_Int_r = (& lizzieLet6_4MQNode_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_4MQNode_3QError_Int_emitted <= (lizzieLet6_4MQNode_3QError_Int_r ? 2'd0 :
                                                 lizzieLet6_4MQNode_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_4MQNode_3QError_Int_1,Go)] > (lizzieLet6_4MQNode_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_4MQNode_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_4MQNode_3QError_Int_1_d[0]}), lizzieLet6_4MQNode_3QError_Int_1_d);
  assign {lizzieLet6_4MQNode_3QError_Int_1_r} = {1 {(lizzieLet6_4MQNode_3QError_Int_1QError_Int_r && lizzieLet6_4MQNode_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4MQNode_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet12_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_4MQNode_3QError_Int_1QError_Int_r = ((! lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                               1'd0};
    else
      if (lizzieLet6_4MQNode_3QError_Int_1QError_Int_r)
        lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d <= lizzieLet6_4MQNode_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_4MQNode_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4MQNode_3QError_Int_2,Go) > (lizzieLet6_4MQNode_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4MQNode_3QError_Int_2_bufchan_d;
  logic lizzieLet6_4MQNode_3QError_Int_2_bufchan_r;
  assign lizzieLet6_4MQNode_3QError_Int_2_r = ((! lizzieLet6_4MQNode_3QError_Int_2_bufchan_d[0]) || lizzieLet6_4MQNode_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4MQNode_3QError_Int_2_r)
        lizzieLet6_4MQNode_3QError_Int_2_bufchan_d <= lizzieLet6_4MQNode_3QError_Int_2_d;
  Go_t lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf;
  assign lizzieLet6_4MQNode_3QError_Int_2_bufchan_r = (! lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_3QError_Int_2_argbuf_d = (lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf[0] ? lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf :
                                                      lizzieLet6_4MQNode_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4MQNode_3QError_Int_2_argbuf_r && lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4MQNode_3QError_Int_2_argbuf_r) && (! lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QError_Int_2_bufchan_buf <= lizzieLet6_4MQNode_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4MQNode_3QNode_Int,Go) > (lizzieLet6_4MQNode_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4MQNode_3QNode_Int_bufchan_d;
  logic lizzieLet6_4MQNode_3QNode_Int_bufchan_r;
  assign lizzieLet6_4MQNode_3QNode_Int_r = ((! lizzieLet6_4MQNode_3QNode_Int_bufchan_d[0]) || lizzieLet6_4MQNode_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4MQNode_3QNode_Int_r)
        lizzieLet6_4MQNode_3QNode_Int_bufchan_d <= lizzieLet6_4MQNode_3QNode_Int_d;
  Go_t lizzieLet6_4MQNode_3QNode_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_3QNode_Int_bufchan_r = (! lizzieLet6_4MQNode_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_3QNode_Int_1_argbuf_d = (lizzieLet6_4MQNode_3QNode_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_3QNode_Int_bufchan_buf :
                                                     lizzieLet6_4MQNode_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4MQNode_3QNode_Int_1_argbuf_r && lizzieLet6_4MQNode_3QNode_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4MQNode_3QNode_Int_1_argbuf_r) && (! lizzieLet6_4MQNode_3QNode_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QNode_Int_bufchan_buf <= lizzieLet6_4MQNode_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4MQNode_3QNone_Int,Go) > [(lizzieLet6_4MQNode_3QNone_Int_1,Go),
                                                     (lizzieLet6_4MQNode_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet6_4MQNode_3QNone_Int_emitted;
  logic [1:0] lizzieLet6_4MQNode_3QNone_Int_done;
  assign lizzieLet6_4MQNode_3QNone_Int_1_d = (lizzieLet6_4MQNode_3QNone_Int_d[0] && (! lizzieLet6_4MQNode_3QNone_Int_emitted[0]));
  assign lizzieLet6_4MQNode_3QNone_Int_2_d = (lizzieLet6_4MQNode_3QNone_Int_d[0] && (! lizzieLet6_4MQNode_3QNone_Int_emitted[1]));
  assign lizzieLet6_4MQNode_3QNone_Int_done = (lizzieLet6_4MQNode_3QNone_Int_emitted | ({lizzieLet6_4MQNode_3QNone_Int_2_d[0],
                                                                                         lizzieLet6_4MQNode_3QNone_Int_1_d[0]} & {lizzieLet6_4MQNode_3QNone_Int_2_r,
                                                                                                                                  lizzieLet6_4MQNode_3QNone_Int_1_r}));
  assign lizzieLet6_4MQNode_3QNone_Int_r = (& lizzieLet6_4MQNode_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4MQNode_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet6_4MQNode_3QNone_Int_emitted <= (lizzieLet6_4MQNode_3QNone_Int_r ? 2'd0 :
                                                lizzieLet6_4MQNode_3QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_4MQNode_3QNone_Int_1,Go)] > (lizzieLet6_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_4MQNode_3QNone_Int_1_d[0]}), lizzieLet6_4MQNode_3QNone_Int_1_d);
  assign {lizzieLet6_4MQNode_3QNone_Int_1_r} = {1 {(lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_r && lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4MQNode_3QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_r = ((! lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= {66'd0,
                                                             1'd0};
    else
      if (lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_r)
        lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d <= lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf :
                                  lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                               1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= {66'd0,
                                                                 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet6_4MQNode_3QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4MQNode_3QNone_Int_2,Go) > (lizzieLet6_4MQNode_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d;
  logic lizzieLet6_4MQNode_3QNone_Int_2_bufchan_r;
  assign lizzieLet6_4MQNode_3QNone_Int_2_r = ((! lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d[0]) || lizzieLet6_4MQNode_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4MQNode_3QNone_Int_2_r)
        lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d <= lizzieLet6_4MQNode_3QNone_Int_2_d;
  Go_t lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf;
  assign lizzieLet6_4MQNode_3QNone_Int_2_bufchan_r = (! lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_3QNone_Int_2_argbuf_d = (lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf[0] ? lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf :
                                                     lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4MQNode_3QNone_Int_2_argbuf_r && lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4MQNode_3QNone_Int_2_argbuf_r) && (! lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QNone_Int_2_bufchan_buf <= lizzieLet6_4MQNode_3QNone_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4MQNode_3QVal_Int,Go) > [(lizzieLet6_4MQNode_3QVal_Int_1,Go),
                                                    (lizzieLet6_4MQNode_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_4MQNode_3QVal_Int_emitted;
  logic [1:0] lizzieLet6_4MQNode_3QVal_Int_done;
  assign lizzieLet6_4MQNode_3QVal_Int_1_d = (lizzieLet6_4MQNode_3QVal_Int_d[0] && (! lizzieLet6_4MQNode_3QVal_Int_emitted[0]));
  assign lizzieLet6_4MQNode_3QVal_Int_2_d = (lizzieLet6_4MQNode_3QVal_Int_d[0] && (! lizzieLet6_4MQNode_3QVal_Int_emitted[1]));
  assign lizzieLet6_4MQNode_3QVal_Int_done = (lizzieLet6_4MQNode_3QVal_Int_emitted | ({lizzieLet6_4MQNode_3QVal_Int_2_d[0],
                                                                                       lizzieLet6_4MQNode_3QVal_Int_1_d[0]} & {lizzieLet6_4MQNode_3QVal_Int_2_r,
                                                                                                                               lizzieLet6_4MQNode_3QVal_Int_1_r}));
  assign lizzieLet6_4MQNode_3QVal_Int_r = (& lizzieLet6_4MQNode_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4MQNode_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_4MQNode_3QVal_Int_emitted <= (lizzieLet6_4MQNode_3QVal_Int_r ? 2'd0 :
                                               lizzieLet6_4MQNode_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_4MQNode_3QVal_Int_1,Go)] > (lizzieLet6_4MQNode_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_4MQNode_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_4MQNode_3QVal_Int_1_d[0]}), lizzieLet6_4MQNode_3QVal_Int_1_d);
  assign {lizzieLet6_4MQNode_3QVal_Int_1_r} = {1 {(lizzieLet6_4MQNode_3QVal_Int_1QError_Int_r && lizzieLet6_4MQNode_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4MQNode_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet10_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_4MQNode_3QVal_Int_1QError_Int_r = ((! lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                             1'd0};
    else
      if (lizzieLet6_4MQNode_3QVal_Int_1QError_Int_r)
        lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet6_4MQNode_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf :
                                   lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                               1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet6_4MQNode_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4MQNode_3QVal_Int_2,Go) > (lizzieLet6_4MQNode_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d;
  logic lizzieLet6_4MQNode_3QVal_Int_2_bufchan_r;
  assign lizzieLet6_4MQNode_3QVal_Int_2_r = ((! lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d[0]) || lizzieLet6_4MQNode_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4MQNode_3QVal_Int_2_r)
        lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d <= lizzieLet6_4MQNode_3QVal_Int_2_d;
  Go_t lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf;
  assign lizzieLet6_4MQNode_3QVal_Int_2_bufchan_r = (! lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_3QVal_Int_2_argbuf_d = (lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf[0] ? lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf :
                                                    lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4MQNode_3QVal_Int_2_argbuf_r && lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4MQNode_3QVal_Int_2_argbuf_r) && (! lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet6_4MQNode_3QVal_Int_2_bufchan_buf <= lizzieLet6_4MQNode_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_4MQNode_4,QTree_Int) (lizzieLet6_6MQNode,Pointer_CTf'''''''''_f'''''''''_Int) > [(lizzieLet6_4MQNode_4QNone_Int,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                              (lizzieLet6_4MQNode_4QVal_Int,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                              (lizzieLet6_4MQNode_4QNode_Int,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                              (lizzieLet6_4MQNode_4QError_Int,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [3:0] lizzieLet6_6MQNode_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_4_d[0] && lizzieLet6_6MQNode_d[0]))
      unique case (lizzieLet6_4MQNode_4_d[2:1])
        2'd0: lizzieLet6_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet6_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet6_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet6_6MQNode_onehotd = 4'd8;
        default: lizzieLet6_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet6_6MQNode_onehotd = 4'd0;
  assign lizzieLet6_4MQNode_4QNone_Int_d = {lizzieLet6_6MQNode_d[16:1],
                                            lizzieLet6_6MQNode_onehotd[0]};
  assign lizzieLet6_4MQNode_4QVal_Int_d = {lizzieLet6_6MQNode_d[16:1],
                                           lizzieLet6_6MQNode_onehotd[1]};
  assign lizzieLet6_4MQNode_4QNode_Int_d = {lizzieLet6_6MQNode_d[16:1],
                                            lizzieLet6_6MQNode_onehotd[2]};
  assign lizzieLet6_4MQNode_4QError_Int_d = {lizzieLet6_6MQNode_d[16:1],
                                             lizzieLet6_6MQNode_onehotd[3]};
  assign lizzieLet6_6MQNode_r = (| (lizzieLet6_6MQNode_onehotd & {lizzieLet6_4MQNode_4QError_Int_r,
                                                                  lizzieLet6_4MQNode_4QNode_Int_r,
                                                                  lizzieLet6_4MQNode_4QVal_Int_r,
                                                                  lizzieLet6_4MQNode_4QNone_Int_r}));
  assign lizzieLet6_4MQNode_4_r = lizzieLet6_6MQNode_r;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_4MQNode_4QError_Int,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet6_4MQNode_4QError_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QError_Int_bufchan_d;
  logic lizzieLet6_4MQNode_4QError_Int_bufchan_r;
  assign lizzieLet6_4MQNode_4QError_Int_r = ((! lizzieLet6_4MQNode_4QError_Int_bufchan_d[0]) || lizzieLet6_4MQNode_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_4MQNode_4QError_Int_r)
        lizzieLet6_4MQNode_4QError_Int_bufchan_d <= lizzieLet6_4MQNode_4QError_Int_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QError_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_4QError_Int_bufchan_r = (! lizzieLet6_4MQNode_4QError_Int_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_4QError_Int_1_argbuf_d = (lizzieLet6_4MQNode_4QError_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_4QError_Int_bufchan_buf :
                                                      lizzieLet6_4MQNode_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_4MQNode_4QError_Int_1_argbuf_r && lizzieLet6_4MQNode_4QError_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_4MQNode_4QError_Int_1_argbuf_r) && (! lizzieLet6_4MQNode_4QError_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_4QError_Int_bufchan_buf <= lizzieLet6_4MQNode_4QError_Int_bufchan_d;
  
  /* dcon (Ty CTf'''''''''_f'''''''''_Int,
      Dcon Lcall_f'''''''''_f'''''''''_Int3) : [(lizzieLet6_4MQNode_4QNode_Int,Pointer_CTf'''''''''_f'''''''''_Int),
                                                (lizzieLet6_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                                (t1aeD_destruct,Pointer_QTree_Int),
                                                (lizzieLet6_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                                (t2aeE_destruct,Pointer_QTree_Int),
                                                (lizzieLet6_4MQNode_7QNode_Int,Pointer_MaskQTree),
                                                (t3aeF_destruct,Pointer_QTree_Int)] > (lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3,CTf'''''''''_f'''''''''_Int) */
  assign \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_d  = \Lcall_f'''''''''_f'''''''''_Int3_dc ((& {lizzieLet6_4MQNode_4QNode_Int_d[0],
                                                                                                                                                                                                                                           lizzieLet6_4MQNode_5QNode_Int_d[0],
                                                                                                                                                                                                                                           t1aeD_destruct_d[0],
                                                                                                                                                                                                                                           lizzieLet6_4MQNode_6QNode_Int_d[0],
                                                                                                                                                                                                                                           t2aeE_destruct_d[0],
                                                                                                                                                                                                                                           lizzieLet6_4MQNode_7QNode_Int_d[0],
                                                                                                                                                                                                                                           t3aeF_destruct_d[0]}), lizzieLet6_4MQNode_4QNode_Int_d, lizzieLet6_4MQNode_5QNode_Int_d, t1aeD_destruct_d, lizzieLet6_4MQNode_6QNode_Int_d, t2aeE_destruct_d, lizzieLet6_4MQNode_7QNode_Int_d, t3aeF_destruct_d);
  assign {lizzieLet6_4MQNode_4QNode_Int_r,
          lizzieLet6_4MQNode_5QNode_Int_r,
          t1aeD_destruct_r,
          lizzieLet6_4MQNode_6QNode_Int_r,
          t2aeE_destruct_r,
          lizzieLet6_4MQNode_7QNode_Int_r,
          t3aeF_destruct_r} = {7 {(\lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_r  && \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_d [0])}};
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3,CTf'''''''''_f'''''''''_Int) > (lizzieLet11_1_argbuf,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d ;
  logic \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_r ;
  assign \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_r  = ((! \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d [0]) || \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d  <= {115'd0,
                                                                                                                                                                                                        1'd0};
    else
      if (\lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_r )
        \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d  <= \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_d ;
  \CTf'''''''''_f'''''''''_Int_t  \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf ;
  assign \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_r  = (! \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0]);
  assign lizzieLet11_1_argbuf_d = (\lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0] ? \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  :
                                   \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                          1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0]))
        \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= {115'd0,
                                                                                                                                                                                                            1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf [0])))
        \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_buf  <= \lizzieLet6_4MQNode_4QNode_Int_1lizzieLet6_4MQNode_5QNode_Int_1t1aeD_1lizzieLet6_4MQNode_6QNode_Int_1t2aeE_1lizzieLet6_4MQNode_7QNode_Int_1t3aeF_1Lcall_f'''''''''_f'''''''''_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_4MQNode_4QNone_Int,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet6_4MQNode_4QNone_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QNone_Int_bufchan_d;
  logic lizzieLet6_4MQNode_4QNone_Int_bufchan_r;
  assign lizzieLet6_4MQNode_4QNone_Int_r = ((! lizzieLet6_4MQNode_4QNone_Int_bufchan_d[0]) || lizzieLet6_4MQNode_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_4MQNode_4QNone_Int_r)
        lizzieLet6_4MQNode_4QNone_Int_bufchan_d <= lizzieLet6_4MQNode_4QNone_Int_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QNone_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_4QNone_Int_bufchan_r = (! lizzieLet6_4MQNode_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_4QNone_Int_1_argbuf_d = (lizzieLet6_4MQNode_4QNone_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_4QNone_Int_bufchan_buf :
                                                     lizzieLet6_4MQNode_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_4MQNode_4QNone_Int_1_argbuf_r && lizzieLet6_4MQNode_4QNone_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_4MQNode_4QNone_Int_1_argbuf_r) && (! lizzieLet6_4MQNode_4QNone_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_4QNone_Int_bufchan_buf <= lizzieLet6_4MQNode_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_4MQNode_4QVal_Int,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet6_4MQNode_4QVal_Int_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QVal_Int_bufchan_d;
  logic lizzieLet6_4MQNode_4QVal_Int_bufchan_r;
  assign lizzieLet6_4MQNode_4QVal_Int_r = ((! lizzieLet6_4MQNode_4QVal_Int_bufchan_d[0]) || lizzieLet6_4MQNode_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_4MQNode_4QVal_Int_r)
        lizzieLet6_4MQNode_4QVal_Int_bufchan_d <= lizzieLet6_4MQNode_4QVal_Int_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_4MQNode_4QVal_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_4QVal_Int_bufchan_r = (! lizzieLet6_4MQNode_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_4QVal_Int_1_argbuf_d = (lizzieLet6_4MQNode_4QVal_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_4QVal_Int_bufchan_buf :
                                                    lizzieLet6_4MQNode_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_4MQNode_4QVal_Int_1_argbuf_r && lizzieLet6_4MQNode_4QVal_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_4MQNode_4QVal_Int_1_argbuf_r) && (! lizzieLet6_4MQNode_4QVal_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_4QVal_Int_bufchan_buf <= lizzieLet6_4MQNode_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet6_4MQNode_5,QTree_Int) (q1aey_destruct,Pointer_MaskQTree) > [(_13,Pointer_MaskQTree),
                                                                                                      (_12,Pointer_MaskQTree),
                                                                                                      (lizzieLet6_4MQNode_5QNode_Int,Pointer_MaskQTree),
                                                                                                      (_11,Pointer_MaskQTree)] */
  logic [3:0] q1aey_destruct_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_5_d[0] && q1aey_destruct_d[0]))
      unique case (lizzieLet6_4MQNode_5_d[2:1])
        2'd0: q1aey_destruct_onehotd = 4'd1;
        2'd1: q1aey_destruct_onehotd = 4'd2;
        2'd2: q1aey_destruct_onehotd = 4'd4;
        2'd3: q1aey_destruct_onehotd = 4'd8;
        default: q1aey_destruct_onehotd = 4'd0;
      endcase
    else q1aey_destruct_onehotd = 4'd0;
  assign _13_d = {q1aey_destruct_d[16:1], q1aey_destruct_onehotd[0]};
  assign _12_d = {q1aey_destruct_d[16:1], q1aey_destruct_onehotd[1]};
  assign lizzieLet6_4MQNode_5QNode_Int_d = {q1aey_destruct_d[16:1],
                                            q1aey_destruct_onehotd[2]};
  assign _11_d = {q1aey_destruct_d[16:1], q1aey_destruct_onehotd[3]};
  assign q1aey_destruct_r = (| (q1aey_destruct_onehotd & {_11_r,
                                                          lizzieLet6_4MQNode_5QNode_Int_r,
                                                          _12_r,
                                                          _13_r}));
  assign lizzieLet6_4MQNode_5_r = q1aey_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet6_4MQNode_6,QTree_Int) (q2aez_destruct,Pointer_MaskQTree) > [(_10,Pointer_MaskQTree),
                                                                                                      (_9,Pointer_MaskQTree),
                                                                                                      (lizzieLet6_4MQNode_6QNode_Int,Pointer_MaskQTree),
                                                                                                      (_8,Pointer_MaskQTree)] */
  logic [3:0] q2aez_destruct_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_6_d[0] && q2aez_destruct_d[0]))
      unique case (lizzieLet6_4MQNode_6_d[2:1])
        2'd0: q2aez_destruct_onehotd = 4'd1;
        2'd1: q2aez_destruct_onehotd = 4'd2;
        2'd2: q2aez_destruct_onehotd = 4'd4;
        2'd3: q2aez_destruct_onehotd = 4'd8;
        default: q2aez_destruct_onehotd = 4'd0;
      endcase
    else q2aez_destruct_onehotd = 4'd0;
  assign _10_d = {q2aez_destruct_d[16:1], q2aez_destruct_onehotd[0]};
  assign _9_d = {q2aez_destruct_d[16:1], q2aez_destruct_onehotd[1]};
  assign lizzieLet6_4MQNode_6QNode_Int_d = {q2aez_destruct_d[16:1],
                                            q2aez_destruct_onehotd[2]};
  assign _8_d = {q2aez_destruct_d[16:1], q2aez_destruct_onehotd[3]};
  assign q2aez_destruct_r = (| (q2aez_destruct_onehotd & {_8_r,
                                                          lizzieLet6_4MQNode_6QNode_Int_r,
                                                          _9_r,
                                                          _10_r}));
  assign lizzieLet6_4MQNode_6_r = q2aez_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet6_4MQNode_7,QTree_Int) (q3aeA_destruct,Pointer_MaskQTree) > [(_7,Pointer_MaskQTree),
                                                                                                      (_6,Pointer_MaskQTree),
                                                                                                      (lizzieLet6_4MQNode_7QNode_Int,Pointer_MaskQTree),
                                                                                                      (_5,Pointer_MaskQTree)] */
  logic [3:0] q3aeA_destruct_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_7_d[0] && q3aeA_destruct_d[0]))
      unique case (lizzieLet6_4MQNode_7_d[2:1])
        2'd0: q3aeA_destruct_onehotd = 4'd1;
        2'd1: q3aeA_destruct_onehotd = 4'd2;
        2'd2: q3aeA_destruct_onehotd = 4'd4;
        2'd3: q3aeA_destruct_onehotd = 4'd8;
        default: q3aeA_destruct_onehotd = 4'd0;
      endcase
    else q3aeA_destruct_onehotd = 4'd0;
  assign _7_d = {q3aeA_destruct_d[16:1], q3aeA_destruct_onehotd[0]};
  assign _6_d = {q3aeA_destruct_d[16:1], q3aeA_destruct_onehotd[1]};
  assign lizzieLet6_4MQNode_7QNode_Int_d = {q3aeA_destruct_d[16:1],
                                            q3aeA_destruct_onehotd[2]};
  assign _5_d = {q3aeA_destruct_d[16:1], q3aeA_destruct_onehotd[3]};
  assign q3aeA_destruct_r = (| (q3aeA_destruct_onehotd & {_5_r,
                                                          lizzieLet6_4MQNode_7QNode_Int_r,
                                                          _6_r,
                                                          _7_r}));
  assign lizzieLet6_4MQNode_7_r = q3aeA_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_MaskQTree) : (lizzieLet6_4MQNode_8,QTree_Int) (q5aeB_destruct,Pointer_MaskQTree) > [(_4,Pointer_MaskQTree),
                                                                                                      (_3,Pointer_MaskQTree),
                                                                                                      (lizzieLet6_4MQNode_8QNode_Int,Pointer_MaskQTree),
                                                                                                      (_2,Pointer_MaskQTree)] */
  logic [3:0] q5aeB_destruct_onehotd;
  always_comb
    if ((lizzieLet6_4MQNode_8_d[0] && q5aeB_destruct_d[0]))
      unique case (lizzieLet6_4MQNode_8_d[2:1])
        2'd0: q5aeB_destruct_onehotd = 4'd1;
        2'd1: q5aeB_destruct_onehotd = 4'd2;
        2'd2: q5aeB_destruct_onehotd = 4'd4;
        2'd3: q5aeB_destruct_onehotd = 4'd8;
        default: q5aeB_destruct_onehotd = 4'd0;
      endcase
    else q5aeB_destruct_onehotd = 4'd0;
  assign _4_d = {q5aeB_destruct_d[16:1], q5aeB_destruct_onehotd[0]};
  assign _3_d = {q5aeB_destruct_d[16:1], q5aeB_destruct_onehotd[1]};
  assign lizzieLet6_4MQNode_8QNode_Int_d = {q5aeB_destruct_d[16:1],
                                            q5aeB_destruct_onehotd[2]};
  assign _2_d = {q5aeB_destruct_d[16:1], q5aeB_destruct_onehotd[3]};
  assign q5aeB_destruct_r = (| (q5aeB_destruct_onehotd & {_2_r,
                                                          lizzieLet6_4MQNode_8QNode_Int_r,
                                                          _3_r,
                                                          _4_r}));
  assign lizzieLet6_4MQNode_8_r = q5aeB_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet6_4MQNode_8QNode_Int,Pointer_MaskQTree) > (lizzieLet6_4MQNode_8QNode_Int_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet6_4MQNode_8QNode_Int_bufchan_d;
  logic lizzieLet6_4MQNode_8QNode_Int_bufchan_r;
  assign lizzieLet6_4MQNode_8QNode_Int_r = ((! lizzieLet6_4MQNode_8QNode_Int_bufchan_d[0]) || lizzieLet6_4MQNode_8QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_8QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_4MQNode_8QNode_Int_r)
        lizzieLet6_4MQNode_8QNode_Int_bufchan_d <= lizzieLet6_4MQNode_8QNode_Int_d;
  Pointer_MaskQTree_t lizzieLet6_4MQNode_8QNode_Int_bufchan_buf;
  assign lizzieLet6_4MQNode_8QNode_Int_bufchan_r = (! lizzieLet6_4MQNode_8QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_4MQNode_8QNode_Int_1_argbuf_d = (lizzieLet6_4MQNode_8QNode_Int_bufchan_buf[0] ? lizzieLet6_4MQNode_8QNode_Int_bufchan_buf :
                                                     lizzieLet6_4MQNode_8QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_4MQNode_8QNode_Int_1_argbuf_r && lizzieLet6_4MQNode_8QNode_Int_bufchan_buf[0]))
        lizzieLet6_4MQNode_8QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_4MQNode_8QNode_Int_1_argbuf_r) && (! lizzieLet6_4MQNode_8QNode_Int_bufchan_buf[0])))
        lizzieLet6_4MQNode_8QNode_Int_bufchan_buf <= lizzieLet6_4MQNode_8QNode_Int_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Int) : (lizzieLet6_5,MaskQTree) (q4'aex_2,Pointer_QTree_Int) > [(_1,Pointer_QTree_Int),
                                                                                        (lizzieLet6_5MQVal,Pointer_QTree_Int),
                                                                                        (_0,Pointer_QTree_Int)] */
  logic [2:0] \q4'aex_2_onehotd ;
  always_comb
    if ((lizzieLet6_5_d[0] && \q4'aex_2_d [0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: \q4'aex_2_onehotd  = 3'd1;
        2'd1: \q4'aex_2_onehotd  = 3'd2;
        2'd2: \q4'aex_2_onehotd  = 3'd4;
        default: \q4'aex_2_onehotd  = 3'd0;
      endcase
    else \q4'aex_2_onehotd  = 3'd0;
  assign _1_d = {\q4'aex_2_d [16:1], \q4'aex_2_onehotd [0]};
  assign lizzieLet6_5MQVal_d = {\q4'aex_2_d [16:1],
                                \q4'aex_2_onehotd [1]};
  assign _0_d = {\q4'aex_2_d [16:1], \q4'aex_2_onehotd [2]};
  assign \q4'aex_2_r  = (| (\q4'aex_2_onehotd  & {_0_r,
                                                  lizzieLet6_5MQVal_r,
                                                  _1_r}));
  assign lizzieLet6_5_r = \q4'aex_2_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet6_5MQVal,Pointer_QTree_Int) > (lizzieLet6_5MQVal_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet6_5MQVal_bufchan_d;
  logic lizzieLet6_5MQVal_bufchan_r;
  assign lizzieLet6_5MQVal_r = ((! lizzieLet6_5MQVal_bufchan_d[0]) || lizzieLet6_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_5MQVal_r)
        lizzieLet6_5MQVal_bufchan_d <= lizzieLet6_5MQVal_d;
  Pointer_QTree_Int_t lizzieLet6_5MQVal_bufchan_buf;
  assign lizzieLet6_5MQVal_bufchan_r = (! lizzieLet6_5MQVal_bufchan_buf[0]);
  assign lizzieLet6_5MQVal_1_argbuf_d = (lizzieLet6_5MQVal_bufchan_buf[0] ? lizzieLet6_5MQVal_bufchan_buf :
                                         lizzieLet6_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_5MQVal_1_argbuf_r && lizzieLet6_5MQVal_bufchan_buf[0]))
        lizzieLet6_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_5MQVal_1_argbuf_r) && (! lizzieLet6_5MQVal_bufchan_buf[0])))
        lizzieLet6_5MQVal_bufchan_buf <= lizzieLet6_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_6,MaskQTree) (sc_0_1_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Int) > [(lizzieLet6_6MQNone,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet6_6MQVal,Pointer_CTf'''''''''_f'''''''''_Int),
                                                                                                                                    (lizzieLet6_6MQNode,Pointer_CTf'''''''''_f'''''''''_Int)] */
  logic [2:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 3'd4;
        default: sc_0_1_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 3'd0;
  assign lizzieLet6_6MQNone_d = {sc_0_1_goMux_mux_d[16:1],
                                 sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_6MQVal_d = {sc_0_1_goMux_mux_d[16:1],
                                sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_6MQNode_d = {sc_0_1_goMux_mux_d[16:1],
                                 sc_0_1_goMux_mux_onehotd[2]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_6MQNode_r,
                                                              lizzieLet6_6MQVal_r,
                                                              lizzieLet6_6MQNone_r}));
  assign lizzieLet6_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_6MQNone,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet6_6MQNone_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQNone_bufchan_d;
  logic lizzieLet6_6MQNone_bufchan_r;
  assign lizzieLet6_6MQNone_r = ((! lizzieLet6_6MQNone_bufchan_d[0]) || lizzieLet6_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6MQNone_r)
        lizzieLet6_6MQNone_bufchan_d <= lizzieLet6_6MQNone_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQNone_bufchan_buf;
  assign lizzieLet6_6MQNone_bufchan_r = (! lizzieLet6_6MQNone_bufchan_buf[0]);
  assign lizzieLet6_6MQNone_1_argbuf_d = (lizzieLet6_6MQNone_bufchan_buf[0] ? lizzieLet6_6MQNone_bufchan_buf :
                                          lizzieLet6_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6MQNone_1_argbuf_r && lizzieLet6_6MQNone_bufchan_buf[0]))
        lizzieLet6_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6MQNone_1_argbuf_r) && (! lizzieLet6_6MQNone_bufchan_buf[0])))
        lizzieLet6_6MQNone_bufchan_buf <= lizzieLet6_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (lizzieLet6_6MQVal,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet6_6MQVal_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQVal_bufchan_d;
  logic lizzieLet6_6MQVal_bufchan_r;
  assign lizzieLet6_6MQVal_r = ((! lizzieLet6_6MQVal_bufchan_d[0]) || lizzieLet6_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6MQVal_r)
        lizzieLet6_6MQVal_bufchan_d <= lizzieLet6_6MQVal_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  lizzieLet6_6MQVal_bufchan_buf;
  assign lizzieLet6_6MQVal_bufchan_r = (! lizzieLet6_6MQVal_bufchan_buf[0]);
  assign lizzieLet6_6MQVal_1_argbuf_d = (lizzieLet6_6MQVal_bufchan_buf[0] ? lizzieLet6_6MQVal_bufchan_buf :
                                         lizzieLet6_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6MQVal_1_argbuf_r && lizzieLet6_6MQVal_bufchan_buf[0]))
        lizzieLet6_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6MQVal_1_argbuf_r) && (! lizzieLet6_6MQVal_bufchan_buf[0])))
        lizzieLet6_6MQVal_bufchan_buf <= lizzieLet6_6MQVal_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (m1ae3_goMux_mux,Pointer_MaskQTree) > (m1ae3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t m1ae3_goMux_mux_bufchan_d;
  logic m1ae3_goMux_mux_bufchan_r;
  assign m1ae3_goMux_mux_r = ((! m1ae3_goMux_mux_bufchan_d[0]) || m1ae3_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae3_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1ae3_goMux_mux_r)
        m1ae3_goMux_mux_bufchan_d <= m1ae3_goMux_mux_d;
  Pointer_MaskQTree_t m1ae3_goMux_mux_bufchan_buf;
  assign m1ae3_goMux_mux_bufchan_r = (! m1ae3_goMux_mux_bufchan_buf[0]);
  assign m1ae3_1_argbuf_d = (m1ae3_goMux_mux_bufchan_buf[0] ? m1ae3_goMux_mux_bufchan_buf :
                             m1ae3_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ae3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1ae3_1_argbuf_r && m1ae3_goMux_mux_bufchan_buf[0]))
        m1ae3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1ae3_1_argbuf_r) && (! m1ae3_goMux_mux_bufchan_buf[0])))
        m1ae3_goMux_mux_bufchan_buf <= m1ae3_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2ae4_1,Pointer_QTree_Int) > (m2ae4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ae4_1_bufchan_d;
  logic m2ae4_1_bufchan_r;
  assign m2ae4_1_r = ((! m2ae4_1_bufchan_d[0]) || m2ae4_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae4_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2ae4_1_r) m2ae4_1_bufchan_d <= m2ae4_1_d;
  Pointer_QTree_Int_t m2ae4_1_bufchan_buf;
  assign m2ae4_1_bufchan_r = (! m2ae4_1_bufchan_buf[0]);
  assign m2ae4_1_argbuf_d = (m2ae4_1_bufchan_buf[0] ? m2ae4_1_bufchan_buf :
                             m2ae4_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae4_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ae4_1_argbuf_r && m2ae4_1_bufchan_buf[0]))
        m2ae4_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ae4_1_argbuf_r) && (! m2ae4_1_bufchan_buf[0])))
        m2ae4_1_bufchan_buf <= m2ae4_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2ae4_goMux_mux,Pointer_QTree_Int) > [(m2ae4_1,Pointer_QTree_Int),
                                                                     (m2ae4_2,Pointer_QTree_Int)] */
  logic [1:0] m2ae4_goMux_mux_emitted;
  logic [1:0] m2ae4_goMux_mux_done;
  assign m2ae4_1_d = {m2ae4_goMux_mux_d[16:1],
                      (m2ae4_goMux_mux_d[0] && (! m2ae4_goMux_mux_emitted[0]))};
  assign m2ae4_2_d = {m2ae4_goMux_mux_d[16:1],
                      (m2ae4_goMux_mux_d[0] && (! m2ae4_goMux_mux_emitted[1]))};
  assign m2ae4_goMux_mux_done = (m2ae4_goMux_mux_emitted | ({m2ae4_2_d[0],
                                                             m2ae4_1_d[0]} & {m2ae4_2_r,
                                                                              m2ae4_1_r}));
  assign m2ae4_goMux_mux_r = (& m2ae4_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ae4_goMux_mux_emitted <= 2'd0;
    else
      m2ae4_goMux_mux_emitted <= (m2ae4_goMux_mux_r ? 2'd0 :
                                  m2ae4_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2aeH_1,Pointer_QTree_Int) > (m2aeH_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2aeH_1_bufchan_d;
  logic m2aeH_1_bufchan_r;
  assign m2aeH_1_r = ((! m2aeH_1_bufchan_d[0]) || m2aeH_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aeH_1_bufchan_d <= {16'd0, 1'd0};
    else if (m2aeH_1_r) m2aeH_1_bufchan_d <= m2aeH_1_d;
  Pointer_QTree_Int_t m2aeH_1_bufchan_buf;
  assign m2aeH_1_bufchan_r = (! m2aeH_1_bufchan_buf[0]);
  assign m2aeH_1_argbuf_d = (m2aeH_1_bufchan_buf[0] ? m2aeH_1_bufchan_buf :
                             m2aeH_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aeH_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2aeH_1_argbuf_r && m2aeH_1_bufchan_buf[0]))
        m2aeH_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2aeH_1_argbuf_r) && (! m2aeH_1_bufchan_buf[0])))
        m2aeH_1_bufchan_buf <= m2aeH_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2aeH_goMux_mux,Pointer_QTree_Int) > [(m2aeH_1,Pointer_QTree_Int),
                                                                     (m2aeH_2,Pointer_QTree_Int)] */
  logic [1:0] m2aeH_goMux_mux_emitted;
  logic [1:0] m2aeH_goMux_mux_done;
  assign m2aeH_1_d = {m2aeH_goMux_mux_d[16:1],
                      (m2aeH_goMux_mux_d[0] && (! m2aeH_goMux_mux_emitted[0]))};
  assign m2aeH_2_d = {m2aeH_goMux_mux_d[16:1],
                      (m2aeH_goMux_mux_d[0] && (! m2aeH_goMux_mux_emitted[1]))};
  assign m2aeH_goMux_mux_done = (m2aeH_goMux_mux_emitted | ({m2aeH_2_d[0],
                                                             m2aeH_1_d[0]} & {m2aeH_2_r,
                                                                              m2aeH_1_r}));
  assign m2aeH_goMux_mux_r = (& m2aeH_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2aeH_goMux_mux_emitted <= 2'd0;
    else
      m2aeH_goMux_mux_emitted <= (m2aeH_goMux_mux_r ? 2'd0 :
                                  m2aeH_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m3ae5_1,Pointer_QTree_Int) > (m3ae5_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m3ae5_1_bufchan_d;
  logic m3ae5_1_bufchan_r;
  assign m3ae5_1_r = ((! m3ae5_1_bufchan_d[0]) || m3ae5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3ae5_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3ae5_1_r) m3ae5_1_bufchan_d <= m3ae5_1_d;
  Pointer_QTree_Int_t m3ae5_1_bufchan_buf;
  assign m3ae5_1_bufchan_r = (! m3ae5_1_bufchan_buf[0]);
  assign m3ae5_1_argbuf_d = (m3ae5_1_bufchan_buf[0] ? m3ae5_1_bufchan_buf :
                             m3ae5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3ae5_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3ae5_1_argbuf_r && m3ae5_1_bufchan_buf[0]))
        m3ae5_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3ae5_1_argbuf_r) && (! m3ae5_1_bufchan_buf[0])))
        m3ae5_1_bufchan_buf <= m3ae5_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m3ae5_goMux_mux,Pointer_QTree_Int) > [(m3ae5_1,Pointer_QTree_Int),
                                                                     (m3ae5_2,Pointer_QTree_Int)] */
  logic [1:0] m3ae5_goMux_mux_emitted;
  logic [1:0] m3ae5_goMux_mux_done;
  assign m3ae5_1_d = {m3ae5_goMux_mux_d[16:1],
                      (m3ae5_goMux_mux_d[0] && (! m3ae5_goMux_mux_emitted[0]))};
  assign m3ae5_2_d = {m3ae5_goMux_mux_d[16:1],
                      (m3ae5_goMux_mux_d[0] && (! m3ae5_goMux_mux_emitted[1]))};
  assign m3ae5_goMux_mux_done = (m3ae5_goMux_mux_emitted | ({m3ae5_2_d[0],
                                                             m3ae5_1_d[0]} & {m3ae5_2_r,
                                                                              m3ae5_1_r}));
  assign m3ae5_goMux_mux_r = (& m3ae5_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3ae5_goMux_mux_emitted <= 2'd0;
    else
      m3ae5_goMux_mux_emitted <= (m3ae5_goMux_mux_r ? 2'd0 :
                                  m3ae5_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m3aeI_1,Pointer_QTree_Int) > (m3aeI_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m3aeI_1_bufchan_d;
  logic m3aeI_1_bufchan_r;
  assign m3aeI_1_r = ((! m3aeI_1_bufchan_d[0]) || m3aeI_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aeI_1_bufchan_d <= {16'd0, 1'd0};
    else if (m3aeI_1_r) m3aeI_1_bufchan_d <= m3aeI_1_d;
  Pointer_QTree_Int_t m3aeI_1_bufchan_buf;
  assign m3aeI_1_bufchan_r = (! m3aeI_1_bufchan_buf[0]);
  assign m3aeI_1_argbuf_d = (m3aeI_1_bufchan_buf[0] ? m3aeI_1_bufchan_buf :
                             m3aeI_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aeI_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m3aeI_1_argbuf_r && m3aeI_1_bufchan_buf[0]))
        m3aeI_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m3aeI_1_argbuf_r) && (! m3aeI_1_bufchan_buf[0])))
        m3aeI_1_bufchan_buf <= m3aeI_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m3aeI_goMux_mux,Pointer_QTree_Int) > [(m3aeI_1,Pointer_QTree_Int),
                                                                     (m3aeI_2,Pointer_QTree_Int)] */
  logic [1:0] m3aeI_goMux_mux_emitted;
  logic [1:0] m3aeI_goMux_mux_done;
  assign m3aeI_1_d = {m3aeI_goMux_mux_d[16:1],
                      (m3aeI_goMux_mux_d[0] && (! m3aeI_goMux_mux_emitted[0]))};
  assign m3aeI_2_d = {m3aeI_goMux_mux_d[16:1],
                      (m3aeI_goMux_mux_d[0] && (! m3aeI_goMux_mux_emitted[1]))};
  assign m3aeI_goMux_mux_done = (m3aeI_goMux_mux_emitted | ({m3aeI_2_d[0],
                                                             m3aeI_1_d[0]} & {m3aeI_2_r,
                                                                              m3aeI_1_r}));
  assign m3aeI_goMux_mux_r = (& m3aeI_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m3aeI_goMux_mux_emitted <= 2'd0;
    else
      m3aeI_goMux_mux_emitted <= (m3aeI_goMux_mux_r ? 2'd0 :
                                  m3aeI_goMux_mux_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addae7_2_2,MyDTInt_Int_Int) > (op_addae7_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addae7_2_2_bufchan_d;
  logic op_addae7_2_2_bufchan_r;
  assign op_addae7_2_2_r = ((! op_addae7_2_2_bufchan_d[0]) || op_addae7_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_2_2_bufchan_d <= 1'd0;
    else
      if (op_addae7_2_2_r) op_addae7_2_2_bufchan_d <= op_addae7_2_2_d;
  MyDTInt_Int_Int_t op_addae7_2_2_bufchan_buf;
  assign op_addae7_2_2_bufchan_r = (! op_addae7_2_2_bufchan_buf[0]);
  assign op_addae7_2_2_argbuf_d = (op_addae7_2_2_bufchan_buf[0] ? op_addae7_2_2_bufchan_buf :
                                   op_addae7_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_addae7_2_2_argbuf_r && op_addae7_2_2_bufchan_buf[0]))
        op_addae7_2_2_bufchan_buf <= 1'd0;
      else if (((! op_addae7_2_2_argbuf_r) && (! op_addae7_2_2_bufchan_buf[0])))
        op_addae7_2_2_bufchan_buf <= op_addae7_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addae7_2_destruct,MyDTInt_Int_Int) > [(op_addae7_2_1,MyDTInt_Int_Int),
                                                                      (op_addae7_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addae7_2_destruct_emitted;
  logic [1:0] op_addae7_2_destruct_done;
  assign op_addae7_2_1_d = (op_addae7_2_destruct_d[0] && (! op_addae7_2_destruct_emitted[0]));
  assign op_addae7_2_2_d = (op_addae7_2_destruct_d[0] && (! op_addae7_2_destruct_emitted[1]));
  assign op_addae7_2_destruct_done = (op_addae7_2_destruct_emitted | ({op_addae7_2_2_d[0],
                                                                       op_addae7_2_1_d[0]} & {op_addae7_2_2_r,
                                                                                              op_addae7_2_1_r}));
  assign op_addae7_2_destruct_r = (& op_addae7_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_2_destruct_emitted <= 2'd0;
    else
      op_addae7_2_destruct_emitted <= (op_addae7_2_destruct_r ? 2'd0 :
                                       op_addae7_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addae7_3_2,MyDTInt_Int_Int) > (op_addae7_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addae7_3_2_bufchan_d;
  logic op_addae7_3_2_bufchan_r;
  assign op_addae7_3_2_r = ((! op_addae7_3_2_bufchan_d[0]) || op_addae7_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_3_2_bufchan_d <= 1'd0;
    else
      if (op_addae7_3_2_r) op_addae7_3_2_bufchan_d <= op_addae7_3_2_d;
  MyDTInt_Int_Int_t op_addae7_3_2_bufchan_buf;
  assign op_addae7_3_2_bufchan_r = (! op_addae7_3_2_bufchan_buf[0]);
  assign op_addae7_3_2_argbuf_d = (op_addae7_3_2_bufchan_buf[0] ? op_addae7_3_2_bufchan_buf :
                                   op_addae7_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_addae7_3_2_argbuf_r && op_addae7_3_2_bufchan_buf[0]))
        op_addae7_3_2_bufchan_buf <= 1'd0;
      else if (((! op_addae7_3_2_argbuf_r) && (! op_addae7_3_2_bufchan_buf[0])))
        op_addae7_3_2_bufchan_buf <= op_addae7_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addae7_3_destruct,MyDTInt_Int_Int) > [(op_addae7_3_1,MyDTInt_Int_Int),
                                                                      (op_addae7_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addae7_3_destruct_emitted;
  logic [1:0] op_addae7_3_destruct_done;
  assign op_addae7_3_1_d = (op_addae7_3_destruct_d[0] && (! op_addae7_3_destruct_emitted[0]));
  assign op_addae7_3_2_d = (op_addae7_3_destruct_d[0] && (! op_addae7_3_destruct_emitted[1]));
  assign op_addae7_3_destruct_done = (op_addae7_3_destruct_emitted | ({op_addae7_3_2_d[0],
                                                                       op_addae7_3_1_d[0]} & {op_addae7_3_2_r,
                                                                                              op_addae7_3_1_r}));
  assign op_addae7_3_destruct_r = (& op_addae7_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_3_destruct_emitted <= 2'd0;
    else
      op_addae7_3_destruct_emitted <= (op_addae7_3_destruct_r ? 2'd0 :
                                       op_addae7_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addae7_4_destruct,MyDTInt_Int_Int) > (op_addae7_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addae7_4_destruct_bufchan_d;
  logic op_addae7_4_destruct_bufchan_r;
  assign op_addae7_4_destruct_r = ((! op_addae7_4_destruct_bufchan_d[0]) || op_addae7_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_addae7_4_destruct_r)
        op_addae7_4_destruct_bufchan_d <= op_addae7_4_destruct_d;
  MyDTInt_Int_Int_t op_addae7_4_destruct_bufchan_buf;
  assign op_addae7_4_destruct_bufchan_r = (! op_addae7_4_destruct_bufchan_buf[0]);
  assign op_addae7_4_1_argbuf_d = (op_addae7_4_destruct_bufchan_buf[0] ? op_addae7_4_destruct_bufchan_buf :
                                   op_addae7_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addae7_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_addae7_4_1_argbuf_r && op_addae7_4_destruct_bufchan_buf[0]))
        op_addae7_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_addae7_4_1_argbuf_r) && (! op_addae7_4_destruct_bufchan_buf[0])))
        op_addae7_4_destruct_bufchan_buf <= op_addae7_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeK_2_2,MyDTInt_Int_Int) > (op_addaeK_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeK_2_2_bufchan_d;
  logic op_addaeK_2_2_bufchan_r;
  assign op_addaeK_2_2_r = ((! op_addaeK_2_2_bufchan_d[0]) || op_addaeK_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_2_2_bufchan_d <= 1'd0;
    else
      if (op_addaeK_2_2_r) op_addaeK_2_2_bufchan_d <= op_addaeK_2_2_d;
  MyDTInt_Int_Int_t op_addaeK_2_2_bufchan_buf;
  assign op_addaeK_2_2_bufchan_r = (! op_addaeK_2_2_bufchan_buf[0]);
  assign op_addaeK_2_2_argbuf_d = (op_addaeK_2_2_bufchan_buf[0] ? op_addaeK_2_2_bufchan_buf :
                                   op_addaeK_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_addaeK_2_2_argbuf_r && op_addaeK_2_2_bufchan_buf[0]))
        op_addaeK_2_2_bufchan_buf <= 1'd0;
      else if (((! op_addaeK_2_2_argbuf_r) && (! op_addaeK_2_2_bufchan_buf[0])))
        op_addaeK_2_2_bufchan_buf <= op_addaeK_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addaeK_2_destruct,MyDTInt_Int_Int) > [(op_addaeK_2_1,MyDTInt_Int_Int),
                                                                      (op_addaeK_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addaeK_2_destruct_emitted;
  logic [1:0] op_addaeK_2_destruct_done;
  assign op_addaeK_2_1_d = (op_addaeK_2_destruct_d[0] && (! op_addaeK_2_destruct_emitted[0]));
  assign op_addaeK_2_2_d = (op_addaeK_2_destruct_d[0] && (! op_addaeK_2_destruct_emitted[1]));
  assign op_addaeK_2_destruct_done = (op_addaeK_2_destruct_emitted | ({op_addaeK_2_2_d[0],
                                                                       op_addaeK_2_1_d[0]} & {op_addaeK_2_2_r,
                                                                                              op_addaeK_2_1_r}));
  assign op_addaeK_2_destruct_r = (& op_addaeK_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_2_destruct_emitted <= 2'd0;
    else
      op_addaeK_2_destruct_emitted <= (op_addaeK_2_destruct_r ? 2'd0 :
                                       op_addaeK_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeK_3_2,MyDTInt_Int_Int) > (op_addaeK_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeK_3_2_bufchan_d;
  logic op_addaeK_3_2_bufchan_r;
  assign op_addaeK_3_2_r = ((! op_addaeK_3_2_bufchan_d[0]) || op_addaeK_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_3_2_bufchan_d <= 1'd0;
    else
      if (op_addaeK_3_2_r) op_addaeK_3_2_bufchan_d <= op_addaeK_3_2_d;
  MyDTInt_Int_Int_t op_addaeK_3_2_bufchan_buf;
  assign op_addaeK_3_2_bufchan_r = (! op_addaeK_3_2_bufchan_buf[0]);
  assign op_addaeK_3_2_argbuf_d = (op_addaeK_3_2_bufchan_buf[0] ? op_addaeK_3_2_bufchan_buf :
                                   op_addaeK_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_addaeK_3_2_argbuf_r && op_addaeK_3_2_bufchan_buf[0]))
        op_addaeK_3_2_bufchan_buf <= 1'd0;
      else if (((! op_addaeK_3_2_argbuf_r) && (! op_addaeK_3_2_bufchan_buf[0])))
        op_addaeK_3_2_bufchan_buf <= op_addaeK_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_addaeK_3_destruct,MyDTInt_Int_Int) > [(op_addaeK_3_1,MyDTInt_Int_Int),
                                                                      (op_addaeK_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_addaeK_3_destruct_emitted;
  logic [1:0] op_addaeK_3_destruct_done;
  assign op_addaeK_3_1_d = (op_addaeK_3_destruct_d[0] && (! op_addaeK_3_destruct_emitted[0]));
  assign op_addaeK_3_2_d = (op_addaeK_3_destruct_d[0] && (! op_addaeK_3_destruct_emitted[1]));
  assign op_addaeK_3_destruct_done = (op_addaeK_3_destruct_emitted | ({op_addaeK_3_2_d[0],
                                                                       op_addaeK_3_1_d[0]} & {op_addaeK_3_2_r,
                                                                                              op_addaeK_3_1_r}));
  assign op_addaeK_3_destruct_r = (& op_addaeK_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_3_destruct_emitted <= 2'd0;
    else
      op_addaeK_3_destruct_emitted <= (op_addaeK_3_destruct_r ? 2'd0 :
                                       op_addaeK_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_addaeK_4_destruct,MyDTInt_Int_Int) > (op_addaeK_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_addaeK_4_destruct_bufchan_d;
  logic op_addaeK_4_destruct_bufchan_r;
  assign op_addaeK_4_destruct_r = ((! op_addaeK_4_destruct_bufchan_d[0]) || op_addaeK_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_addaeK_4_destruct_r)
        op_addaeK_4_destruct_bufchan_d <= op_addaeK_4_destruct_d;
  MyDTInt_Int_Int_t op_addaeK_4_destruct_bufchan_buf;
  assign op_addaeK_4_destruct_bufchan_r = (! op_addaeK_4_destruct_bufchan_buf[0]);
  assign op_addaeK_4_1_argbuf_d = (op_addaeK_4_destruct_bufchan_buf[0] ? op_addaeK_4_destruct_bufchan_buf :
                                   op_addaeK_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_addaeK_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_addaeK_4_1_argbuf_r && op_addaeK_4_destruct_bufchan_buf[0]))
        op_addaeK_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_addaeK_4_1_argbuf_r) && (! op_addaeK_4_destruct_bufchan_buf[0])))
        op_addaeK_4_destruct_bufchan_buf <= op_addaeK_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1'aen_3_destruct,Pointer_QTree_Int) > (q1'aen_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \q1'aen_3_destruct_bufchan_d ;
  logic \q1'aen_3_destruct_bufchan_r ;
  assign \q1'aen_3_destruct_r  = ((! \q1'aen_3_destruct_bufchan_d [0]) || \q1'aen_3_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q1'aen_3_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q1'aen_3_destruct_r )
        \q1'aen_3_destruct_bufchan_d  <= \q1'aen_3_destruct_d ;
  Pointer_QTree_Int_t \q1'aen_3_destruct_bufchan_buf ;
  assign \q1'aen_3_destruct_bufchan_r  = (! \q1'aen_3_destruct_bufchan_buf [0]);
  assign \q1'aen_3_1_argbuf_d  = (\q1'aen_3_destruct_bufchan_buf [0] ? \q1'aen_3_destruct_bufchan_buf  :
                                  \q1'aen_3_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q1'aen_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q1'aen_3_1_argbuf_r  && \q1'aen_3_destruct_bufchan_buf [0]))
        \q1'aen_3_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q1'aen_3_1_argbuf_r ) && (! \q1'aen_3_destruct_bufchan_buf [0])))
        \q1'aen_3_destruct_bufchan_buf  <= \q1'aen_3_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a85_destruct,Pointer_QTree_Int) > (q1a85_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a85_destruct_bufchan_d;
  logic q1a85_destruct_bufchan_r;
  assign q1a85_destruct_r = ((! q1a85_destruct_bufchan_d[0]) || q1a85_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a85_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a85_destruct_r) q1a85_destruct_bufchan_d <= q1a85_destruct_d;
  Pointer_QTree_Int_t q1a85_destruct_bufchan_buf;
  assign q1a85_destruct_bufchan_r = (! q1a85_destruct_bufchan_buf[0]);
  assign q1a85_1_argbuf_d = (q1a85_destruct_bufchan_buf[0] ? q1a85_destruct_bufchan_buf :
                             q1a85_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a85_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a85_1_argbuf_r && q1a85_destruct_bufchan_buf[0]))
        q1a85_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a85_1_argbuf_r) && (! q1a85_destruct_bufchan_buf[0])))
        q1a85_destruct_bufchan_buf <= q1a85_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1ae8_3_destruct,Pointer_MaskQTree) > (q1ae8_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1ae8_3_destruct_bufchan_d;
  logic q1ae8_3_destruct_bufchan_r;
  assign q1ae8_3_destruct_r = ((! q1ae8_3_destruct_bufchan_d[0]) || q1ae8_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ae8_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ae8_3_destruct_r)
        q1ae8_3_destruct_bufchan_d <= q1ae8_3_destruct_d;
  Pointer_MaskQTree_t q1ae8_3_destruct_bufchan_buf;
  assign q1ae8_3_destruct_bufchan_r = (! q1ae8_3_destruct_bufchan_buf[0]);
  assign q1ae8_3_1_argbuf_d = (q1ae8_3_destruct_bufchan_buf[0] ? q1ae8_3_destruct_bufchan_buf :
                               q1ae8_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ae8_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ae8_3_1_argbuf_r && q1ae8_3_destruct_bufchan_buf[0]))
        q1ae8_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ae8_3_1_argbuf_r) && (! q1ae8_3_destruct_bufchan_buf[0])))
        q1ae8_3_destruct_bufchan_buf <= q1ae8_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1aeR_3_destruct,Pointer_QTree_Int) > (q1aeR_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1aeR_3_destruct_bufchan_d;
  logic q1aeR_3_destruct_bufchan_r;
  assign q1aeR_3_destruct_r = ((! q1aeR_3_destruct_bufchan_d[0]) || q1aeR_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aeR_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1aeR_3_destruct_r)
        q1aeR_3_destruct_bufchan_d <= q1aeR_3_destruct_d;
  Pointer_QTree_Int_t q1aeR_3_destruct_bufchan_buf;
  assign q1aeR_3_destruct_bufchan_r = (! q1aeR_3_destruct_bufchan_buf[0]);
  assign q1aeR_3_1_argbuf_d = (q1aeR_3_destruct_bufchan_buf[0] ? q1aeR_3_destruct_bufchan_buf :
                               q1aeR_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aeR_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1aeR_3_1_argbuf_r && q1aeR_3_destruct_bufchan_buf[0]))
        q1aeR_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1aeR_3_1_argbuf_r) && (! q1aeR_3_destruct_bufchan_buf[0])))
        q1aeR_3_destruct_bufchan_buf <= q1aeR_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1aey_3_destruct,Pointer_MaskQTree) > (q1aey_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1aey_3_destruct_bufchan_d;
  logic q1aey_3_destruct_bufchan_r;
  assign q1aey_3_destruct_r = ((! q1aey_3_destruct_bufchan_d[0]) || q1aey_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aey_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1aey_3_destruct_r)
        q1aey_3_destruct_bufchan_d <= q1aey_3_destruct_d;
  Pointer_MaskQTree_t q1aey_3_destruct_bufchan_buf;
  assign q1aey_3_destruct_bufchan_r = (! q1aey_3_destruct_bufchan_buf[0]);
  assign q1aey_3_1_argbuf_d = (q1aey_3_destruct_bufchan_buf[0] ? q1aey_3_destruct_bufchan_buf :
                               q1aey_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aey_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1aey_3_1_argbuf_r && q1aey_3_destruct_bufchan_buf[0]))
        q1aey_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1aey_3_1_argbuf_r) && (! q1aey_3_destruct_bufchan_buf[0])))
        q1aey_3_destruct_bufchan_buf <= q1aey_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2'aeo_2_destruct,Pointer_QTree_Int) > (q2'aeo_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \q2'aeo_2_destruct_bufchan_d ;
  logic \q2'aeo_2_destruct_bufchan_r ;
  assign \q2'aeo_2_destruct_r  = ((! \q2'aeo_2_destruct_bufchan_d [0]) || \q2'aeo_2_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q2'aeo_2_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q2'aeo_2_destruct_r )
        \q2'aeo_2_destruct_bufchan_d  <= \q2'aeo_2_destruct_d ;
  Pointer_QTree_Int_t \q2'aeo_2_destruct_bufchan_buf ;
  assign \q2'aeo_2_destruct_bufchan_r  = (! \q2'aeo_2_destruct_bufchan_buf [0]);
  assign \q2'aeo_2_1_argbuf_d  = (\q2'aeo_2_destruct_bufchan_buf [0] ? \q2'aeo_2_destruct_bufchan_buf  :
                                  \q2'aeo_2_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q2'aeo_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q2'aeo_2_1_argbuf_r  && \q2'aeo_2_destruct_bufchan_buf [0]))
        \q2'aeo_2_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q2'aeo_2_1_argbuf_r ) && (! \q2'aeo_2_destruct_bufchan_buf [0])))
        \q2'aeo_2_destruct_bufchan_buf  <= \q2'aeo_2_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a86_1_destruct,Pointer_QTree_Int) > (q2a86_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a86_1_destruct_bufchan_d;
  logic q2a86_1_destruct_bufchan_r;
  assign q2a86_1_destruct_r = ((! q2a86_1_destruct_bufchan_d[0]) || q2a86_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a86_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a86_1_destruct_r)
        q2a86_1_destruct_bufchan_d <= q2a86_1_destruct_d;
  Pointer_QTree_Int_t q2a86_1_destruct_bufchan_buf;
  assign q2a86_1_destruct_bufchan_r = (! q2a86_1_destruct_bufchan_buf[0]);
  assign q2a86_1_1_argbuf_d = (q2a86_1_destruct_bufchan_buf[0] ? q2a86_1_destruct_bufchan_buf :
                               q2a86_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a86_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a86_1_1_argbuf_r && q2a86_1_destruct_bufchan_buf[0]))
        q2a86_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a86_1_1_argbuf_r) && (! q2a86_1_destruct_bufchan_buf[0])))
        q2a86_1_destruct_bufchan_buf <= q2a86_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2ae9_2_destruct,Pointer_MaskQTree) > (q2ae9_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2ae9_2_destruct_bufchan_d;
  logic q2ae9_2_destruct_bufchan_r;
  assign q2ae9_2_destruct_r = ((! q2ae9_2_destruct_bufchan_d[0]) || q2ae9_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ae9_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2ae9_2_destruct_r)
        q2ae9_2_destruct_bufchan_d <= q2ae9_2_destruct_d;
  Pointer_MaskQTree_t q2ae9_2_destruct_bufchan_buf;
  assign q2ae9_2_destruct_bufchan_r = (! q2ae9_2_destruct_bufchan_buf[0]);
  assign q2ae9_2_1_argbuf_d = (q2ae9_2_destruct_bufchan_buf[0] ? q2ae9_2_destruct_bufchan_buf :
                               q2ae9_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ae9_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2ae9_2_1_argbuf_r && q2ae9_2_destruct_bufchan_buf[0]))
        q2ae9_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2ae9_2_1_argbuf_r) && (! q2ae9_2_destruct_bufchan_buf[0])))
        q2ae9_2_destruct_bufchan_buf <= q2ae9_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2aeS_2_destruct,Pointer_QTree_Int) > (q2aeS_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2aeS_2_destruct_bufchan_d;
  logic q2aeS_2_destruct_bufchan_r;
  assign q2aeS_2_destruct_r = ((! q2aeS_2_destruct_bufchan_d[0]) || q2aeS_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aeS_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2aeS_2_destruct_r)
        q2aeS_2_destruct_bufchan_d <= q2aeS_2_destruct_d;
  Pointer_QTree_Int_t q2aeS_2_destruct_bufchan_buf;
  assign q2aeS_2_destruct_bufchan_r = (! q2aeS_2_destruct_bufchan_buf[0]);
  assign q2aeS_2_1_argbuf_d = (q2aeS_2_destruct_bufchan_buf[0] ? q2aeS_2_destruct_bufchan_buf :
                               q2aeS_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aeS_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2aeS_2_1_argbuf_r && q2aeS_2_destruct_bufchan_buf[0]))
        q2aeS_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2aeS_2_1_argbuf_r) && (! q2aeS_2_destruct_bufchan_buf[0])))
        q2aeS_2_destruct_bufchan_buf <= q2aeS_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2aez_2_destruct,Pointer_MaskQTree) > (q2aez_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2aez_2_destruct_bufchan_d;
  logic q2aez_2_destruct_bufchan_r;
  assign q2aez_2_destruct_r = ((! q2aez_2_destruct_bufchan_d[0]) || q2aez_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aez_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2aez_2_destruct_r)
        q2aez_2_destruct_bufchan_d <= q2aez_2_destruct_d;
  Pointer_MaskQTree_t q2aez_2_destruct_bufchan_buf;
  assign q2aez_2_destruct_bufchan_r = (! q2aez_2_destruct_bufchan_buf[0]);
  assign q2aez_2_1_argbuf_d = (q2aez_2_destruct_bufchan_buf[0] ? q2aez_2_destruct_bufchan_buf :
                               q2aez_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aez_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2aez_2_1_argbuf_r && q2aez_2_destruct_bufchan_buf[0]))
        q2aez_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2aez_2_1_argbuf_r) && (! q2aez_2_destruct_bufchan_buf[0])))
        q2aez_2_destruct_bufchan_buf <= q2aez_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3'aep_1_destruct,Pointer_QTree_Int) > (q3'aep_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \q3'aep_1_destruct_bufchan_d ;
  logic \q3'aep_1_destruct_bufchan_r ;
  assign \q3'aep_1_destruct_r  = ((! \q3'aep_1_destruct_bufchan_d [0]) || \q3'aep_1_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q3'aep_1_destruct_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\q3'aep_1_destruct_r )
        \q3'aep_1_destruct_bufchan_d  <= \q3'aep_1_destruct_d ;
  Pointer_QTree_Int_t \q3'aep_1_destruct_bufchan_buf ;
  assign \q3'aep_1_destruct_bufchan_r  = (! \q3'aep_1_destruct_bufchan_buf [0]);
  assign \q3'aep_1_1_argbuf_d  = (\q3'aep_1_destruct_bufchan_buf [0] ? \q3'aep_1_destruct_bufchan_buf  :
                                  \q3'aep_1_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \q3'aep_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q3'aep_1_1_argbuf_r  && \q3'aep_1_destruct_bufchan_buf [0]))
        \q3'aep_1_destruct_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q3'aep_1_1_argbuf_r ) && (! \q3'aep_1_destruct_bufchan_buf [0])))
        \q3'aep_1_destruct_bufchan_buf  <= \q3'aep_1_destruct_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a87_2_destruct,Pointer_QTree_Int) > (q3a87_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a87_2_destruct_bufchan_d;
  logic q3a87_2_destruct_bufchan_r;
  assign q3a87_2_destruct_r = ((! q3a87_2_destruct_bufchan_d[0]) || q3a87_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a87_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a87_2_destruct_r)
        q3a87_2_destruct_bufchan_d <= q3a87_2_destruct_d;
  Pointer_QTree_Int_t q3a87_2_destruct_bufchan_buf;
  assign q3a87_2_destruct_bufchan_r = (! q3a87_2_destruct_bufchan_buf[0]);
  assign q3a87_2_1_argbuf_d = (q3a87_2_destruct_bufchan_buf[0] ? q3a87_2_destruct_bufchan_buf :
                               q3a87_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a87_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a87_2_1_argbuf_r && q3a87_2_destruct_bufchan_buf[0]))
        q3a87_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a87_2_1_argbuf_r) && (! q3a87_2_destruct_bufchan_buf[0])))
        q3a87_2_destruct_bufchan_buf <= q3a87_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3aeA_1_destruct,Pointer_MaskQTree) > (q3aeA_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3aeA_1_destruct_bufchan_d;
  logic q3aeA_1_destruct_bufchan_r;
  assign q3aeA_1_destruct_r = ((! q3aeA_1_destruct_bufchan_d[0]) || q3aeA_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aeA_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aeA_1_destruct_r)
        q3aeA_1_destruct_bufchan_d <= q3aeA_1_destruct_d;
  Pointer_MaskQTree_t q3aeA_1_destruct_bufchan_buf;
  assign q3aeA_1_destruct_bufchan_r = (! q3aeA_1_destruct_bufchan_buf[0]);
  assign q3aeA_1_1_argbuf_d = (q3aeA_1_destruct_bufchan_buf[0] ? q3aeA_1_destruct_bufchan_buf :
                               q3aeA_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aeA_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aeA_1_1_argbuf_r && q3aeA_1_destruct_bufchan_buf[0]))
        q3aeA_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aeA_1_1_argbuf_r) && (! q3aeA_1_destruct_bufchan_buf[0])))
        q3aeA_1_destruct_bufchan_buf <= q3aeA_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3aeT_1_destruct,Pointer_QTree_Int) > (q3aeT_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3aeT_1_destruct_bufchan_d;
  logic q3aeT_1_destruct_bufchan_r;
  assign q3aeT_1_destruct_r = ((! q3aeT_1_destruct_bufchan_d[0]) || q3aeT_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aeT_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aeT_1_destruct_r)
        q3aeT_1_destruct_bufchan_d <= q3aeT_1_destruct_d;
  Pointer_QTree_Int_t q3aeT_1_destruct_bufchan_buf;
  assign q3aeT_1_destruct_bufchan_r = (! q3aeT_1_destruct_bufchan_buf[0]);
  assign q3aeT_1_1_argbuf_d = (q3aeT_1_destruct_bufchan_buf[0] ? q3aeT_1_destruct_bufchan_buf :
                               q3aeT_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aeT_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aeT_1_1_argbuf_r && q3aeT_1_destruct_bufchan_buf[0]))
        q3aeT_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aeT_1_1_argbuf_r) && (! q3aeT_1_destruct_bufchan_buf[0])))
        q3aeT_1_destruct_bufchan_buf <= q3aeT_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3aea_1_destruct,Pointer_MaskQTree) > (q3aea_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3aea_1_destruct_bufchan_d;
  logic q3aea_1_destruct_bufchan_r;
  assign q3aea_1_destruct_r = ((! q3aea_1_destruct_bufchan_d[0]) || q3aea_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aea_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aea_1_destruct_r)
        q3aea_1_destruct_bufchan_d <= q3aea_1_destruct_d;
  Pointer_MaskQTree_t q3aea_1_destruct_bufchan_buf;
  assign q3aea_1_destruct_bufchan_r = (! q3aea_1_destruct_bufchan_buf[0]);
  assign q3aea_1_1_argbuf_d = (q3aea_1_destruct_bufchan_buf[0] ? q3aea_1_destruct_bufchan_buf :
                               q3aea_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aea_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aea_1_1_argbuf_r && q3aea_1_destruct_bufchan_buf[0]))
        q3aea_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aea_1_1_argbuf_r) && (! q3aea_1_destruct_bufchan_buf[0])))
        q3aea_1_destruct_bufchan_buf <= q3aea_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4'aex_1,Pointer_QTree_Int) > (q4'aex_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \q4'aex_1_bufchan_d ;
  logic \q4'aex_1_bufchan_r ;
  assign \q4'aex_1_r  = ((! \q4'aex_1_bufchan_d [0]) || \q4'aex_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'aex_1_bufchan_d  <= {16'd0, 1'd0};
    else if (\q4'aex_1_r ) \q4'aex_1_bufchan_d  <= \q4'aex_1_d ;
  Pointer_QTree_Int_t \q4'aex_1_bufchan_buf ;
  assign \q4'aex_1_bufchan_r  = (! \q4'aex_1_bufchan_buf [0]);
  assign \q4'aex_1_argbuf_d  = (\q4'aex_1_bufchan_buf [0] ? \q4'aex_1_bufchan_buf  :
                                \q4'aex_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'aex_1_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\q4'aex_1_argbuf_r  && \q4'aex_1_bufchan_buf [0]))
        \q4'aex_1_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \q4'aex_1_argbuf_r ) && (! \q4'aex_1_bufchan_buf [0])))
        \q4'aex_1_bufchan_buf  <= \q4'aex_1_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (q4'aex_goMux_mux,Pointer_QTree_Int) > [(q4'aex_1,Pointer_QTree_Int),
                                                                      (q4'aex_2,Pointer_QTree_Int)] */
  logic [1:0] \q4'aex_goMux_mux_emitted ;
  logic [1:0] \q4'aex_goMux_mux_done ;
  assign \q4'aex_1_d  = {\q4'aex_goMux_mux_d [16:1],
                         (\q4'aex_goMux_mux_d [0] && (! \q4'aex_goMux_mux_emitted [0]))};
  assign \q4'aex_2_d  = {\q4'aex_goMux_mux_d [16:1],
                         (\q4'aex_goMux_mux_d [0] && (! \q4'aex_goMux_mux_emitted [1]))};
  assign \q4'aex_goMux_mux_done  = (\q4'aex_goMux_mux_emitted  | ({\q4'aex_2_d [0],
                                                                   \q4'aex_1_d [0]} & {\q4'aex_2_r ,
                                                                                       \q4'aex_1_r }));
  assign \q4'aex_goMux_mux_r  = (& \q4'aex_goMux_mux_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \q4'aex_goMux_mux_emitted  <= 2'd0;
    else
      \q4'aex_goMux_mux_emitted  <= (\q4'aex_goMux_mux_r  ? 2'd0 :
                                     \q4'aex_goMux_mux_done );
  
  /* buf (Ty Pointer_QTree_Int) : (q4a88_3_destruct,Pointer_QTree_Int) > (q4a88_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a88_3_destruct_bufchan_d;
  logic q4a88_3_destruct_bufchan_r;
  assign q4a88_3_destruct_r = ((! q4a88_3_destruct_bufchan_d[0]) || q4a88_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a88_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a88_3_destruct_r)
        q4a88_3_destruct_bufchan_d <= q4a88_3_destruct_d;
  Pointer_QTree_Int_t q4a88_3_destruct_bufchan_buf;
  assign q4a88_3_destruct_bufchan_r = (! q4a88_3_destruct_bufchan_buf[0]);
  assign q4a88_3_1_argbuf_d = (q4a88_3_destruct_bufchan_buf[0] ? q4a88_3_destruct_bufchan_buf :
                               q4a88_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a88_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a88_3_1_argbuf_r && q4a88_3_destruct_bufchan_buf[0]))
        q4a88_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a88_3_1_argbuf_r) && (! q4a88_3_destruct_bufchan_buf[0])))
        q4a88_3_destruct_bufchan_buf <= q4a88_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q4aew_goMux_mux,Pointer_MaskQTree) > (q4aew_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q4aew_goMux_mux_bufchan_d;
  logic q4aew_goMux_mux_bufchan_r;
  assign q4aew_goMux_mux_r = ((! q4aew_goMux_mux_bufchan_d[0]) || q4aew_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4aew_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4aew_goMux_mux_r)
        q4aew_goMux_mux_bufchan_d <= q4aew_goMux_mux_d;
  Pointer_MaskQTree_t q4aew_goMux_mux_bufchan_buf;
  assign q4aew_goMux_mux_bufchan_r = (! q4aew_goMux_mux_bufchan_buf[0]);
  assign q4aew_1_argbuf_d = (q4aew_goMux_mux_bufchan_buf[0] ? q4aew_goMux_mux_bufchan_buf :
                             q4aew_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4aew_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4aew_1_argbuf_r && q4aew_goMux_mux_bufchan_buf[0]))
        q4aew_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4aew_1_argbuf_r) && (! q4aew_goMux_mux_bufchan_buf[0])))
        q4aew_goMux_mux_bufchan_buf <= q4aew_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int) > (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) */
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                             1'd0};
    else
      if (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf :
                                                           readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                               1'd0};
    else
      if ((readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
      else if (((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) > [(lizzieLet46_1,CT$wnnz_Int),
                                                                                      (lizzieLet46_2,CT$wnnz_Int),
                                                                                      (lizzieLet46_3,CT$wnnz_Int),
                                                                                      (lizzieLet46_4,CT$wnnz_Int)] */
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet46_1_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet46_2_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet46_3_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet46_4_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet46_4_d[0],
                                                                                                                       lizzieLet46_3_d[0],
                                                                                                                       lizzieLet46_2_d[0],
                                                                                                                       lizzieLet46_1_d[0]} & {lizzieLet46_4_r,
                                                                                                                                              lizzieLet46_3_r,
                                                                                                                                              lizzieLet46_2_r,
                                                                                                                                              lizzieLet46_1_r}));
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTf'''''''''_f'''''''''_Int) : (readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf,CTf'''''''''_f'''''''''_Int) > (readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb,CTf'''''''''_f'''''''''_Int) */
  \CTf'''''''''_f'''''''''_Int_t  \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d  <= {115'd0,
                                                                                 1'd0};
    else
      if (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_r )
        \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_d ;
  \CTf'''''''''_f'''''''''_Int_t  \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  :
                                                                               \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                   1'd0};
    else
      if ((\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {115'd0,
                                                                                     1'd0};
      else if (((! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf'''''''''_f'''''''''_Int) : (readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb,CTf'''''''''_f'''''''''_Int) > [(lizzieLet50_1,CTf'''''''''_f'''''''''_Int),
                                                                                                                                        (lizzieLet50_2,CTf'''''''''_f'''''''''_Int),
                                                                                                                                        (lizzieLet50_3,CTf'''''''''_f'''''''''_Int),
                                                                                                                                        (lizzieLet50_4,CTf'''''''''_f'''''''''_Int)] */
  logic [3:0] \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet50_1_d = {\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet50_2_d = {\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet50_3_d = {\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet50_4_d = {\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet50_4_d[0],
                                                                                                                                                               lizzieLet50_3_d[0],
                                                                                                                                                               lizzieLet50_2_d[0],
                                                                                                                                                               lizzieLet50_1_d[0]} & {lizzieLet50_4_r,
                                                                                                                                                                                      lizzieLet50_3_r,
                                                                                                                                                                                      lizzieLet50_2_r,
                                                                                                                                                                                      lizzieLet50_1_r}));
  assign \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                                   \readPointer_CTf'''''''''_f'''''''''_Intscfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf'_f'_Int) : (readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf,CTf'_f'_Int) > (readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb,CTf'_f'_Int) */
  \CTf'_f'_Int_t  \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d  <= {115'd0,
                                                                 1'd0};
    else
      if (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_r )
        \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_d ;
  \CTf'_f'_Int_t  \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf  :
                                                               \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf  <= {115'd0,
                                                                   1'd0};
    else
      if ((\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf  <= {115'd0,
                                                                     1'd0};
      else if (((! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf'_f'_Int) : (readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb,CTf'_f'_Int) > [(lizzieLet55_1,CTf'_f'_Int),
                                                                                        (lizzieLet55_2,CTf'_f'_Int),
                                                                                        (lizzieLet55_3,CTf'_f'_Int),
                                                                                        (lizzieLet55_4,CTf'_f'_Int)] */
  logic [3:0] \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet55_1_d = {\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet55_2_d = {\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet55_3_d = {\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet55_4_d = {\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [115:1],
                            (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet55_4_d[0],
                                                                                                                               lizzieLet55_3_d[0],
                                                                                                                               lizzieLet55_2_d[0],
                                                                                                                               lizzieLet55_1_d[0]} & {lizzieLet55_4_r,
                                                                                                                                                      lizzieLet55_3_r,
                                                                                                                                                      lizzieLet55_2_r,
                                                                                                                                                      lizzieLet55_1_r}));
  assign \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                   \readPointer_CTf'_f'_Intscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty CTf_f_Int) : (readPointer_CTf_f_Intscfarg_0_3_1_argbuf,CTf_f_Int) > (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb,CTf_f_Int) */
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d;
  logic readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_r;
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_r = ((! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d[0]) || readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d <= {163'd0,
                                                             1'd0};
    else
      if (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_r)
        readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d <= readPointer_CTf_f_Intscfarg_0_3_1_argbuf_d;
  CTf_f_Int_t readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf;
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_r = (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d = (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf[0] ? readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf :
                                                           readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf <= {163'd0,
                                                               1'd0};
    else
      if ((readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_r && readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf[0]))
        readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf <= {163'd0,
                                                                 1'd0};
      else if (((! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_r) && (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf[0])))
        readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_buf <= readPointer_CTf_f_Intscfarg_0_3_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf_f_Int) : (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb,CTf_f_Int) > [(lizzieLet60_1,CTf_f_Int),
                                                                                  (lizzieLet60_2,CTf_f_Int),
                                                                                  (lizzieLet60_3,CTf_f_Int),
                                                                                  (lizzieLet60_4,CTf_f_Int)] */
  logic [3:0] readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_done;
  assign lizzieLet60_1_d = {readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet60_2_d = {readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet60_3_d = {readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet60_4_d = {readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[163:1],
                            (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_done = (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted | ({lizzieLet60_4_d[0],
                                                                                                                       lizzieLet60_3_d[0],
                                                                                                                       lizzieLet60_2_d[0],
                                                                                                                       lizzieLet60_1_d[0]} & {lizzieLet60_4_r,
                                                                                                                                              lizzieLet60_3_r,
                                                                                                                                              lizzieLet60_2_r,
                                                                                                                                              lizzieLet60_1_r}));
  assign readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_r = (& readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_emitted <= (readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CTf_f_Intscfarg_0_3_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreem1ae3_1_argbuf,MaskQTree) > (readPointer_MaskQTreem1ae3_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreem1ae3_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreem1ae3_1_argbuf_r = ((! readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreem1ae3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreem1ae3_1_argbuf_r)
        readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d <= readPointer_MaskQTreem1ae3_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreem1ae3_1_argbuf_bufchan_r = (! readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreem1ae3_1_argbuf_rwb_d = (readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf :
                                                      readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreem1ae3_1_argbuf_rwb_r && readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreem1ae3_1_argbuf_rwb_r) && (! readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreem1ae3_1_argbuf_bufchan_buf <= readPointer_MaskQTreem1ae3_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreem1ae3_1_argbuf_rwb,MaskQTree) > [(lizzieLet24_1,MaskQTree),
                                                                             (lizzieLet24_2,MaskQTree),
                                                                             (lizzieLet24_3,MaskQTree),
                                                                             (lizzieLet24_4,MaskQTree),
                                                                             (lizzieLet24_5,MaskQTree),
                                                                             (lizzieLet24_6,MaskQTree),
                                                                             (lizzieLet24_7,MaskQTree),
                                                                             (lizzieLet24_8,MaskQTree),
                                                                             (lizzieLet24_9,MaskQTree),
                                                                             (lizzieLet24_10,MaskQTree)] */
  logic [9:0] readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted;
  logic [9:0] readPointer_MaskQTreem1ae3_1_argbuf_rwb_done;
  assign lizzieLet24_1_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet24_2_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet24_3_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet24_4_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet24_5_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet24_6_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet24_7_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet24_8_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet24_9_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                            (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[8]))};
  assign lizzieLet24_10_d = {readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[66:1],
                             (readPointer_MaskQTreem1ae3_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted[9]))};
  assign readPointer_MaskQTreem1ae3_1_argbuf_rwb_done = (readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted | ({lizzieLet24_10_d[0],
                                                                                                             lizzieLet24_9_d[0],
                                                                                                             lizzieLet24_8_d[0],
                                                                                                             lizzieLet24_7_d[0],
                                                                                                             lizzieLet24_6_d[0],
                                                                                                             lizzieLet24_5_d[0],
                                                                                                             lizzieLet24_4_d[0],
                                                                                                             lizzieLet24_3_d[0],
                                                                                                             lizzieLet24_2_d[0],
                                                                                                             lizzieLet24_1_d[0]} & {lizzieLet24_10_r,
                                                                                                                                    lizzieLet24_9_r,
                                                                                                                                    lizzieLet24_8_r,
                                                                                                                                    lizzieLet24_7_r,
                                                                                                                                    lizzieLet24_6_r,
                                                                                                                                    lizzieLet24_5_r,
                                                                                                                                    lizzieLet24_4_r,
                                                                                                                                    lizzieLet24_3_r,
                                                                                                                                    lizzieLet24_2_r,
                                                                                                                                    lizzieLet24_1_r}));
  assign readPointer_MaskQTreem1ae3_1_argbuf_rwb_r = (& readPointer_MaskQTreem1ae3_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted <= 10'd0;
    else
      readPointer_MaskQTreem1ae3_1_argbuf_rwb_emitted <= (readPointer_MaskQTreem1ae3_1_argbuf_rwb_r ? 10'd0 :
                                                          readPointer_MaskQTreem1ae3_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreeq4aew_1_argbuf,MaskQTree) > (readPointer_MaskQTreeq4aew_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreeq4aew_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreeq4aew_1_argbuf_r = ((! readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreeq4aew_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreeq4aew_1_argbuf_r)
        readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d <= readPointer_MaskQTreeq4aew_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreeq4aew_1_argbuf_bufchan_r = (! readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreeq4aew_1_argbuf_rwb_d = (readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf :
                                                      readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreeq4aew_1_argbuf_rwb_r && readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreeq4aew_1_argbuf_rwb_r) && (! readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreeq4aew_1_argbuf_bufchan_buf <= readPointer_MaskQTreeq4aew_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreeq4aew_1_argbuf_rwb,MaskQTree) > [(lizzieLet6_1,MaskQTree),
                                                                             (lizzieLet6_2,MaskQTree),
                                                                             (lizzieLet6_3,MaskQTree),
                                                                             (lizzieLet6_4,MaskQTree),
                                                                             (lizzieLet6_5,MaskQTree),
                                                                             (lizzieLet6_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreeq4aew_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[66:1],
                           (readPointer_MaskQTreeq4aew_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreeq4aew_1_argbuf_rwb_done = (readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted | ({lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_MaskQTreeq4aew_1_argbuf_rwb_r = (& readPointer_MaskQTreeq4aew_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreeq4aew_1_argbuf_rwb_emitted <= (readPointer_MaskQTreeq4aew_1_argbuf_rwb_r ? 6'd0 :
                                                          readPointer_MaskQTreeq4aew_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2ae4_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2ae4_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2ae4_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2ae4_1_argbuf_r = ((! readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2ae4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2ae4_1_argbuf_r)
        readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d <= readPointer_QTree_Intm2ae4_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2ae4_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2ae4_1_argbuf_rwb_d = (readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2ae4_1_argbuf_rwb_r && readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2ae4_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2ae4_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2ae4_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2aeH_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2aeH_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2aeH_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2aeH_1_argbuf_r = ((! readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2aeH_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2aeH_1_argbuf_r)
        readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d <= readPointer_QTree_Intm2aeH_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2aeH_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2aeH_1_argbuf_rwb_d = (readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2aeH_1_argbuf_rwb_r && readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2aeH_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2aeH_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2aeH_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm2aeH_1_argbuf_rwb,QTree_Int) > [(lizzieLet13_1,QTree_Int),
                                                                             (lizzieLet13_2,QTree_Int),
                                                                             (lizzieLet13_3,QTree_Int),
                                                                             (lizzieLet13_4,QTree_Int),
                                                                             (lizzieLet13_5,QTree_Int),
                                                                             (lizzieLet13_6,QTree_Int),
                                                                             (lizzieLet13_7,QTree_Int),
                                                                             (lizzieLet13_8,QTree_Int),
                                                                             (lizzieLet13_9,QTree_Int)] */
  logic [8:0] readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Intm2aeH_1_argbuf_rwb_done;
  assign lizzieLet13_1_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet13_2_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet13_3_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet13_4_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet13_5_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet13_6_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet13_7_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet13_8_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet13_9_d = {readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intm2aeH_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Intm2aeH_1_argbuf_rwb_done = (readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted | ({lizzieLet13_9_d[0],
                                                                                                             lizzieLet13_8_d[0],
                                                                                                             lizzieLet13_7_d[0],
                                                                                                             lizzieLet13_6_d[0],
                                                                                                             lizzieLet13_5_d[0],
                                                                                                             lizzieLet13_4_d[0],
                                                                                                             lizzieLet13_3_d[0],
                                                                                                             lizzieLet13_2_d[0],
                                                                                                             lizzieLet13_1_d[0]} & {lizzieLet13_9_r,
                                                                                                                                    lizzieLet13_8_r,
                                                                                                                                    lizzieLet13_7_r,
                                                                                                                                    lizzieLet13_6_r,
                                                                                                                                    lizzieLet13_5_r,
                                                                                                                                    lizzieLet13_4_r,
                                                                                                                                    lizzieLet13_3_r,
                                                                                                                                    lizzieLet13_2_r,
                                                                                                                                    lizzieLet13_1_r}));
  assign readPointer_QTree_Intm2aeH_1_argbuf_rwb_r = (& readPointer_QTree_Intm2aeH_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Intm2aeH_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm2aeH_1_argbuf_rwb_r ? 9'd0 :
                                                          readPointer_QTree_Intm2aeH_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm3ae5_1_argbuf,QTree_Int) > (readPointer_QTree_Intm3ae5_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm3ae5_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm3ae5_1_argbuf_r = ((! readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm3ae5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm3ae5_1_argbuf_r)
        readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d <= readPointer_QTree_Intm3ae5_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm3ae5_1_argbuf_bufchan_r = (! readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm3ae5_1_argbuf_rwb_d = (readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm3ae5_1_argbuf_rwb_r && readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm3ae5_1_argbuf_rwb_r) && (! readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm3ae5_1_argbuf_bufchan_buf <= readPointer_QTree_Intm3ae5_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm3aeI_1_argbuf,QTree_Int) > (readPointer_QTree_Intm3aeI_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm3aeI_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm3aeI_1_argbuf_r = ((! readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm3aeI_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm3aeI_1_argbuf_r)
        readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d <= readPointer_QTree_Intm3aeI_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm3aeI_1_argbuf_bufchan_r = (! readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm3aeI_1_argbuf_rwb_d = (readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm3aeI_1_argbuf_rwb_r && readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm3aeI_1_argbuf_rwb_r) && (! readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm3aeI_1_argbuf_bufchan_buf <= readPointer_QTree_Intm3aeI_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intq4'aex_1_argbuf,QTree_Int) > (readPointer_QTree_Intq4'aex_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d ;
  logic \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_r ;
  assign \readPointer_QTree_Intq4'aex_1_argbuf_r  = ((! \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d [0]) || \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d  <= {66'd0, 1'd0};
    else
      if (\readPointer_QTree_Intq4'aex_1_argbuf_r )
        \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d  <= \readPointer_QTree_Intq4'aex_1_argbuf_d ;
  QTree_Int_t \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf ;
  assign \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_r  = (! \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf [0]);
  assign \readPointer_QTree_Intq4'aex_1_argbuf_rwb_d  = (\readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf [0] ? \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf  :
                                                         \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf  <= {66'd0,
                                                             1'd0};
    else
      if ((\readPointer_QTree_Intq4'aex_1_argbuf_rwb_r  && \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf [0]))
        \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf  <= {66'd0,
                                                               1'd0};
      else if (((! \readPointer_QTree_Intq4'aex_1_argbuf_rwb_r ) && (! \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf [0])))
        \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_buf  <= \readPointer_QTree_Intq4'aex_1_argbuf_bufchan_d ;
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntwsjQ_1_1_argbuf,QTree_Int) > (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_r = ((! readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntwsjQ_1_1_argbuf_r)
        readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d <= readPointer_QTree_IntwsjQ_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_r = (! readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d = (readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_r && readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_r) && (! readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_buf <= readPointer_QTree_IntwsjQ_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_done = (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_r = (& readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_emitted <= (readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_IntwsjQ_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (sc_0_11_destruct,Pointer_CTf'''''''''_f'''''''''_Int) > (sc_0_11_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_11_destruct_bufchan_d;
  logic sc_0_11_destruct_bufchan_r;
  assign sc_0_11_destruct_r = ((! sc_0_11_destruct_bufchan_d[0]) || sc_0_11_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_11_destruct_r)
        sc_0_11_destruct_bufchan_d <= sc_0_11_destruct_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  sc_0_11_destruct_bufchan_buf;
  assign sc_0_11_destruct_bufchan_r = (! sc_0_11_destruct_bufchan_buf[0]);
  assign sc_0_11_1_argbuf_d = (sc_0_11_destruct_bufchan_buf[0] ? sc_0_11_destruct_bufchan_buf :
                               sc_0_11_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_11_1_argbuf_r && sc_0_11_destruct_bufchan_buf[0]))
        sc_0_11_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_11_1_argbuf_r) && (! sc_0_11_destruct_bufchan_buf[0])))
        sc_0_11_destruct_bufchan_buf <= sc_0_11_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (sc_0_15_destruct,Pointer_CTf'_f'_Int) > (sc_0_15_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  sc_0_15_destruct_bufchan_d;
  logic sc_0_15_destruct_bufchan_r;
  assign sc_0_15_destruct_r = ((! sc_0_15_destruct_bufchan_d[0]) || sc_0_15_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_15_destruct_r)
        sc_0_15_destruct_bufchan_d <= sc_0_15_destruct_d;
  \Pointer_CTf'_f'_Int_t  sc_0_15_destruct_bufchan_buf;
  assign sc_0_15_destruct_bufchan_r = (! sc_0_15_destruct_bufchan_buf[0]);
  assign sc_0_15_1_argbuf_d = (sc_0_15_destruct_bufchan_buf[0] ? sc_0_15_destruct_bufchan_buf :
                               sc_0_15_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_15_1_argbuf_r && sc_0_15_destruct_bufchan_buf[0]))
        sc_0_15_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_15_1_argbuf_r) && (! sc_0_15_destruct_bufchan_buf[0])))
        sc_0_15_destruct_bufchan_buf <= sc_0_15_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (sc_0_19_destruct,Pointer_CTf_f_Int) > (sc_0_19_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t sc_0_19_destruct_bufchan_d;
  logic sc_0_19_destruct_bufchan_r;
  assign sc_0_19_destruct_r = ((! sc_0_19_destruct_bufchan_d[0]) || sc_0_19_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_19_destruct_r)
        sc_0_19_destruct_bufchan_d <= sc_0_19_destruct_d;
  Pointer_CTf_f_Int_t sc_0_19_destruct_bufchan_buf;
  assign sc_0_19_destruct_bufchan_r = (! sc_0_19_destruct_bufchan_buf[0]);
  assign sc_0_19_1_argbuf_d = (sc_0_19_destruct_bufchan_buf[0] ? sc_0_19_destruct_bufchan_buf :
                               sc_0_19_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_19_1_argbuf_r && sc_0_19_destruct_bufchan_buf[0]))
        sc_0_19_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_19_1_argbuf_r) && (! sc_0_19_destruct_bufchan_buf[0])))
        sc_0_19_destruct_bufchan_buf <= sc_0_19_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (sc_0_7_destruct,Pointer_CT$wnnz_Int) > (sc_0_7_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_d;
  logic sc_0_7_destruct_bufchan_r;
  assign sc_0_7_destruct_r = ((! sc_0_7_destruct_bufchan_d[0]) || sc_0_7_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_7_destruct_r)
        sc_0_7_destruct_bufchan_d <= sc_0_7_destruct_d;
  Pointer_CT$wnnz_Int_t sc_0_7_destruct_bufchan_buf;
  assign sc_0_7_destruct_bufchan_r = (! sc_0_7_destruct_bufchan_buf[0]);
  assign sc_0_7_1_argbuf_d = (sc_0_7_destruct_bufchan_buf[0] ? sc_0_7_destruct_bufchan_buf :
                              sc_0_7_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_7_1_argbuf_r && sc_0_7_destruct_bufchan_buf[0]))
        sc_0_7_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_7_1_argbuf_r) && (! sc_0_7_destruct_bufchan_buf[0])))
        sc_0_7_destruct_bufchan_buf <= sc_0_7_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (scfarg_0_1_goMux_mux,Pointer_CTf'''''''''_f'''''''''_Int) > (scfarg_0_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (scfarg_0_2_goMux_mux,Pointer_CTf'_f'_Int) > (scfarg_0_2_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTf'_f'_Int_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (scfarg_0_3_goMux_mux,Pointer_CTf_f_Int) > (scfarg_0_3_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t scfarg_0_3_goMux_mux_bufchan_d;
  logic scfarg_0_3_goMux_mux_bufchan_r;
  assign scfarg_0_3_goMux_mux_r = ((! scfarg_0_3_goMux_mux_bufchan_d[0]) || scfarg_0_3_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_3_goMux_mux_r)
        scfarg_0_3_goMux_mux_bufchan_d <= scfarg_0_3_goMux_mux_d;
  Pointer_CTf_f_Int_t scfarg_0_3_goMux_mux_bufchan_buf;
  assign scfarg_0_3_goMux_mux_bufchan_r = (! scfarg_0_3_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_3_1_argbuf_d = (scfarg_0_3_goMux_mux_bufchan_buf[0] ? scfarg_0_3_goMux_mux_bufchan_buf :
                                  scfarg_0_3_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_3_1_argbuf_r && scfarg_0_3_goMux_mux_bufchan_buf[0]))
        scfarg_0_3_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_3_1_argbuf_r) && (! scfarg_0_3_goMux_mux_bufchan_buf[0])))
        scfarg_0_3_goMux_mux_bufchan_buf <= scfarg_0_3_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) > (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aeD_3_destruct,Pointer_QTree_Int) > (t1aeD_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aeD_3_destruct_bufchan_d;
  logic t1aeD_3_destruct_bufchan_r;
  assign t1aeD_3_destruct_r = ((! t1aeD_3_destruct_bufchan_d[0]) || t1aeD_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeD_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aeD_3_destruct_r)
        t1aeD_3_destruct_bufchan_d <= t1aeD_3_destruct_d;
  Pointer_QTree_Int_t t1aeD_3_destruct_bufchan_buf;
  assign t1aeD_3_destruct_bufchan_r = (! t1aeD_3_destruct_bufchan_buf[0]);
  assign t1aeD_3_1_argbuf_d = (t1aeD_3_destruct_bufchan_buf[0] ? t1aeD_3_destruct_bufchan_buf :
                               t1aeD_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeD_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aeD_3_1_argbuf_r && t1aeD_3_destruct_bufchan_buf[0]))
        t1aeD_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aeD_3_1_argbuf_r) && (! t1aeD_3_destruct_bufchan_buf[0])))
        t1aeD_3_destruct_bufchan_buf <= t1aeD_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aeW_3_destruct,Pointer_QTree_Int) > (t1aeW_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aeW_3_destruct_bufchan_d;
  logic t1aeW_3_destruct_bufchan_r;
  assign t1aeW_3_destruct_r = ((! t1aeW_3_destruct_bufchan_d[0]) || t1aeW_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeW_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aeW_3_destruct_r)
        t1aeW_3_destruct_bufchan_d <= t1aeW_3_destruct_d;
  Pointer_QTree_Int_t t1aeW_3_destruct_bufchan_buf;
  assign t1aeW_3_destruct_bufchan_r = (! t1aeW_3_destruct_bufchan_buf[0]);
  assign t1aeW_3_1_argbuf_d = (t1aeW_3_destruct_bufchan_buf[0] ? t1aeW_3_destruct_bufchan_buf :
                               t1aeW_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aeW_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aeW_3_1_argbuf_r && t1aeW_3_destruct_bufchan_buf[0]))
        t1aeW_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aeW_3_1_argbuf_r) && (! t1aeW_3_destruct_bufchan_buf[0])))
        t1aeW_3_destruct_bufchan_buf <= t1aeW_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aed_destruct,Pointer_QTree_Int) > (t1aed_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aed_destruct_bufchan_d;
  logic t1aed_destruct_bufchan_r;
  assign t1aed_destruct_r = ((! t1aed_destruct_bufchan_d[0]) || t1aed_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aed_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aed_destruct_r) t1aed_destruct_bufchan_d <= t1aed_destruct_d;
  Pointer_QTree_Int_t t1aed_destruct_bufchan_buf;
  assign t1aed_destruct_bufchan_r = (! t1aed_destruct_bufchan_buf[0]);
  assign t1aed_1_argbuf_d = (t1aed_destruct_bufchan_buf[0] ? t1aed_destruct_bufchan_buf :
                             t1aed_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aed_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aed_1_argbuf_r && t1aed_destruct_bufchan_buf[0]))
        t1aed_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aed_1_argbuf_r) && (! t1aed_destruct_bufchan_buf[0])))
        t1aed_destruct_bufchan_buf <= t1aed_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1aes_3_destruct,Pointer_QTree_Int) > (t1aes_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1aes_3_destruct_bufchan_d;
  logic t1aes_3_destruct_bufchan_r;
  assign t1aes_3_destruct_r = ((! t1aes_3_destruct_bufchan_d[0]) || t1aes_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aes_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1aes_3_destruct_r)
        t1aes_3_destruct_bufchan_d <= t1aes_3_destruct_d;
  Pointer_QTree_Int_t t1aes_3_destruct_bufchan_buf;
  assign t1aes_3_destruct_bufchan_r = (! t1aes_3_destruct_bufchan_buf[0]);
  assign t1aes_3_1_argbuf_d = (t1aes_3_destruct_bufchan_buf[0] ? t1aes_3_destruct_bufchan_buf :
                               t1aes_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1aes_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1aes_3_1_argbuf_r && t1aes_3_destruct_bufchan_buf[0]))
        t1aes_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1aes_3_1_argbuf_r) && (! t1aes_3_destruct_bufchan_buf[0])))
        t1aes_3_destruct_bufchan_buf <= t1aes_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aeE_2_destruct,Pointer_QTree_Int) > (t2aeE_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aeE_2_destruct_bufchan_d;
  logic t2aeE_2_destruct_bufchan_r;
  assign t2aeE_2_destruct_r = ((! t2aeE_2_destruct_bufchan_d[0]) || t2aeE_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeE_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aeE_2_destruct_r)
        t2aeE_2_destruct_bufchan_d <= t2aeE_2_destruct_d;
  Pointer_QTree_Int_t t2aeE_2_destruct_bufchan_buf;
  assign t2aeE_2_destruct_bufchan_r = (! t2aeE_2_destruct_bufchan_buf[0]);
  assign t2aeE_2_1_argbuf_d = (t2aeE_2_destruct_bufchan_buf[0] ? t2aeE_2_destruct_bufchan_buf :
                               t2aeE_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeE_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aeE_2_1_argbuf_r && t2aeE_2_destruct_bufchan_buf[0]))
        t2aeE_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aeE_2_1_argbuf_r) && (! t2aeE_2_destruct_bufchan_buf[0])))
        t2aeE_2_destruct_bufchan_buf <= t2aeE_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aeX_2_destruct,Pointer_QTree_Int) > (t2aeX_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aeX_2_destruct_bufchan_d;
  logic t2aeX_2_destruct_bufchan_r;
  assign t2aeX_2_destruct_r = ((! t2aeX_2_destruct_bufchan_d[0]) || t2aeX_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeX_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aeX_2_destruct_r)
        t2aeX_2_destruct_bufchan_d <= t2aeX_2_destruct_d;
  Pointer_QTree_Int_t t2aeX_2_destruct_bufchan_buf;
  assign t2aeX_2_destruct_bufchan_r = (! t2aeX_2_destruct_bufchan_buf[0]);
  assign t2aeX_2_1_argbuf_d = (t2aeX_2_destruct_bufchan_buf[0] ? t2aeX_2_destruct_bufchan_buf :
                               t2aeX_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aeX_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aeX_2_1_argbuf_r && t2aeX_2_destruct_bufchan_buf[0]))
        t2aeX_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aeX_2_1_argbuf_r) && (! t2aeX_2_destruct_bufchan_buf[0])))
        t2aeX_2_destruct_bufchan_buf <= t2aeX_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aee_destruct,Pointer_QTree_Int) > (t2aee_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aee_destruct_bufchan_d;
  logic t2aee_destruct_bufchan_r;
  assign t2aee_destruct_r = ((! t2aee_destruct_bufchan_d[0]) || t2aee_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aee_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aee_destruct_r) t2aee_destruct_bufchan_d <= t2aee_destruct_d;
  Pointer_QTree_Int_t t2aee_destruct_bufchan_buf;
  assign t2aee_destruct_bufchan_r = (! t2aee_destruct_bufchan_buf[0]);
  assign t2aee_1_argbuf_d = (t2aee_destruct_bufchan_buf[0] ? t2aee_destruct_bufchan_buf :
                             t2aee_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aee_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aee_1_argbuf_r && t2aee_destruct_bufchan_buf[0]))
        t2aee_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aee_1_argbuf_r) && (! t2aee_destruct_bufchan_buf[0])))
        t2aee_destruct_bufchan_buf <= t2aee_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2aet_2_destruct,Pointer_QTree_Int) > (t2aet_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2aet_2_destruct_bufchan_d;
  logic t2aet_2_destruct_bufchan_r;
  assign t2aet_2_destruct_r = ((! t2aet_2_destruct_bufchan_d[0]) || t2aet_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aet_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2aet_2_destruct_r)
        t2aet_2_destruct_bufchan_d <= t2aet_2_destruct_d;
  Pointer_QTree_Int_t t2aet_2_destruct_bufchan_buf;
  assign t2aet_2_destruct_bufchan_r = (! t2aet_2_destruct_bufchan_buf[0]);
  assign t2aet_2_1_argbuf_d = (t2aet_2_destruct_bufchan_buf[0] ? t2aet_2_destruct_bufchan_buf :
                               t2aet_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2aet_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2aet_2_1_argbuf_r && t2aet_2_destruct_bufchan_buf[0]))
        t2aet_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2aet_2_1_argbuf_r) && (! t2aet_2_destruct_bufchan_buf[0])))
        t2aet_2_destruct_bufchan_buf <= t2aet_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aeF_1_destruct,Pointer_QTree_Int) > (t3aeF_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aeF_1_destruct_bufchan_d;
  logic t3aeF_1_destruct_bufchan_r;
  assign t3aeF_1_destruct_r = ((! t3aeF_1_destruct_bufchan_d[0]) || t3aeF_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeF_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aeF_1_destruct_r)
        t3aeF_1_destruct_bufchan_d <= t3aeF_1_destruct_d;
  Pointer_QTree_Int_t t3aeF_1_destruct_bufchan_buf;
  assign t3aeF_1_destruct_bufchan_r = (! t3aeF_1_destruct_bufchan_buf[0]);
  assign t3aeF_1_1_argbuf_d = (t3aeF_1_destruct_bufchan_buf[0] ? t3aeF_1_destruct_bufchan_buf :
                               t3aeF_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeF_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aeF_1_1_argbuf_r && t3aeF_1_destruct_bufchan_buf[0]))
        t3aeF_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aeF_1_1_argbuf_r) && (! t3aeF_1_destruct_bufchan_buf[0])))
        t3aeF_1_destruct_bufchan_buf <= t3aeF_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aeY_1_destruct,Pointer_QTree_Int) > (t3aeY_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aeY_1_destruct_bufchan_d;
  logic t3aeY_1_destruct_bufchan_r;
  assign t3aeY_1_destruct_r = ((! t3aeY_1_destruct_bufchan_d[0]) || t3aeY_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeY_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aeY_1_destruct_r)
        t3aeY_1_destruct_bufchan_d <= t3aeY_1_destruct_d;
  Pointer_QTree_Int_t t3aeY_1_destruct_bufchan_buf;
  assign t3aeY_1_destruct_bufchan_r = (! t3aeY_1_destruct_bufchan_buf[0]);
  assign t3aeY_1_1_argbuf_d = (t3aeY_1_destruct_bufchan_buf[0] ? t3aeY_1_destruct_bufchan_buf :
                               t3aeY_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeY_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aeY_1_1_argbuf_r && t3aeY_1_destruct_bufchan_buf[0]))
        t3aeY_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aeY_1_1_argbuf_r) && (! t3aeY_1_destruct_bufchan_buf[0])))
        t3aeY_1_destruct_bufchan_buf <= t3aeY_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aef_destruct,Pointer_QTree_Int) > (t3aef_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aef_destruct_bufchan_d;
  logic t3aef_destruct_bufchan_r;
  assign t3aef_destruct_r = ((! t3aef_destruct_bufchan_d[0]) || t3aef_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aef_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aef_destruct_r) t3aef_destruct_bufchan_d <= t3aef_destruct_d;
  Pointer_QTree_Int_t t3aef_destruct_bufchan_buf;
  assign t3aef_destruct_bufchan_r = (! t3aef_destruct_bufchan_buf[0]);
  assign t3aef_1_argbuf_d = (t3aef_destruct_bufchan_buf[0] ? t3aef_destruct_bufchan_buf :
                             t3aef_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aef_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aef_1_argbuf_r && t3aef_destruct_bufchan_buf[0]))
        t3aef_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aef_1_argbuf_r) && (! t3aef_destruct_bufchan_buf[0])))
        t3aef_destruct_bufchan_buf <= t3aef_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3aeu_1_destruct,Pointer_QTree_Int) > (t3aeu_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3aeu_1_destruct_bufchan_d;
  logic t3aeu_1_destruct_bufchan_r;
  assign t3aeu_1_destruct_r = ((! t3aeu_1_destruct_bufchan_d[0]) || t3aeu_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeu_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3aeu_1_destruct_r)
        t3aeu_1_destruct_bufchan_d <= t3aeu_1_destruct_d;
  Pointer_QTree_Int_t t3aeu_1_destruct_bufchan_buf;
  assign t3aeu_1_destruct_bufchan_r = (! t3aeu_1_destruct_bufchan_buf[0]);
  assign t3aeu_1_1_argbuf_d = (t3aeu_1_destruct_bufchan_buf[0] ? t3aeu_1_destruct_bufchan_buf :
                               t3aeu_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3aeu_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3aeu_1_1_argbuf_r && t3aeu_1_destruct_bufchan_buf[0]))
        t3aeu_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3aeu_1_1_argbuf_r) && (! t3aeu_1_destruct_bufchan_buf[0])))
        t3aeu_1_destruct_bufchan_buf <= t3aeu_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aeG_destruct,Pointer_QTree_Int) > (t4aeG_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aeG_destruct_bufchan_d;
  logic t4aeG_destruct_bufchan_r;
  assign t4aeG_destruct_r = ((! t4aeG_destruct_bufchan_d[0]) || t4aeG_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeG_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aeG_destruct_r) t4aeG_destruct_bufchan_d <= t4aeG_destruct_d;
  Pointer_QTree_Int_t t4aeG_destruct_bufchan_buf;
  assign t4aeG_destruct_bufchan_r = (! t4aeG_destruct_bufchan_buf[0]);
  assign t4aeG_1_argbuf_d = (t4aeG_destruct_bufchan_buf[0] ? t4aeG_destruct_bufchan_buf :
                             t4aeG_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeG_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aeG_1_argbuf_r && t4aeG_destruct_bufchan_buf[0]))
        t4aeG_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aeG_1_argbuf_r) && (! t4aeG_destruct_bufchan_buf[0])))
        t4aeG_destruct_bufchan_buf <= t4aeG_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aeZ_destruct,Pointer_QTree_Int) > (t4aeZ_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aeZ_destruct_bufchan_d;
  logic t4aeZ_destruct_bufchan_r;
  assign t4aeZ_destruct_r = ((! t4aeZ_destruct_bufchan_d[0]) || t4aeZ_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeZ_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aeZ_destruct_r) t4aeZ_destruct_bufchan_d <= t4aeZ_destruct_d;
  Pointer_QTree_Int_t t4aeZ_destruct_bufchan_buf;
  assign t4aeZ_destruct_bufchan_r = (! t4aeZ_destruct_bufchan_buf[0]);
  assign t4aeZ_1_argbuf_d = (t4aeZ_destruct_bufchan_buf[0] ? t4aeZ_destruct_bufchan_buf :
                             t4aeZ_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeZ_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aeZ_1_argbuf_r && t4aeZ_destruct_bufchan_buf[0]))
        t4aeZ_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aeZ_1_argbuf_r) && (! t4aeZ_destruct_bufchan_buf[0])))
        t4aeZ_destruct_bufchan_buf <= t4aeZ_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aeg_destruct,Pointer_QTree_Int) > (t4aeg_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aeg_destruct_bufchan_d;
  logic t4aeg_destruct_bufchan_r;
  assign t4aeg_destruct_r = ((! t4aeg_destruct_bufchan_d[0]) || t4aeg_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeg_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aeg_destruct_r) t4aeg_destruct_bufchan_d <= t4aeg_destruct_d;
  Pointer_QTree_Int_t t4aeg_destruct_bufchan_buf;
  assign t4aeg_destruct_bufchan_r = (! t4aeg_destruct_bufchan_buf[0]);
  assign t4aeg_1_argbuf_d = (t4aeg_destruct_bufchan_buf[0] ? t4aeg_destruct_bufchan_buf :
                             t4aeg_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aeg_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aeg_1_argbuf_r && t4aeg_destruct_bufchan_buf[0]))
        t4aeg_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aeg_1_argbuf_r) && (! t4aeg_destruct_bufchan_buf[0])))
        t4aeg_destruct_bufchan_buf <= t4aeg_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4aev_destruct,Pointer_QTree_Int) > (t4aev_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4aev_destruct_bufchan_d;
  logic t4aev_destruct_bufchan_r;
  assign t4aev_destruct_r = ((! t4aev_destruct_bufchan_d[0]) || t4aev_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aev_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4aev_destruct_r) t4aev_destruct_bufchan_d <= t4aev_destruct_d;
  Pointer_QTree_Int_t t4aev_destruct_bufchan_buf;
  assign t4aev_destruct_bufchan_r = (! t4aev_destruct_bufchan_buf[0]);
  assign t4aev_1_argbuf_d = (t4aev_destruct_bufchan_buf[0] ? t4aev_destruct_bufchan_buf :
                             t4aev_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4aev_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4aev_1_argbuf_r && t4aev_destruct_bufchan_buf[0]))
        t4aev_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4aev_1_argbuf_r) && (! t4aev_destruct_bufchan_buf[0])))
        t4aev_destruct_bufchan_buf <= t4aev_destruct_bufchan_d;
  
  /* buf (Ty Int) : (vaeM_1,Int) > (vaeM_1_argbuf,Int) */
  Int_t vaeM_1_bufchan_d;
  logic vaeM_1_bufchan_r;
  assign vaeM_1_r = ((! vaeM_1_bufchan_d[0]) || vaeM_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeM_1_bufchan_d <= {32'd0, 1'd0};
    else if (vaeM_1_r) vaeM_1_bufchan_d <= vaeM_1_d;
  Int_t vaeM_1_bufchan_buf;
  assign vaeM_1_bufchan_r = (! vaeM_1_bufchan_buf[0]);
  assign vaeM_1_argbuf_d = (vaeM_1_bufchan_buf[0] ? vaeM_1_bufchan_buf :
                            vaeM_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeM_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vaeM_1_argbuf_r && vaeM_1_bufchan_buf[0]))
        vaeM_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vaeM_1_argbuf_r) && (! vaeM_1_bufchan_buf[0])))
        vaeM_1_bufchan_buf <= vaeM_1_bufchan_d;
  
  /* fork (Ty Int) : (vaeM_destruct,Int) > [(vaeM_1,Int),(vaeM_2,Int)] */
  logic [1:0] vaeM_destruct_emitted;
  logic [1:0] vaeM_destruct_done;
  assign vaeM_1_d = {vaeM_destruct_d[32:1],
                     (vaeM_destruct_d[0] && (! vaeM_destruct_emitted[0]))};
  assign vaeM_2_d = {vaeM_destruct_d[32:1],
                     (vaeM_destruct_d[0] && (! vaeM_destruct_emitted[1]))};
  assign vaeM_destruct_done = (vaeM_destruct_emitted | ({vaeM_2_d[0],
                                                         vaeM_1_d[0]} & {vaeM_2_r, vaeM_1_r}));
  assign vaeM_destruct_r = (& vaeM_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaeM_destruct_emitted <= 2'd0;
    else
      vaeM_destruct_emitted <= (vaeM_destruct_r ? 2'd0 :
                                vaeM_destruct_done);
  
  /* buf (Ty Int) : (vaei_destruct,Int) > (vaei_1_argbuf,Int) */
  Int_t vaei_destruct_bufchan_d;
  logic vaei_destruct_bufchan_r;
  assign vaei_destruct_r = ((! vaei_destruct_bufchan_d[0]) || vaei_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaei_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vaei_destruct_r) vaei_destruct_bufchan_d <= vaei_destruct_d;
  Int_t vaei_destruct_bufchan_buf;
  assign vaei_destruct_bufchan_r = (! vaei_destruct_bufchan_buf[0]);
  assign vaei_1_argbuf_d = (vaei_destruct_bufchan_buf[0] ? vaei_destruct_bufchan_buf :
                            vaei_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vaei_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vaei_1_argbuf_r && vaei_destruct_bufchan_buf[0]))
        vaei_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vaei_1_argbuf_r) && (! vaei_destruct_bufchan_buf[0])))
        vaei_destruct_bufchan_buf <= vaei_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (lizzieLet30_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet47_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet47_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet47_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet47_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca2_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet47_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet48_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet48_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet48_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet48_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet48_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet49_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet49_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet49_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet49_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet49_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca3_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > (writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf  :
                                                                         \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) > (sca3_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet11_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > (writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf  :
                                                                         \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) > (lizzieLet4_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet4_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet43_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > (writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf  :
                                                                         \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) > (sca2_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet51_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > (writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf  :
                                                                         \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) > (sca1_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet52_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) > (writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_d  = (\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf  :
                                                                         \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_r  && \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_r ) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'''''''''_f'''''''''_Int) : (writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb,Pointer_CTf'''''''''_f'''''''''_Int) > (sca0_1_1_argbuf,Pointer_CTf'''''''''_f'''''''''_Int) */
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_r  = ((! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_r )
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_d ;
  \Pointer_CTf'''''''''_f'''''''''_Int_t  \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_r  = (! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_buf  <= \writeCTf'''''''''_f'''''''''_IntlizzieLet53_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet21_1_argbuf,Pointer_CTf'_f'_Int) > (writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_r  = ((! \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet21_1_argbuf_r )
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d  <= \writeCTf'_f'_IntlizzieLet21_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_d  = (\writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf  :
                                                         \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_r  && \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_r ) && (! \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet21_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb,Pointer_CTf'_f'_Int) > (sca3_2_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_r  = ((! \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_r )
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet21_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet44_1_argbuf,Pointer_CTf'_f'_Int) > (writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_r  = ((! \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet44_1_argbuf_r )
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d  <= \writeCTf'_f'_IntlizzieLet44_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_d  = (\writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf  :
                                                         \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_r  && \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_r ) && (! \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet44_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb,Pointer_CTf'_f'_Int) > (lizzieLet12_1_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_r  = ((! \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_r )
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet12_1_1_argbuf_d = (\writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf  :
                                     \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet44_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet56_1_argbuf,Pointer_CTf'_f'_Int) > (writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_r  = ((! \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet56_1_argbuf_r )
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d  <= \writeCTf'_f'_IntlizzieLet56_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_d  = (\writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf  :
                                                         \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_r  && \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_r ) && (! \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet56_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb,Pointer_CTf'_f'_Int) > (sca2_2_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_r  = ((! \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_r )
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet56_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet57_1_argbuf,Pointer_CTf'_f'_Int) > (writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_r  = ((! \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet57_1_argbuf_r )
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d  <= \writeCTf'_f'_IntlizzieLet57_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_d  = (\writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf  :
                                                         \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_r  && \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_r ) && (! \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet57_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb,Pointer_CTf'_f'_Int) > (sca1_2_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_r  = ((! \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_r )
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet57_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet58_1_argbuf,Pointer_CTf'_f'_Int) > (writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_r  = ((! \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet58_1_argbuf_r )
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d  <= \writeCTf'_f'_IntlizzieLet58_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_d  = (\writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf  :
                                                         \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_r  && \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_r ) && (! \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet58_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int) : (writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb,Pointer_CTf'_f'_Int) > (sca0_2_1_argbuf,Pointer_CTf'_f'_Int) */
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_r  = ((! \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                               1'd0};
    else
      if (\writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_r )
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_t  \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                 1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                   1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_IntlizzieLet58_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet40_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet40_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet40_1_argbuf_r = ((! writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet40_1_argbuf_r)
        writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet40_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet40_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet40_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet40_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet40_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet40_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca3_3_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet40_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet40_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet40_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_3_1_argbuf_d = (writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca3_3_1_argbuf_r && writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca3_3_1_argbuf_r) && (! writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet40_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet45_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet45_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet45_1_argbuf_r = ((! writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet45_1_argbuf_r)
        writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet45_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet45_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet45_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet45_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet45_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet45_1_argbuf_rwb,Pointer_CTf_f_Int) > (lizzieLet27_1_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet45_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet45_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet45_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet27_1_1_argbuf_d = (writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf :
                                     writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet27_1_1_argbuf_r && writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet27_1_1_argbuf_r) && (! writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet45_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet61_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet61_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet61_1_argbuf_r = ((! writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet61_1_argbuf_r)
        writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet61_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet61_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet61_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet61_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet61_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet61_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca2_3_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet61_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet61_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet61_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_3_1_argbuf_d = (writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca2_3_1_argbuf_r && writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca2_3_1_argbuf_r) && (! writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet61_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet62_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet62_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet62_1_argbuf_r = ((! writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet62_1_argbuf_r)
        writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet62_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet62_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet62_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet62_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet62_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet62_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca1_3_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet62_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet62_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet62_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_3_1_argbuf_d = (writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca1_3_1_argbuf_r && writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca1_3_1_argbuf_r) && (! writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet62_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet63_1_argbuf,Pointer_CTf_f_Int) > (writeCTf_f_IntlizzieLet63_1_argbuf_rwb,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d;
  logic writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_r;
  assign writeCTf_f_IntlizzieLet63_1_argbuf_r = ((! writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d[0]) || writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet63_1_argbuf_r)
        writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d <= writeCTf_f_IntlizzieLet63_1_argbuf_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf;
  assign writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_r = (! writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_IntlizzieLet63_1_argbuf_rwb_d = (writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf[0] ? writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf :
                                                     writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCTf_f_IntlizzieLet63_1_argbuf_rwb_r && writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCTf_f_IntlizzieLet63_1_argbuf_rwb_r) && (! writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_buf <= writeCTf_f_IntlizzieLet63_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int) : (writeCTf_f_IntlizzieLet63_1_argbuf_rwb,Pointer_CTf_f_Int) > (sca0_3_1_argbuf,Pointer_CTf_f_Int) */
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_IntlizzieLet63_1_argbuf_rwb_r = ((! writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCTf_f_IntlizzieLet63_1_argbuf_rwb_r)
        writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d <= writeCTf_f_IntlizzieLet63_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_t writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_r = (! writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_3_1_argbuf_d = (writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((sca0_3_1_argbuf_r && writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! sca0_3_1_argbuf_r) && (! writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_buf <= writeCTf_f_IntlizzieLet63_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_r = ((! writeQTree_IntlizzieLet10_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_r)
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_d = (writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet10_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet10_1_argbuf_rwb_r && writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet10_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet12_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_argbuf_r = ((! writeQTree_IntlizzieLet12_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_argbuf_r)
        writeQTree_IntlizzieLet12_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet12_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet12_1_argbuf_rwb_d = (writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet12_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet12_1_argbuf_rwb_r && writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet12_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet12_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet12_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet12_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_r = ((! writeQTree_IntlizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_r)
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_d = (writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet15_1_argbuf_rwb_r && writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet15_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet15_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet15_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_r = ((! writeQTree_IntlizzieLet16_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_r)
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_d = (writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet16_1_argbuf_rwb_r && writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet16_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_r = ((! writeQTree_IntlizzieLet17_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_r)
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_d = (writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet17_1_argbuf_rwb_r && writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet17_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet17_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet17_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet17_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_r = ((! writeQTree_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_r)
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_d = (writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet18_1_argbuf_rwb_r && writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet18_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet18_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet18_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_r = ((! writeQTree_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_r)
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_d = (writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet20_1_argbuf_rwb_r && writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet20_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet20_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet20_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_r = ((! writeQTree_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_r)
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_d = (writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet22_1_argbuf_rwb_r && writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet22_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet22_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet22_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet23_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet23_1_argbuf_r = ((! writeQTree_IntlizzieLet23_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet23_1_argbuf_r)
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet23_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet23_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_d = (writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet23_1_argbuf_rwb_r && writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet23_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet23_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet23_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet23_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet25_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_argbuf_r = ((! writeQTree_IntlizzieLet25_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_argbuf_r)
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet25_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_d = (writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet25_1_argbuf_rwb_r && writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet25_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet25_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet25_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet25_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_2_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet28_2_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet28_2_1_argbuf_r = ((! writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_2_1_argbuf_r)
        writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet28_2_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet28_2_1_argbuf_rwb_d = (writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet28_2_1_argbuf_rwb_r && writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet28_2_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet28_2_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_2_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet15_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet28_2_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet28_2_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet28_2_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet15_1_1_argbuf_d = (writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet15_1_1_argbuf_r && writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet15_1_1_argbuf_r) && (! writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet28_2_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet29_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet29_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet29_1_1_argbuf_r = ((! writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet29_1_1_argbuf_r)
        writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet29_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet29_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet29_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet29_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet29_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet29_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet16_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet29_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet29_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet29_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet16_1_1_argbuf_d = (writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet16_1_1_argbuf_r && writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet16_1_1_argbuf_r) && (! writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet29_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet30_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet30_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet30_1_1_argbuf_r = ((! writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet30_1_1_argbuf_r)
        writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet30_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet30_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet30_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet30_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet30_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet30_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet17_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet30_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet30_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet30_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet17_1_1_argbuf_d = (writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet17_1_1_argbuf_r && writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet17_1_1_argbuf_r) && (! writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet30_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_r = ((! writeQTree_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_r)
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_d = (writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet31_1_argbuf_rwb_r && writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet31_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet31_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet18_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet31_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet18_1_1_argbuf_d = (writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet18_1_1_argbuf_r && writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet18_1_1_argbuf_r) && (! writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet33_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_1_argbuf_r = ((! writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_1_argbuf_r)
        writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet33_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet33_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet33_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet33_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet33_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet19_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet33_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_1_argbuf_d = (writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet19_1_1_argbuf_r && writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet19_1_1_argbuf_r) && (! writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet33_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_r = ((! writeQTree_IntlizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_r)
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_d = (writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet33_1_argbuf_rwb_r && writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet33_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet33_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet19_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet33_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_r = ((! writeQTree_IntlizzieLet34_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_r)
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_d = (writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet34_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet34_1_argbuf_rwb_r && writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet34_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet34_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet20_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet34_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet34_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet20_1_1_argbuf_d = (writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet20_1_1_argbuf_r && writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet20_1_1_argbuf_r) && (! writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet34_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet35_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet35_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet35_1_argbuf_r = ((! writeQTree_IntlizzieLet35_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet35_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet35_1_argbuf_r)
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet35_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet35_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_d = (writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet35_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet35_1_argbuf_rwb_r && writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet35_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet35_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet35_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet35_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet21_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet35_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet35_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet21_1_1_argbuf_d = (writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet21_1_1_argbuf_r && writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet21_1_1_argbuf_r) && (! writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet35_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet36_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet36_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet36_1_argbuf_r = ((! writeQTree_IntlizzieLet36_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet36_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet36_1_argbuf_r)
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet36_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet36_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_d = (writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet36_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet36_1_argbuf_rwb_r && writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet36_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet36_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet36_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet36_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet22_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet36_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet36_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet22_1_1_argbuf_d = (writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet22_1_1_argbuf_r && writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet22_1_1_argbuf_r) && (! writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet36_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet38_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_argbuf_r = ((! writeQTree_IntlizzieLet38_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_argbuf_r)
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet38_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_d = (writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet38_1_argbuf_rwb_r && writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet38_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet38_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet23_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet38_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet38_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet23_1_1_argbuf_d = (writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet23_1_1_argbuf_r && writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet23_1_1_argbuf_r) && (! writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet39_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_argbuf_r = ((! writeQTree_IntlizzieLet39_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_argbuf_r)
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet39_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_d = (writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet39_1_argbuf_rwb_r && writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet39_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet39_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet39_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet24_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet39_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet39_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet24_1_1_argbuf_d = (writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet24_1_1_argbuf_r && writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet24_1_1_argbuf_r) && (! writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet39_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet41_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet41_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet41_1_argbuf_r = ((! writeQTree_IntlizzieLet41_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet41_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet41_1_argbuf_r)
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet41_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet41_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_d = (writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet41_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet41_1_argbuf_rwb_r && writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet41_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet41_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet41_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet41_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet25_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet41_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet41_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet25_1_1_argbuf_d = (writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet25_1_1_argbuf_r && writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet25_1_1_argbuf_r) && (! writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet41_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet42_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet42_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet42_1_argbuf_r = ((! writeQTree_IntlizzieLet42_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet42_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet42_1_argbuf_r)
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet42_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet42_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_d = (writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet42_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet42_1_argbuf_rwb_r && writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet42_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet42_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet42_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet42_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet26_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet42_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet42_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet26_1_1_argbuf_d = (writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet26_1_1_argbuf_r && writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet26_1_1_argbuf_r) && (! writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet42_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet54_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet54_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet54_1_argbuf_r = ((! writeQTree_IntlizzieLet54_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet54_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet54_1_argbuf_r)
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet54_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet54_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_d = (writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet54_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet54_1_argbuf_rwb_r && writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet54_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet54_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet54_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet54_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet54_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet54_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet54_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet59_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet59_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet59_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet59_1_argbuf_r = ((! writeQTree_IntlizzieLet59_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet59_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet59_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet59_1_argbuf_r)
        writeQTree_IntlizzieLet59_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet59_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet59_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet59_1_argbuf_rwb_d = (writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet59_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet59_1_argbuf_rwb_r && writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet59_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet59_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet59_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet59_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet59_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet59_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet59_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet59_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet64_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet64_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet64_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet64_1_argbuf_r = ((! writeQTree_IntlizzieLet64_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet64_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet64_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet64_1_argbuf_r)
        writeQTree_IntlizzieLet64_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet64_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet64_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet64_1_argbuf_rwb_d = (writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet64_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet64_1_argbuf_rwb_r && writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet64_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet64_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet64_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet64_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet64_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet64_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet64_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_3_1_argbuf_d = (writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_3_1_argbuf_r && writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_3_1_argbuf_r) && (! writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet64_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wsjQ_1_goMux_mux,Pointer_QTree_Int) > (wsjQ_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wsjQ_1_goMux_mux_bufchan_d;
  logic wsjQ_1_goMux_mux_bufchan_r;
  assign wsjQ_1_goMux_mux_r = ((! wsjQ_1_goMux_mux_bufchan_d[0]) || wsjQ_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsjQ_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wsjQ_1_goMux_mux_r)
        wsjQ_1_goMux_mux_bufchan_d <= wsjQ_1_goMux_mux_d;
  Pointer_QTree_Int_t wsjQ_1_goMux_mux_bufchan_buf;
  assign wsjQ_1_goMux_mux_bufchan_r = (! wsjQ_1_goMux_mux_bufchan_buf[0]);
  assign wsjQ_1_1_argbuf_d = (wsjQ_1_goMux_mux_bufchan_buf[0] ? wsjQ_1_goMux_mux_bufchan_buf :
                              wsjQ_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsjQ_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wsjQ_1_1_argbuf_r && wsjQ_1_goMux_mux_bufchan_buf[0]))
        wsjQ_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wsjQ_1_1_argbuf_r) && (! wsjQ_1_goMux_mux_bufchan_buf[0])))
        wsjQ_1_goMux_mux_bufchan_buf <= wsjQ_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) > (lizzieLet48_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d;
  logic wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_r;
  assign wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_r = ((! wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d[0]) || wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_r)
        wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d <= wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_d;
  CT$wnnz_Int_t wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf;
  assign wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_r = (! wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet48_1_argbuf_d = (wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf[0] ? wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf :
                                   wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet48_1_argbuf_r && wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf[0]))
        wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet48_1_argbuf_r) && (! wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf[0])))
        wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_buf <= wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int1) : [(wwsjT_2_destruct,Int#),
                                (lizzieLet46_4Lcall_$wnnz_Int2,Int#),
                                (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                (q4a88_2_destruct,Pointer_QTree_Int)] > (wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) */
  assign wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_d = Lcall_$wnnz_Int1_dc((& {wwsjT_2_destruct_d[0],
                                                                                                               lizzieLet46_4Lcall_$wnnz_Int2_d[0],
                                                                                                               sc_0_5_destruct_d[0],
                                                                                                               q4a88_2_destruct_d[0]}), wwsjT_2_destruct_d, lizzieLet46_4Lcall_$wnnz_Int2_d, sc_0_5_destruct_d, q4a88_2_destruct_d);
  assign {wwsjT_2_destruct_r,
          lizzieLet46_4Lcall_$wnnz_Int2_r,
          sc_0_5_destruct_r,
          q4a88_2_destruct_r} = {4 {(wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_r && wwsjT_2_1lizzieLet46_4Lcall_$wnnz_Int2_1sc_0_5_1q4a88_2_1Lcall_$wnnz_Int1_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) > (lizzieLet49_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  logic wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r;
  assign wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r = ((! wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d[0]) || wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= {115'd0,
                                                                                               1'd0};
    else
      if (wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r)
        wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d <= wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d;
  CT$wnnz_Int_t wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf;
  assign wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_r = (! wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet49_1_argbuf_d = (wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0] ? wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf :
                                   wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet49_1_argbuf_r && wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0]))
        wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet49_1_argbuf_r) && (! wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf[0])))
        wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_buf <= wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int0) : [(wwsjT_3_destruct,Int#),
                                (ww1Xkr_1_destruct,Int#),
                                (lizzieLet46_4Lcall_$wnnz_Int1,Int#),
                                (sc_0_6_destruct,Pointer_CT$wnnz_Int)] > (wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0,CT$wnnz_Int) */
  assign wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d = Lcall_$wnnz_Int0_dc((& {wwsjT_3_destruct_d[0],
                                                                                                                ww1Xkr_1_destruct_d[0],
                                                                                                                lizzieLet46_4Lcall_$wnnz_Int1_d[0],
                                                                                                                sc_0_6_destruct_d[0]}), wwsjT_3_destruct_d, ww1Xkr_1_destruct_d, lizzieLet46_4Lcall_$wnnz_Int1_d, sc_0_6_destruct_d);
  assign {wwsjT_3_destruct_r,
          ww1Xkr_1_destruct_r,
          lizzieLet46_4Lcall_$wnnz_Int1_r,
          sc_0_6_destruct_r} = {4 {(wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_r && wwsjT_3_1ww1Xkr_1_1lizzieLet46_4Lcall_$wnnz_Int1_1sc_0_6_1Lcall_$wnnz_Int0_d[0])}};
  
  /* op_add (Ty Int#) : (wwsjT_4_1ww1Xkr_2_1_Add32,Int#) (ww2Xku_1_destruct,Int#) > (es_6_2_1ww2Xku_1_1_Add32,Int#) */
  assign es_6_2_1ww2Xku_1_1_Add32_d = {(wwsjT_4_1ww1Xkr_2_1_Add32_d[32:1] + ww2Xku_1_destruct_d[32:1]),
                                       (wwsjT_4_1ww1Xkr_2_1_Add32_d[0] && ww2Xku_1_destruct_d[0])};
  assign {wwsjT_4_1ww1Xkr_2_1_Add32_r,
          ww2Xku_1_destruct_r} = {2 {(es_6_2_1ww2Xku_1_1_Add32_r && es_6_2_1ww2Xku_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwsjT_4_destruct,Int#) (ww1Xkr_2_destruct,Int#) > (wwsjT_4_1ww1Xkr_2_1_Add32,Int#) */
  assign wwsjT_4_1ww1Xkr_2_1_Add32_d = {(wwsjT_4_destruct_d[32:1] + ww1Xkr_2_destruct_d[32:1]),
                                        (wwsjT_4_destruct_d[0] && ww1Xkr_2_destruct_d[0])};
  assign {wwsjT_4_destruct_r,
          ww1Xkr_2_destruct_r} = {2 {(wwsjT_4_1ww1Xkr_2_1_Add32_r && wwsjT_4_1ww1Xkr_2_1_Add32_d[0])}};
endmodule