`timescale 1ns/1ns
import mMapAdd_package::*;

module mMapAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t w1sm4_1_1_d,
  output logic w1sm4_1_1_r,
  input Pointer_QTree_Int_t wsm3_1_0_d,
  output logic wsm3_1_0_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_0_1I#_dout ,
  input logic \es_0_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (w1sm4_1_1, 16, 65536, Pointer_QTree_Int), (wsm3_1_0, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_0_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wmAdd_Int 16 3 (0,[0]) (1,[16p,0,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,0,16p,16p,16p,16p]) (3,[16p,16p,16p,0,16p,16p]) (4,[16p,16p,16p,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CT__024wnnz 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTmain_map__027_Int_Bool 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p]) (3,[16p,16p,16p,0,0,16p]) (4,[16p,16p,16p,16p])
TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,0,16p,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Bool 16 0 (0,[0,16p])
TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT__024wmAdd_Int 16 0 (0,[0,0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_CT__024wnnz 16 0 (0,[0,16p,16p])
TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map__027_Int_Bool 16 0 (0,[0,0,0,16p,16p])
TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int 16 0 (0,[0,0,0,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t goFork_d;
  logic goFork_r;
  Go_t goFor_2_d;
  logic goFor_2_r;
  Go_t goFor_3_d;
  logic goFor_3_r;
  Go_t goFor_4_d;
  logic goFor_4_r;
  Go_t goFor_5_d;
  logic goFor_5_r;
  Go_t goFor_6_d;
  logic goFor_6_r;
  Go_t goFor_7_d;
  logic goFor_7_r;
  Go_t goFor_8_d;
  logic goFor_8_r;
  Go_t goFor_9_d;
  logic goFor_9_r;
  \Word16#_t  initHP_CT$wmAdd_Int_d;
  logic initHP_CT$wmAdd_Int_r;
  \Word16#_t  incrHP_CT$wmAdd_Int_d;
  logic incrHP_CT$wmAdd_Int_r;
  Go_t incrHP_mergeCT$wmAdd_Int_d;
  logic incrHP_mergeCT$wmAdd_Int_r;
  Go_t incrHP_CT$wmAdd_Int1_d;
  logic incrHP_CT$wmAdd_Int1_r;
  Go_t incrHP_CT$wmAdd_Int2_d;
  logic incrHP_CT$wmAdd_Int2_r;
  \Word16#_t  addHP_CT$wmAdd_Int_d;
  logic addHP_CT$wmAdd_Int_r;
  \Word16#_t  mergeHP_CT$wmAdd_Int_d;
  logic mergeHP_CT$wmAdd_Int_r;
  Go_t incrHP_mergeCT$wmAdd_Int_buf_d;
  logic incrHP_mergeCT$wmAdd_Int_buf_r;
  \Word16#_t  mergeHP_CT$wmAdd_Int_buf_d;
  logic mergeHP_CT$wmAdd_Int_buf_r;
  \Word16#_t  forkHP1_CT$wmAdd_Int_d;
  logic forkHP1_CT$wmAdd_Int_r;
  \Word16#_t  forkHP1_CT$wmAdd_In2_d;
  logic forkHP1_CT$wmAdd_In2_r;
  \Word16#_t  forkHP1_CT$wmAdd_In3_d;
  logic forkHP1_CT$wmAdd_In3_r;
  C2_t memMergeChoice_CT$wmAdd_Int_d;
  logic memMergeChoice_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_d;
  logic memMergeIn_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_d;
  logic memOut_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memReadOut_CT$wmAdd_Int_d;
  logic memReadOut_CT$wmAdd_Int_r;
  MemOut_CT$wmAdd_Int_t memWriteOut_CT$wmAdd_Int_d;
  logic memWriteOut_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_dbuf_d;
  logic memMergeIn_CT$wmAdd_Int_dbuf_r;
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_rbuf_d;
  logic memMergeIn_CT$wmAdd_Int_rbuf_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_dbuf_d;
  logic memOut_CT$wmAdd_Int_dbuf_r;
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_rbuf_d;
  logic memOut_CT$wmAdd_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wmAdd_Int_d;
  logic destructReadIn_CT$wmAdd_Int_r;
  MemIn_CT$wmAdd_Int_t dconReadIn_CT$wmAdd_Int_d;
  logic dconReadIn_CT$wmAdd_Int_r;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wmAdd_Int_d;
  logic writeMerge_choice_CT$wmAdd_Int_r;
  CT$wmAdd_Int_t writeMerge_data_CT$wmAdd_Int_d;
  logic writeMerge_data_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet12_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet26_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_d;
  logic writeCT$wmAdd_IntlizzieLet27_1_argbuf_r;
  MemIn_CT$wmAdd_Int_t dconWriteIn_CT$wmAdd_Int_d;
  logic dconWriteIn_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t dconPtr_CT$wmAdd_Int_d;
  logic dconPtr_CT$wmAdd_Int_r;
  Pointer_CT$wmAdd_Int_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  Pointer_CT$wmAdd_Int_t demuxWriteResult_CT$wmAdd_Int_d;
  logic demuxWriteResult_CT$wmAdd_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C3_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intma8M_1_argbuf_d;
  logic readPointer_QTree_Intma8M_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intw1slS_1_1_argbuf_d;
  logic readPointer_QTree_Intw1slS_1_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intw2slT_1_1_argbuf_d;
  logic readPointer_QTree_Intw2slT_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C8_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet14_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  initHP_CT$wnnz_d;
  logic initHP_CT$wnnz_r;
  \Word16#_t  incrHP_CT$wnnz_d;
  logic incrHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_d;
  logic incrHP_mergeCT$wnnz_r;
  Go_t incrHP_CT$wnnz1_d;
  logic incrHP_CT$wnnz1_r;
  Go_t incrHP_CT$wnnz2_d;
  logic incrHP_CT$wnnz2_r;
  \Word16#_t  addHP_CT$wnnz_d;
  logic addHP_CT$wnnz_r;
  \Word16#_t  mergeHP_CT$wnnz_d;
  logic mergeHP_CT$wnnz_r;
  Go_t incrHP_mergeCT$wnnz_buf_d;
  logic incrHP_mergeCT$wnnz_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_buf_d;
  logic mergeHP_CT$wnnz_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_d;
  logic forkHP1_CT$wnnz_r;
  \Word16#_t  forkHP1_CT$wnn2_d;
  logic forkHP1_CT$wnn2_r;
  \Word16#_t  forkHP1_CT$wnn3_d;
  logic forkHP1_CT$wnn3_r;
  C2_t memMergeChoice_CT$wnnz_d;
  logic memMergeChoice_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_d;
  logic memMergeIn_CT$wnnz_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_d;
  logic memOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memReadOut_CT$wnnz_d;
  logic memReadOut_CT$wnnz_r;
  MemOut_CT$wnnz_t memWriteOut_CT$wnnz_d;
  logic memWriteOut_CT$wnnz_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_dbuf_d;
  logic memMergeIn_CT$wnnz_dbuf_r;
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_rbuf_d;
  logic memMergeIn_CT$wnnz_rbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_dbuf_d;
  logic memOut_CT$wnnz_dbuf_r;
  MemOut_CT$wnnz_t memOut_CT$wnnz_rbuf_d;
  logic memOut_CT$wnnz_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_d;
  logic destructReadIn_CT$wnnz_r;
  MemIn_CT$wnnz_t dconReadIn_CT$wnnz_d;
  logic dconReadIn_CT$wnnz_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_1_argbuf_d;
  logic readPointer_CT$wnnzscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_d;
  logic writeMerge_choice_CT$wnnz_r;
  CT$wnnz_t writeMerge_data_CT$wnnz_d;
  logic writeMerge_data_CT$wnnz_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_d;
  logic writeCT$wnnzlizzieLet16_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_d;
  logic writeCT$wnnzlizzieLet1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_d;
  logic writeCT$wnnzlizzieLet30_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_d;
  logic writeCT$wnnzlizzieLet31_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_d;
  logic writeCT$wnnzlizzieLet32_1_argbuf_r;
  MemIn_CT$wnnz_t dconWriteIn_CT$wnnz_d;
  logic dconWriteIn_CT$wnnz_r;
  Pointer_CT$wnnz_t dconPtr_CT$wnnz_d;
  logic dconPtr_CT$wnnz_r;
  Pointer_CT$wnnz_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Pointer_CT$wnnz_t demuxWriteResult_CT$wnnz_d;
  logic demuxWriteResult_CT$wnnz_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Boo2_d;
  logic forkHP1_QTree_Boo2_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_BoolwslW_1_1_argbuf_d;
  logic readPointer_QTree_BoolwslW_1_1_argbuf_r;
  C5_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_d;
  logic writeQTree_BoollizzieLet20_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_d;
  logic writeQTree_BoollizzieLet22_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  \initHP_CTmain_map'_Int_Bool_d ;
  logic \initHP_CTmain_map'_Int_Bool_r ;
  \Word16#_t  \incrHP_CTmain_map'_Int_Bool_d ;
  logic \incrHP_CTmain_map'_Int_Bool_r ;
  Go_t \incrHP_mergeCTmain_map'_Int_Bool_d ;
  logic \incrHP_mergeCTmain_map'_Int_Bool_r ;
  Go_t \incrHP_CTmain_map'_Int_Bool1_d ;
  logic \incrHP_CTmain_map'_Int_Bool1_r ;
  Go_t \incrHP_CTmain_map'_Int_Bool2_d ;
  logic \incrHP_CTmain_map'_Int_Bool2_r ;
  \Word16#_t  \addHP_CTmain_map'_Int_Bool_d ;
  logic \addHP_CTmain_map'_Int_Bool_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Bool_d ;
  logic \mergeHP_CTmain_map'_Int_Bool_r ;
  Go_t \incrHP_mergeCTmain_map'_Int_Bool_buf_d ;
  logic \incrHP_mergeCTmain_map'_Int_Bool_buf_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Bool_buf_d ;
  logic \mergeHP_CTmain_map'_Int_Bool_buf_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_Bool_d ;
  logic \forkHP1_CTmain_map'_Int_Bool_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_Boo2_d ;
  logic \forkHP1_CTmain_map'_Int_Boo2_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Int_Boo3_d ;
  logic \forkHP1_CTmain_map'_Int_Boo3_r ;
  C2_t \memMergeChoice_CTmain_map'_Int_Bool_d ;
  logic \memMergeChoice_CTmain_map'_Int_Bool_r ;
  \MemIn_CTmain_map'_Int_Bool_t  \memMergeIn_CTmain_map'_Int_Bool_d ;
  logic \memMergeIn_CTmain_map'_Int_Bool_r ;
  \MemOut_CTmain_map'_Int_Bool_t  \memOut_CTmain_map'_Int_Bool_d ;
  logic \memOut_CTmain_map'_Int_Bool_r ;
  \MemOut_CTmain_map'_Int_Bool_t  \memReadOut_CTmain_map'_Int_Bool_d ;
  logic \memReadOut_CTmain_map'_Int_Bool_r ;
  \MemOut_CTmain_map'_Int_Bool_t  \memWriteOut_CTmain_map'_Int_Bool_d ;
  logic \memWriteOut_CTmain_map'_Int_Bool_r ;
  \MemIn_CTmain_map'_Int_Bool_t  \memMergeIn_CTmain_map'_Int_Bool_dbuf_d ;
  logic \memMergeIn_CTmain_map'_Int_Bool_dbuf_r ;
  \MemIn_CTmain_map'_Int_Bool_t  \memMergeIn_CTmain_map'_Int_Bool_rbuf_d ;
  logic \memMergeIn_CTmain_map'_Int_Bool_rbuf_r ;
  \MemOut_CTmain_map'_Int_Bool_t  \memOut_CTmain_map'_Int_Bool_dbuf_d ;
  logic \memOut_CTmain_map'_Int_Bool_dbuf_r ;
  \MemOut_CTmain_map'_Int_Bool_t  \memOut_CTmain_map'_Int_Bool_rbuf_d ;
  logic \memOut_CTmain_map'_Int_Bool_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmain_map'_Int_Bool_d ;
  logic \destructReadIn_CTmain_map'_Int_Bool_r ;
  \MemIn_CTmain_map'_Int_Bool_t  \dconReadIn_CTmain_map'_Int_Bool_d ;
  logic \dconReadIn_CTmain_map'_Int_Bool_r ;
  \CTmain_map'_Int_Bool_t  \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmain_map'_Int_Bool_d ;
  logic \writeMerge_choice_CTmain_map'_Int_Bool_r ;
  \CTmain_map'_Int_Bool_t  \writeMerge_data_CTmain_map'_Int_Bool_d ;
  logic \writeMerge_data_CTmain_map'_Int_Bool_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_r ;
  \MemIn_CTmain_map'_Int_Bool_t  \dconWriteIn_CTmain_map'_Int_Bool_d ;
  logic \dconWriteIn_CTmain_map'_Int_Bool_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \dconPtr_CTmain_map'_Int_Bool_d ;
  logic \dconPtr_CTmain_map'_Int_Bool_r ;
  \Pointer_CTmain_map'_Int_Bool_t  _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  \Pointer_CTmain_map'_Int_Bool_t  \demuxWriteResult_CTmain_map'_Int_Bool_d ;
  logic \demuxWriteResult_CTmain_map'_Int_Bool_r ;
  Go_t go_1_argbuf_d;
  logic go_1_argbuf_r;
  Go_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_r ;
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_r ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_r ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_r ;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Int_t w1slS_1_argbuf_d;
  logic w1slS_1_argbuf_r;
  Pointer_QTree_Int_t w2slT_1_argbuf_d;
  logic w2slT_1_argbuf_r;
  MyDTInt_Int_Int_t wslR_1_argbuf_d;
  logic wslR_1_argbuf_r;
  Pointer_QTree_Int_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_r ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_r ;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  Go_t go_7_3_d;
  logic go_7_3_r;
  Go_t go_7_4_d;
  logic go_7_4_r;
  Go_t go_7_5_d;
  logic go_7_5_r;
  Go_t go_7_6_d;
  logic go_7_6_r;
  Pointer_QTree_Int_t w1sm4_1_argbuf_d;
  logic w1sm4_1_argbuf_r;
  Pointer_QTree_Int_t wsm3_1_argbuf_d;
  logic wsm3_1_argbuf_r;
  Int_t \es_0_1I#_d ;
  logic \es_0_1I#_r ;
  Go_t \$wnnzTupGo___Pointer_QTree_Boolgo_8_d ;
  logic \$wnnzTupGo___Pointer_QTree_Boolgo_8_r ;
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwslW_d ;
  logic \$wnnzTupGo___Pointer_QTree_BoolwslW_r ;
  Go_t go_8_1_d;
  logic go_8_1_r;
  Go_t go_8_2_d;
  logic go_8_2_r;
  Pointer_QTree_Bool_t wslW_1_argbuf_d;
  logic wslW_1_argbuf_r;
  \Int#_t  \$wmain_resbuf_d ;
  logic \$wmain_resbuf_r ;
  Go_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_r;
  MyDTBool_Bool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r;
  MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r;
  MyDTBool_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTBool_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTBool_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t es_0_4_1_d;
  logic es_0_4_1_r;
  MyBool_t es_0_4_2_d;
  logic es_0_4_2_r;
  MyBool_t es_0_4_3_d;
  logic es_0_4_3_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_r;
  MyDTInt_Bool_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Bool_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Bool_t arg0_2_3_d;
  logic arg0_2_3_r;
  MyBool_t xa88_1_d;
  logic xa88_1_r;
  MyBool_t xa88_2_d;
  logic xa88_2_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r;
  MyDTInt_Int_Int_t arg0_4_1_d;
  logic arg0_4_1_r;
  MyDTInt_Int_Int_t arg0_4_2_d;
  logic arg0_4_2_r;
  MyDTInt_Int_Int_t arg0_4_3_d;
  logic arg0_4_3_r;
  QTree_Int_t es_0_3_1QVal_Int_d;
  logic es_0_3_1QVal_Int_r;
  MyBool_t arg0_1Dcon_main2_d;
  logic arg0_1Dcon_main2_r;
  MyBool_t arg0_1Dcon_main2_1_d;
  logic arg0_1Dcon_main2_1_r;
  MyBool_t arg0_1Dcon_main2_2_d;
  logic arg0_1Dcon_main2_2_r;
  Go_t arg0_1Dcon_main2_1MyFalse_d;
  logic arg0_1Dcon_main2_1MyFalse_r;
  Go_t arg0_1Dcon_main2_1MyTrue_d;
  logic arg0_1Dcon_main2_1MyTrue_r;
  MyBool_t arg0_1Dcon_main2_1MyFalse_1MyTrue_d;
  logic arg0_1Dcon_main2_1MyFalse_1MyTrue_r;
  MyBool_t applyfnBool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_5_resbuf_r;
  MyBool_t arg0_1Dcon_main2_1MyTrue_1MyFalse_d;
  logic arg0_1Dcon_main2_1MyTrue_1MyFalse_r;
  MyBool_t arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d;
  logic arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_r;
  Go_t arg0_2Dcon_main2_d;
  logic arg0_2Dcon_main2_r;
  Int_t arg0_2_1Dcon_main1_d;
  logic arg0_2_1Dcon_main1_r;
  Int_t arg0_2_1Dcon_main1_1_d;
  logic arg0_2_1Dcon_main1_1_r;
  Int_t arg0_2_1Dcon_main1_2_d;
  logic arg0_2_1Dcon_main1_2_r;
  Int_t arg0_2_1Dcon_main1_3_d;
  logic arg0_2_1Dcon_main1_3_r;
  Int_t arg0_2_1Dcon_main1_4_d;
  logic arg0_2_1Dcon_main1_4_r;
  \Int#_t  x1ajF_destruct_d;
  logic x1ajF_destruct_r;
  Int_t \arg0_2_1Dcon_main1_1I#_d ;
  logic \arg0_2_1Dcon_main1_1I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_d ;
  logic \arg0_2_1Dcon_main1_3I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_2_d ;
  logic \arg0_2_1Dcon_main1_3I#_2_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_3_d ;
  logic \arg0_2_1Dcon_main1_3I#_3_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_2_1Dcon_main1_3I#_1_argbuf_0_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet2_1wild1XF_1_Eq_d;
  logic lizzieLet2_1wild1XF_1_Eq_r;
  Go_t \arg0_2_1Dcon_main1_3I#_2_argbuf_d ;
  logic \arg0_2_1Dcon_main1_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d;
  logic lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_r;
  Go_t arg0_2_2Dcon_main1_d;
  logic arg0_2_2Dcon_main1_r;
  MyBool_t lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_d;
  logic lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_r;
  MyBool_t arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_d;
  logic arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_r;
  Int_t \arg0_4_1Dcon_$fNumInt_$c+_d ;
  logic \arg0_4_1Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_4_r ;
  \Int#_t  xa1lV_destruct_d;
  logic xa1lV_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_1I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r ;
  \Int#_t  ya1lW_destruct_d;
  logic ya1lW_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d ;
  logic \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r ;
  Int_t \es_0_2_1I#_d ;
  logic \es_0_2_1I#_r ;
  Int_t \es_0_2_1I#_mux_d ;
  logic \es_0_2_1I#_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_mux_r ;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  MyBool_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_r;
  MyDTInt_Int_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_r;
  Pointer_QTree_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_r;
  Pointer_QTree_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_r;
  Pointer_CT$wmAdd_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r;
  Go_t call_$wmAdd_Int_initBufi_d;
  logic call_$wmAdd_Int_initBufi_r;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t call_$wmAdd_Int_unlockFork1_d;
  logic call_$wmAdd_Int_unlockFork1_r;
  Go_t call_$wmAdd_Int_unlockFork2_d;
  logic call_$wmAdd_Int_unlockFork2_r;
  Go_t call_$wmAdd_Int_unlockFork3_d;
  logic call_$wmAdd_Int_unlockFork3_r;
  Go_t call_$wmAdd_Int_unlockFork4_d;
  logic call_$wmAdd_Int_unlockFork4_r;
  Go_t call_$wmAdd_Int_unlockFork5_d;
  logic call_$wmAdd_Int_unlockFork5_r;
  Go_t call_$wmAdd_Int_initBuf_d;
  logic call_$wmAdd_Int_initBuf_r;
  Go_t call_$wmAdd_Int_goMux1_d;
  logic call_$wmAdd_Int_goMux1_r;
  MyDTInt_Int_Int_t call_$wmAdd_Int_goMux2_d;
  logic call_$wmAdd_Int_goMux2_r;
  Pointer_QTree_Int_t call_$wmAdd_Int_goMux3_d;
  logic call_$wmAdd_Int_goMux3_r;
  Pointer_QTree_Int_t call_$wmAdd_Int_goMux4_d;
  logic call_$wmAdd_Int_goMux4_r;
  Pointer_CT$wmAdd_Int_t call_$wmAdd_Int_goMux5_d;
  logic call_$wmAdd_Int_goMux5_r;
  Go_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_r;
  Pointer_QTree_Bool_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_r;
  Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_r;
  Go_t call_$wnnz_initBufi_d;
  logic call_$wnnz_initBufi_r;
  C5_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t call_$wnnz_unlockFork1_d;
  logic call_$wnnz_unlockFork1_r;
  Go_t call_$wnnz_unlockFork2_d;
  logic call_$wnnz_unlockFork2_r;
  Go_t call_$wnnz_unlockFork3_d;
  logic call_$wnnz_unlockFork3_r;
  Go_t call_$wnnz_initBuf_d;
  logic call_$wnnz_initBuf_r;
  Go_t call_$wnnz_goMux1_d;
  logic call_$wnnz_goMux1_r;
  Pointer_QTree_Bool_t call_$wnnz_goMux2_d;
  logic call_$wnnz_goMux2_r;
  Pointer_CT$wnnz_t call_$wnnz_goMux3_d;
  logic call_$wnnz_goMux3_r;
  Go_t \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_r ;
  MyDTBool_Bool_t \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_r ;
  MyDTInt_Bool_t \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_r ;
  Pointer_QTree_Int_t \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_r ;
  Go_t \call_main_map'_Int_Bool_initBufi_d ;
  logic \call_main_map'_Int_Bool_initBufi_r ;
  C5_t go_13_goMux_choice_d;
  logic go_13_goMux_choice_r;
  Go_t go_13_goMux_data_d;
  logic go_13_goMux_data_r;
  Go_t \call_main_map'_Int_Bool_unlockFork1_d ;
  logic \call_main_map'_Int_Bool_unlockFork1_r ;
  Go_t \call_main_map'_Int_Bool_unlockFork2_d ;
  logic \call_main_map'_Int_Bool_unlockFork2_r ;
  Go_t \call_main_map'_Int_Bool_unlockFork3_d ;
  logic \call_main_map'_Int_Bool_unlockFork3_r ;
  Go_t \call_main_map'_Int_Bool_unlockFork4_d ;
  logic \call_main_map'_Int_Bool_unlockFork4_r ;
  Go_t \call_main_map'_Int_Bool_unlockFork5_d ;
  logic \call_main_map'_Int_Bool_unlockFork5_r ;
  Go_t \call_main_map'_Int_Bool_initBuf_d ;
  logic \call_main_map'_Int_Bool_initBuf_r ;
  Go_t \call_main_map'_Int_Bool_goMux1_d ;
  logic \call_main_map'_Int_Bool_goMux1_r ;
  MyDTBool_Bool_t \call_main_map'_Int_Bool_goMux2_d ;
  logic \call_main_map'_Int_Bool_goMux2_r ;
  MyDTInt_Bool_t \call_main_map'_Int_Bool_goMux3_d ;
  logic \call_main_map'_Int_Bool_goMux3_r ;
  Pointer_QTree_Int_t \call_main_map'_Int_Bool_goMux4_d ;
  logic \call_main_map'_Int_Bool_goMux4_r ;
  \Pointer_CTmain_map'_Int_Bool_t  \call_main_map'_Int_Bool_goMux5_d ;
  logic \call_main_map'_Int_Bool_goMux5_r ;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Go_t es_0_4_1MyFalse_d;
  logic es_0_4_1MyFalse_r;
  Go_t es_0_4_1MyTrue_d;
  logic es_0_4_1MyTrue_r;
  Go_t es_0_4_1MyFalse_1_argbuf_d;
  logic es_0_4_1MyFalse_1_argbuf_r;
  Go_t es_0_4_1MyTrue_1_d;
  logic es_0_4_1MyTrue_1_r;
  Go_t es_0_4_1MyTrue_2_d;
  logic es_0_4_1MyTrue_2_r;
  QTree_Bool_t es_0_4_1MyTrue_1QNone_Bool_d;
  logic es_0_4_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Go_t es_0_4_1MyTrue_2_argbuf_d;
  logic es_0_4_1MyTrue_2_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyFalse_d;
  logic es_0_4_2MyFalse_r;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyTrue_d;
  logic es_0_4_2MyTrue_r;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyFalse_1_argbuf_d;
  logic es_0_4_2MyFalse_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyTrue_1_argbuf_d;
  logic es_0_4_2MyTrue_1_argbuf_r;
  MyBool_t es_0_4_3MyFalse_d;
  logic es_0_4_3MyFalse_r;
  MyBool_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  QTree_Bool_t es_0_4_3MyFalse_1QVal_Bool_d;
  logic es_0_4_3MyFalse_1QVal_Bool_r;
  QTree_Bool_t lizzieLet19_1_argbuf_d;
  logic lizzieLet19_1_argbuf_r;
  \Int#_t  contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  \Int#_t  es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_d;
  logic es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_r;
  MyDTInt_Bool_t ga8L_2_2_argbuf_d;
  logic ga8L_2_2_argbuf_r;
  MyDTInt_Bool_t ga8L_2_1_d;
  logic ga8L_2_1_r;
  MyDTInt_Bool_t ga8L_2_2_d;
  logic ga8L_2_2_r;
  MyDTInt_Bool_t ga8L_3_2_argbuf_d;
  logic ga8L_3_2_argbuf_r;
  MyDTInt_Bool_t ga8L_3_1_d;
  logic ga8L_3_1_r;
  MyDTInt_Bool_t ga8L_3_2_d;
  logic ga8L_3_2_r;
  MyDTInt_Bool_t ga8L_4_1_argbuf_d;
  logic ga8L_4_1_argbuf_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  C5_t go_11_goMux_choice_3_d;
  logic go_11_goMux_choice_3_r;
  C5_t go_11_goMux_choice_4_d;
  logic go_11_goMux_choice_4_r;
  MyDTInt_Int_Int_t wslR_1_goMux_mux_d;
  logic wslR_1_goMux_mux_r;
  Pointer_QTree_Int_t w1slS_1_goMux_mux_d;
  logic w1slS_1_goMux_mux_r;
  Pointer_QTree_Int_t w2slT_1_goMux_mux_d;
  logic w2slT_1_goMux_mux_r;
  Pointer_CT$wmAdd_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C5_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  Pointer_QTree_Bool_t wslW_1_goMux_mux_d;
  logic wslW_1_goMux_mux_r;
  Pointer_CT$wnnz_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_13_goMux_choice_1_d;
  logic go_13_goMux_choice_1_r;
  C5_t go_13_goMux_choice_2_d;
  logic go_13_goMux_choice_2_r;
  C5_t go_13_goMux_choice_3_d;
  logic go_13_goMux_choice_3_r;
  C5_t go_13_goMux_choice_4_d;
  logic go_13_goMux_choice_4_r;
  MyDTBool_Bool_t isZa8K_goMux_mux_d;
  logic isZa8K_goMux_mux_r;
  MyDTInt_Bool_t ga8L_goMux_mux_d;
  logic ga8L_goMux_mux_r;
  Pointer_QTree_Int_t ma8M_goMux_mux_d;
  logic ma8M_goMux_mux_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  \CTmain_map'_Int_Bool_t  \go_14_1Lmain_map'_Int_Boolsbos_d ;
  logic \go_14_1Lmain_map'_Int_Boolsbos_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t go_14_2_argbuf_d;
  logic go_14_2_argbuf_r;
  \TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_t  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d ;
  logic \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_r ;
  C10_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C10_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C4_t go_16_goMux_choice_1_d;
  logic go_16_goMux_choice_1_r;
  C4_t go_16_goMux_choice_2_d;
  logic go_16_goMux_choice_2_r;
  \Int#_t  srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CT$wnnz_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C5_t go_17_goMux_choice_1_d;
  logic go_17_goMux_choice_1_r;
  C5_t go_17_goMux_choice_2_d;
  logic go_17_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTmain_map'_Int_Bool_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r ;
  CT$wmAdd_Int_t go_6_1L$wmAdd_Intsbos_d;
  logic go_6_1L$wmAdd_Intsbos_r;
  CT$wmAdd_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_t call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d;
  logic call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r;
  MyDTInt_Bool_t go_7_1Dcon_main1_d;
  logic go_7_1Dcon_main1_r;
  MyDTInt_Bool_t es_2_1_argbuf_d;
  logic es_2_1_argbuf_r;
  MyDTBool_Bool_t go_7_2Dcon_main2_d;
  logic go_7_2Dcon_main2_r;
  MyDTBool_Bool_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$c+_d ;
  logic \go_7_3Dcon_$fNumInt_$c+_r ;
  MyDTInt_Int_Int_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  Go_t go_7_4_argbuf_d;
  logic go_7_4_argbuf_r;
  TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r ;
  Go_t go_7_5_argbuf_d;
  logic go_7_5_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_r ;
  Go_t go_7_6_argbuf_d;
  logic go_7_6_argbuf_r;
  TupGo___Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_Bool_1_d ;
  logic \$wnnzTupGo___Pointer_QTree_Bool_1_r ;
  CT$wnnz_t go_8_1L$wnnzsbos_d;
  logic go_8_1L$wnnzsbos_r;
  CT$wnnz_t lizzieLet1_1_argbuf_d;
  logic lizzieLet1_1_argbuf_r;
  Go_t go_8_2_argbuf_d;
  logic go_8_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_t call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d;
  logic call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r;
  MyDTBool_Bool_t isZa8K_2_2_argbuf_d;
  logic isZa8K_2_2_argbuf_r;
  MyDTBool_Bool_t isZa8K_2_1_d;
  logic isZa8K_2_1_r;
  MyDTBool_Bool_t isZa8K_2_2_d;
  logic isZa8K_2_2_r;
  MyDTBool_Bool_t isZa8K_3_2_argbuf_d;
  logic isZa8K_3_2_argbuf_r;
  MyDTBool_Bool_t isZa8K_3_1_d;
  logic isZa8K_3_1_r;
  MyDTBool_Bool_t isZa8K_3_2_d;
  logic isZa8K_3_2_r;
  MyDTBool_Bool_t isZa8K_4_1_argbuf_d;
  logic isZa8K_4_1_argbuf_r;
  Pointer_QTree_Bool_t q1a92_destruct_d;
  logic q1a92_destruct_r;
  Pointer_QTree_Bool_t q2a93_destruct_d;
  logic q2a93_destruct_r;
  Pointer_QTree_Bool_t q3a94_destruct_d;
  logic q3a94_destruct_r;
  Pointer_QTree_Bool_t q4a95_destruct_d;
  logic q4a95_destruct_r;
  QTree_Bool_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  QTree_Bool_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  QTree_Bool_t lizzieLet15_1QNode_Bool_d;
  logic lizzieLet15_1QNode_Bool_r;
  QTree_Bool_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Go_t lizzieLet15_3QNone_Bool_d;
  logic lizzieLet15_3QNone_Bool_r;
  Go_t lizzieLet15_3QVal_Bool_d;
  logic lizzieLet15_3QVal_Bool_r;
  Go_t lizzieLet15_3QNode_Bool_d;
  logic lizzieLet15_3QNode_Bool_r;
  Go_t lizzieLet15_3QError_Bool_d;
  logic lizzieLet15_3QError_Bool_r;
  Go_t lizzieLet15_3QError_Bool_1_d;
  logic lizzieLet15_3QError_Bool_1_r;
  Go_t lizzieLet15_3QError_Bool_2_d;
  logic lizzieLet15_3QError_Bool_2_r;
  Go_t lizzieLet15_3QError_Bool_1_argbuf_d;
  logic lizzieLet15_3QError_Bool_1_argbuf_r;
  \Int#_t  lizzieLet15_3QError_Bool_1_argbuf_0_d;
  logic lizzieLet15_3QError_Bool_1_argbuf_0_r;
  \Int#_t  lizzieLet5_2_1_argbuf_d;
  logic lizzieLet5_2_1_argbuf_r;
  Go_t lizzieLet15_3QError_Bool_2_argbuf_d;
  logic lizzieLet15_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet15_3QNode_Bool_1_argbuf_d;
  logic lizzieLet15_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet15_3QNone_Bool_1_d;
  logic lizzieLet15_3QNone_Bool_1_r;
  Go_t lizzieLet15_3QNone_Bool_2_d;
  logic lizzieLet15_3QNone_Bool_2_r;
  Go_t lizzieLet15_3QNone_Bool_1_argbuf_d;
  logic lizzieLet15_3QNone_Bool_1_argbuf_r;
  \Int#_t  lizzieLet15_3QNone_Bool_1_argbuf_0_d;
  logic lizzieLet15_3QNone_Bool_1_argbuf_0_r;
  \Int#_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Go_t lizzieLet15_3QNone_Bool_2_argbuf_d;
  logic lizzieLet15_3QNone_Bool_2_argbuf_r;
  C4_t go_16_goMux_choice_d;
  logic go_16_goMux_choice_r;
  Go_t go_16_goMux_data_d;
  logic go_16_goMux_data_r;
  Go_t lizzieLet15_3QVal_Bool_1_d;
  logic lizzieLet15_3QVal_Bool_1_r;
  Go_t lizzieLet15_3QVal_Bool_2_d;
  logic lizzieLet15_3QVal_Bool_2_r;
  Go_t lizzieLet15_3QVal_Bool_1_argbuf_d;
  logic lizzieLet15_3QVal_Bool_1_argbuf_r;
  \Int#_t  lizzieLet15_3QVal_Bool_1_argbuf_1_d;
  logic lizzieLet15_3QVal_Bool_1_argbuf_1_r;
  \Int#_t  lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Go_t lizzieLet15_3QVal_Bool_2_argbuf_d;
  logic lizzieLet15_3QVal_Bool_2_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet15_4QNone_Bool_d;
  logic lizzieLet15_4QNone_Bool_r;
  Pointer_CT$wnnz_t lizzieLet15_4QVal_Bool_d;
  logic lizzieLet15_4QVal_Bool_r;
  Pointer_CT$wnnz_t lizzieLet15_4QNode_Bool_d;
  logic lizzieLet15_4QNode_Bool_r;
  Pointer_CT$wnnz_t lizzieLet15_4QError_Bool_d;
  logic lizzieLet15_4QError_Bool_r;
  Pointer_CT$wnnz_t lizzieLet15_4QError_Bool_1_argbuf_d;
  logic lizzieLet15_4QError_Bool_1_argbuf_r;
  CT$wnnz_t lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_d;
  logic lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet15_4QNone_Bool_1_argbuf_d;
  logic lizzieLet15_4QNone_Bool_1_argbuf_r;
  Pointer_CT$wnnz_t lizzieLet15_4QVal_Bool_1_argbuf_d;
  logic lizzieLet15_4QVal_Bool_1_argbuf_r;
  Pointer_QTree_Int_t q1a8O_destruct_d;
  logic q1a8O_destruct_r;
  Pointer_QTree_Int_t q2a8P_destruct_d;
  logic q2a8P_destruct_r;
  Pointer_QTree_Int_t q3a8Q_destruct_d;
  logic q3a8Q_destruct_r;
  Pointer_QTree_Int_t q4a8R_destruct_d;
  logic q4a8R_destruct_r;
  Int_t va8N_destruct_d;
  logic va8N_destruct_r;
  QTree_Int_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  QTree_Int_t lizzieLet17_1QVal_Int_d;
  logic lizzieLet17_1QVal_Int_r;
  QTree_Int_t lizzieLet17_1QNode_Int_d;
  logic lizzieLet17_1QNode_Int_r;
  QTree_Int_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  MyDTInt_Bool_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_3QVal_Int_d;
  logic lizzieLet17_3QVal_Int_r;
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_d;
  logic lizzieLet17_3QNode_Int_r;
  MyDTInt_Bool_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_1_d;
  logic lizzieLet17_3QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_2_d;
  logic lizzieLet17_3QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_2_argbuf_d;
  logic lizzieLet17_3QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet17_3QVal_Int_1_argbuf_d;
  logic lizzieLet17_3QVal_Int_1_argbuf_r;
  Go_t lizzieLet17_4QNone_Int_d;
  logic lizzieLet17_4QNone_Int_r;
  Go_t lizzieLet17_4QVal_Int_d;
  logic lizzieLet17_4QVal_Int_r;
  Go_t lizzieLet17_4QNode_Int_d;
  logic lizzieLet17_4QNode_Int_r;
  Go_t lizzieLet17_4QError_Int_d;
  logic lizzieLet17_4QError_Int_r;
  Go_t lizzieLet17_4QError_Int_1_d;
  logic lizzieLet17_4QError_Int_1_r;
  Go_t lizzieLet17_4QError_Int_2_d;
  logic lizzieLet17_4QError_Int_2_r;
  QTree_Bool_t lizzieLet17_4QError_Int_1QError_Bool_d;
  logic lizzieLet17_4QError_Int_1QError_Bool_r;
  QTree_Bool_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t lizzieLet17_4QError_Int_2_argbuf_d;
  logic lizzieLet17_4QError_Int_2_argbuf_r;
  Go_t lizzieLet17_4QNode_Int_1_argbuf_d;
  logic lizzieLet17_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet17_4QNone_Int_1_d;
  logic lizzieLet17_4QNone_Int_1_r;
  Go_t lizzieLet17_4QNone_Int_2_d;
  logic lizzieLet17_4QNone_Int_2_r;
  QTree_Bool_t lizzieLet17_4QNone_Int_1QNone_Bool_d;
  logic lizzieLet17_4QNone_Int_1QNone_Bool_r;
  QTree_Bool_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t lizzieLet17_4QNone_Int_2_argbuf_d;
  logic lizzieLet17_4QNone_Int_2_argbuf_r;
  C5_t go_17_goMux_choice_d;
  logic go_17_goMux_choice_r;
  Go_t go_17_goMux_data_d;
  logic go_17_goMux_data_r;
  Go_t lizzieLet17_4QVal_Int_1_d;
  logic lizzieLet17_4QVal_Int_1_r;
  Go_t lizzieLet17_4QVal_Int_2_d;
  logic lizzieLet17_4QVal_Int_2_r;
  Go_t lizzieLet17_4QVal_Int_3_d;
  logic lizzieLet17_4QVal_Int_3_r;
  Go_t lizzieLet17_4QVal_Int_1_argbuf_d;
  logic lizzieLet17_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  Go_t lizzieLet17_4QVal_Int_2_argbuf_d;
  logic lizzieLet17_4QVal_Int_2_argbuf_r;
  TupGo___MyDTBool_Bool___MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r;
  MyDTBool_Bool_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  MyDTBool_Bool_t lizzieLet17_5QVal_Int_d;
  logic lizzieLet17_5QVal_Int_r;
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_d;
  logic lizzieLet17_5QNode_Int_r;
  MyDTBool_Bool_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_1_d;
  logic lizzieLet17_5QNode_Int_1_r;
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_2_d;
  logic lizzieLet17_5QNode_Int_2_r;
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_2_argbuf_d;
  logic lizzieLet17_5QNode_Int_2_argbuf_r;
  MyDTBool_Bool_t lizzieLet17_5QVal_Int_1_argbuf_d;
  logic lizzieLet17_5QVal_Int_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QNone_Int_d;
  logic lizzieLet17_6QNone_Int_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QVal_Int_d;
  logic lizzieLet17_6QVal_Int_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QNode_Int_d;
  logic lizzieLet17_6QNode_Int_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QError_Int_d;
  logic lizzieLet17_6QError_Int_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QError_Int_1_argbuf_d;
  logic lizzieLet17_6QError_Int_1_argbuf_r;
  \CTmain_map'_Int_Bool_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_d ;
  logic \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QNone_Int_1_argbuf_d;
  logic lizzieLet17_6QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_QTree_Int_t es_4_3_destruct_d;
  logic es_4_3_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Int_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_QTree_Int_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  MyDTInt_Int_Int_t wslR_4_destruct_d;
  logic wslR_4_destruct_r;
  Pointer_QTree_Int_t q1a8j_3_destruct_d;
  logic q1a8j_3_destruct_r;
  Pointer_QTree_Int_t t1a8o_3_destruct_d;
  logic t1a8o_3_destruct_r;
  Pointer_QTree_Int_t es_4_1_destruct_d;
  logic es_4_1_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  MyDTInt_Int_Int_t wslR_3_destruct_d;
  logic wslR_3_destruct_r;
  Pointer_QTree_Int_t q1a8j_2_destruct_d;
  logic q1a8j_2_destruct_r;
  Pointer_QTree_Int_t t1a8o_2_destruct_d;
  logic t1a8o_2_destruct_r;
  Pointer_QTree_Int_t q2a8k_2_destruct_d;
  logic q2a8k_2_destruct_r;
  Pointer_QTree_Int_t t2a8p_2_destruct_d;
  logic t2a8p_2_destruct_r;
  Pointer_CT$wmAdd_Int_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  MyDTInt_Int_Int_t wslR_2_destruct_d;
  logic wslR_2_destruct_r;
  Pointer_QTree_Int_t q1a8j_1_destruct_d;
  logic q1a8j_1_destruct_r;
  Pointer_QTree_Int_t t1a8o_1_destruct_d;
  logic t1a8o_1_destruct_r;
  Pointer_QTree_Int_t q2a8k_1_destruct_d;
  logic q2a8k_1_destruct_r;
  Pointer_QTree_Int_t t2a8p_1_destruct_d;
  logic t2a8p_1_destruct_r;
  Pointer_QTree_Int_t q3a8l_1_destruct_d;
  logic q3a8l_1_destruct_r;
  Pointer_QTree_Int_t t3a8q_1_destruct_d;
  logic t3a8q_1_destruct_r;
  CT$wmAdd_Int_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  CT$wmAdd_Int_t lizzieLet24_1Lcall_$wmAdd_Int3_d;
  logic lizzieLet24_1Lcall_$wmAdd_Int3_r;
  CT$wmAdd_Int_t lizzieLet24_1Lcall_$wmAdd_Int2_d;
  logic lizzieLet24_1Lcall_$wmAdd_Int2_r;
  CT$wmAdd_Int_t lizzieLet24_1Lcall_$wmAdd_Int1_d;
  logic lizzieLet24_1Lcall_$wmAdd_Int1_r;
  CT$wmAdd_Int_t lizzieLet24_1Lcall_$wmAdd_Int0_d;
  logic lizzieLet24_1Lcall_$wmAdd_Int0_r;
  Go_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int3_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int3_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int2_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int2_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int1_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int1_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int0_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int0_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet24_4L$wmAdd_Intsbos_d;
  logic lizzieLet24_4L$wmAdd_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int3_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int3_r;
  Pointer_QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int2_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int2_r;
  Pointer_QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int1_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int1_r;
  Pointer_QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int0_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int0_r;
  Pointer_QTree_Int_t lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wmAdd_Int_goConst_d;
  logic call_$wmAdd_Int_goConst_r;
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_d ;
  logic \$wmAdd_Int_resbuf_r ;
  QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_r;
  QTree_Int_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_r;
  CT$wmAdd_Int_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_r;
  CT$wmAdd_Int_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_r;
  CT$wmAdd_Int_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  \Int#_t  wwslZ_3_destruct_d;
  logic wwslZ_3_destruct_r;
  \Int#_t  ww1XmJ_2_destruct_d;
  logic ww1XmJ_2_destruct_r;
  \Int#_t  ww2XmM_1_destruct_d;
  logic ww2XmM_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  \Int#_t  wwslZ_2_destruct_d;
  logic wwslZ_2_destruct_r;
  \Int#_t  ww1XmJ_1_destruct_d;
  logic ww1XmJ_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Bool_t q4a95_3_destruct_d;
  logic q4a95_3_destruct_r;
  \Int#_t  wwslZ_1_destruct_d;
  logic wwslZ_1_destruct_r;
  Pointer_CT$wnnz_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Bool_t q4a95_2_destruct_d;
  logic q4a95_2_destruct_r;
  Pointer_QTree_Bool_t q3a94_2_destruct_d;
  logic q3a94_2_destruct_r;
  Pointer_CT$wnnz_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Bool_t q4a95_1_destruct_d;
  logic q4a95_1_destruct_r;
  Pointer_QTree_Bool_t q3a94_1_destruct_d;
  logic q3a94_1_destruct_r;
  Pointer_QTree_Bool_t q2a93_1_destruct_d;
  logic q2a93_1_destruct_r;
  CT$wnnz_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  CT$wnnz_t lizzieLet29_1Lcall_$wnnz3_d;
  logic lizzieLet29_1Lcall_$wnnz3_r;
  CT$wnnz_t lizzieLet29_1Lcall_$wnnz2_d;
  logic lizzieLet29_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet29_1Lcall_$wnnz1_d;
  logic lizzieLet29_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet29_1Lcall_$wnnz0_d;
  logic lizzieLet29_1Lcall_$wnnz0_r;
  Go_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Go_t lizzieLet29_3Lcall_$wnnz3_d;
  logic lizzieLet29_3Lcall_$wnnz3_r;
  Go_t lizzieLet29_3Lcall_$wnnz2_d;
  logic lizzieLet29_3Lcall_$wnnz2_r;
  Go_t lizzieLet29_3Lcall_$wnnz1_d;
  logic lizzieLet29_3Lcall_$wnnz1_r;
  Go_t lizzieLet29_3Lcall_$wnnz0_d;
  logic lizzieLet29_3Lcall_$wnnz0_r;
  Go_t lizzieLet29_3Lcall_$wnnz0_1_argbuf_d;
  logic lizzieLet29_3Lcall_$wnnz0_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_$wnnz1_1_argbuf_d;
  logic lizzieLet29_3Lcall_$wnnz1_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_$wnnz2_1_argbuf_d;
  logic lizzieLet29_3Lcall_$wnnz2_1_argbuf_r;
  Go_t lizzieLet29_3Lcall_$wnnz3_1_argbuf_d;
  logic lizzieLet29_3Lcall_$wnnz3_1_argbuf_r;
  \Int#_t  lizzieLet29_4L$wnnzsbos_d;
  logic lizzieLet29_4L$wnnzsbos_r;
  \Int#_t  lizzieLet29_4Lcall_$wnnz3_d;
  logic lizzieLet29_4Lcall_$wnnz3_r;
  \Int#_t  lizzieLet29_4Lcall_$wnnz2_d;
  logic lizzieLet29_4Lcall_$wnnz2_r;
  \Int#_t  lizzieLet29_4Lcall_$wnnz1_d;
  logic lizzieLet29_4Lcall_$wnnz1_r;
  \Int#_t  lizzieLet29_4Lcall_$wnnz0_d;
  logic lizzieLet29_4Lcall_$wnnz0_r;
  \Int#_t  lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_d;
  logic lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_d;
  logic lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_goConst_d;
  logic call_$wnnz_goConst_r;
  \Int#_t  \$wnnz_resbuf_d ;
  logic \$wnnz_resbuf_r ;
  CT$wnnz_t lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_d;
  logic lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_r;
  CT$wnnz_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Bool_t lizzieLet3_1_argbuf_d;
  logic lizzieLet3_1_argbuf_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_QTree_Bool_t es_4_7_destruct_d;
  logic es_4_7_destruct_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_QTree_Bool_t es_4_6_destruct_d;
  logic es_4_6_destruct_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  MyDTBool_Bool_t isZa8K_4_destruct_d;
  logic isZa8K_4_destruct_r;
  MyDTInt_Bool_t ga8L_4_destruct_d;
  logic ga8L_4_destruct_r;
  Pointer_QTree_Int_t q1a8O_3_destruct_d;
  logic q1a8O_3_destruct_r;
  Pointer_QTree_Bool_t es_4_5_destruct_d;
  logic es_4_5_destruct_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  MyDTBool_Bool_t isZa8K_3_destruct_d;
  logic isZa8K_3_destruct_r;
  MyDTInt_Bool_t ga8L_3_destruct_d;
  logic ga8L_3_destruct_r;
  Pointer_QTree_Int_t q1a8O_2_destruct_d;
  logic q1a8O_2_destruct_r;
  Pointer_QTree_Int_t q2a8P_2_destruct_d;
  logic q2a8P_2_destruct_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  MyDTBool_Bool_t isZa8K_2_destruct_d;
  logic isZa8K_2_destruct_r;
  MyDTInt_Bool_t ga8L_2_destruct_d;
  logic ga8L_2_destruct_r;
  Pointer_QTree_Int_t q1a8O_1_destruct_d;
  logic q1a8O_1_destruct_r;
  Pointer_QTree_Int_t q2a8P_1_destruct_d;
  logic q2a8P_1_destruct_r;
  Pointer_QTree_Int_t q3a8Q_1_destruct_d;
  logic q3a8Q_1_destruct_r;
  \CTmain_map'_Int_Bool_t  _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_1Lcall_main_map'_Int_Bool3_d ;
  logic \lizzieLet33_1Lcall_main_map'_Int_Bool3_r ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_1Lcall_main_map'_Int_Bool2_d ;
  logic \lizzieLet33_1Lcall_main_map'_Int_Bool2_r ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_1Lcall_main_map'_Int_Bool1_d ;
  logic \lizzieLet33_1Lcall_main_map'_Int_Bool1_r ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_1Lcall_main_map'_Int_Bool0_d ;
  logic \lizzieLet33_1Lcall_main_map'_Int_Bool0_r ;
  Go_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool3_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool3_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool2_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool2_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool1_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool1_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool0_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool0_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_r ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lmain_map'_Int_Boolsbos_d ;
  logic \lizzieLet33_4Lmain_map'_Int_Boolsbos_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool3_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool3_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool2_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool2_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool1_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool1_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool0_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool0_r ;
  QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet34_1_argbuf_d;
  logic lizzieLet34_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_r ;
  Go_t \call_main_map'_Int_Bool_goConst_d ;
  logic \call_main_map'_Int_Bool_goConst_r ;
  Pointer_QTree_Bool_t \main_map'_Int_Bool_resbuf_d ;
  logic \main_map'_Int_Bool_resbuf_r ;
  Go_t lizzieLet4_1MyFalse_d;
  logic lizzieLet4_1MyFalse_r;
  Go_t lizzieLet4_1MyTrue_d;
  logic lizzieLet4_1MyTrue_r;
  MyBool_t lizzieLet4_1MyFalse_1MyTrue_d;
  logic lizzieLet4_1MyFalse_1MyTrue_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t lizzieLet4_1MyTrue_1MyFalse_d;
  logic lizzieLet4_1MyTrue_1MyFalse_r;
  MyBool_t lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d;
  logic lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_r;
  Pointer_QTree_Int_t q1a8j_destruct_d;
  logic q1a8j_destruct_r;
  Pointer_QTree_Int_t q2a8k_destruct_d;
  logic q2a8k_destruct_r;
  Pointer_QTree_Int_t q3a8l_destruct_d;
  logic q3a8l_destruct_r;
  Pointer_QTree_Int_t q4a8m_destruct_d;
  logic q4a8m_destruct_r;
  Int_t v1a8d_destruct_d;
  logic v1a8d_destruct_r;
  QTree_Int_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  QTree_Int_t lizzieLet5_1QVal_Int_d;
  logic lizzieLet5_1QVal_Int_r;
  QTree_Int_t lizzieLet5_1QNode_Int_d;
  logic lizzieLet5_1QNode_Int_r;
  QTree_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Go_t lizzieLet5_3QNone_Int_d;
  logic lizzieLet5_3QNone_Int_r;
  Go_t lizzieLet5_3QVal_Int_d;
  logic lizzieLet5_3QVal_Int_r;
  Go_t lizzieLet5_3QNode_Int_d;
  logic lizzieLet5_3QNode_Int_r;
  Go_t lizzieLet5_3QError_Int_d;
  logic lizzieLet5_3QError_Int_r;
  Go_t lizzieLet5_3QError_Int_1_d;
  logic lizzieLet5_3QError_Int_1_r;
  Go_t lizzieLet5_3QError_Int_2_d;
  logic lizzieLet5_3QError_Int_2_r;
  QTree_Int_t lizzieLet5_3QError_Int_1QError_Int_d;
  logic lizzieLet5_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Go_t lizzieLet5_3QError_Int_2_argbuf_d;
  logic lizzieLet5_3QError_Int_2_argbuf_r;
  Go_t lizzieLet5_3QNone_Int_1_argbuf_d;
  logic lizzieLet5_3QNone_Int_1_argbuf_r;
  C10_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  QTree_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  QTree_Int_t lizzieLet5_4QVal_Int_d;
  logic lizzieLet5_4QVal_Int_r;
  QTree_Int_t lizzieLet5_4QNode_Int_d;
  logic lizzieLet5_4QNode_Int_r;
  QTree_Int_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  QTree_Int_t lizzieLet5_4QNode_Int_1_d;
  logic lizzieLet5_4QNode_Int_1_r;
  QTree_Int_t lizzieLet5_4QNode_Int_2_d;
  logic lizzieLet5_4QNode_Int_2_r;
  QTree_Int_t lizzieLet5_4QNode_Int_3_d;
  logic lizzieLet5_4QNode_Int_3_r;
  QTree_Int_t lizzieLet5_4QNode_Int_4_d;
  logic lizzieLet5_4QNode_Int_4_r;
  QTree_Int_t lizzieLet5_4QNode_Int_5_d;
  logic lizzieLet5_4QNode_Int_5_r;
  QTree_Int_t lizzieLet5_4QNode_Int_6_d;
  logic lizzieLet5_4QNode_Int_6_r;
  QTree_Int_t lizzieLet5_4QNode_Int_7_d;
  logic lizzieLet5_4QNode_Int_7_r;
  QTree_Int_t lizzieLet5_4QNode_Int_8_d;
  logic lizzieLet5_4QNode_Int_8_r;
  QTree_Int_t lizzieLet5_4QNode_Int_9_d;
  logic lizzieLet5_4QNode_Int_9_r;
  QTree_Int_t lizzieLet5_4QNode_Int_10_d;
  logic lizzieLet5_4QNode_Int_10_r;
  Pointer_QTree_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_QTree_Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_10QNode_Int_d;
  logic lizzieLet5_4QNode_Int_10QNode_Int_r;
  Pointer_QTree_Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_r;
  Pointer_QTree_Int_t t1a8o_destruct_d;
  logic t1a8o_destruct_r;
  Pointer_QTree_Int_t t2a8p_destruct_d;
  logic t2a8p_destruct_r;
  Pointer_QTree_Int_t t3a8q_destruct_d;
  logic t3a8q_destruct_r;
  Pointer_QTree_Int_t t4a8r_destruct_d;
  logic t4a8r_destruct_r;
  QTree_Int_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  QTree_Int_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  QTree_Int_t lizzieLet5_4QNode_Int_1QNode_Int_d;
  logic lizzieLet5_4QNode_Int_1QNode_Int_r;
  QTree_Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Go_t lizzieLet5_4QNode_Int_3QNone_Int_d;
  logic lizzieLet5_4QNode_Int_3QNone_Int_r;
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_r;
  Go_t lizzieLet5_4QNode_Int_3QNode_Int_d;
  logic lizzieLet5_4QNode_Int_3QNode_Int_r;
  Go_t lizzieLet5_4QNode_Int_3QError_Int_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_r;
  Go_t lizzieLet5_4QNode_Int_3QError_Int_1_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_1_r;
  Go_t lizzieLet5_4QNode_Int_3QError_Int_2_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Go_t lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_1_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_1_r;
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_2_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_2_r;
  QTree_Int_t lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_r;
  QTree_Int_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNone_Int_d;
  logic lizzieLet5_4QNode_Int_4QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QVal_Int_d;
  logic lizzieLet5_4QNode_Int_4QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNode_Int_d;
  logic lizzieLet5_4QNode_Int_4QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QError_Int_d;
  logic lizzieLet5_4QNode_Int_4QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_r;
  CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_d;
  logic lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_r;
  CT$wmAdd_Int_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_5QNone_Int_d;
  logic lizzieLet5_4QNode_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_QTree_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  Pointer_QTree_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTInt_Int_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_d;
  logic lizzieLet5_4QNode_Int_6QNode_Int_r;
  MyDTInt_Int_Int_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_1_d;
  logic lizzieLet5_4QNode_Int_6QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_2_d;
  logic lizzieLet5_4QNode_Int_6QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_d;
  logic lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Int_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_7QNode_Int_d;
  logic lizzieLet5_4QNode_Int_7QNode_Int_r;
  Pointer_QTree_Int_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_8QNode_Int_d;
  logic lizzieLet5_4QNode_Int_8QNode_Int_r;
  Pointer_QTree_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Pointer_QTree_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Pointer_QTree_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_9QNode_Int_d;
  logic lizzieLet5_4QNode_Int_9QNode_Int_r;
  Pointer_QTree_Int_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  QTree_Int_t lizzieLet5_4QVal_Int_1_d;
  logic lizzieLet5_4QVal_Int_1_r;
  QTree_Int_t lizzieLet5_4QVal_Int_2_d;
  logic lizzieLet5_4QVal_Int_2_r;
  QTree_Int_t lizzieLet5_4QVal_Int_3_d;
  logic lizzieLet5_4QVal_Int_3_r;
  QTree_Int_t lizzieLet5_4QVal_Int_4_d;
  logic lizzieLet5_4QVal_Int_4_r;
  QTree_Int_t lizzieLet5_4QVal_Int_5_d;
  logic lizzieLet5_4QVal_Int_5_r;
  QTree_Int_t lizzieLet5_4QVal_Int_6_d;
  logic lizzieLet5_4QVal_Int_6_r;
  QTree_Int_t lizzieLet5_4QVal_Int_7_d;
  logic lizzieLet5_4QVal_Int_7_r;
  Int_t va8e_destruct_d;
  logic va8e_destruct_r;
  QTree_Int_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  QTree_Int_t lizzieLet5_4QVal_Int_1QVal_Int_d;
  logic lizzieLet5_4QVal_Int_1QVal_Int_r;
  QTree_Int_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  QTree_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Go_t lizzieLet5_4QVal_Int_3QNone_Int_d;
  logic lizzieLet5_4QVal_Int_3QNone_Int_r;
  Go_t lizzieLet5_4QVal_Int_3QVal_Int_d;
  logic lizzieLet5_4QVal_Int_3QVal_Int_r;
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_r;
  Go_t lizzieLet5_4QVal_Int_3QError_Int_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_r;
  Go_t lizzieLet5_4QVal_Int_3QError_Int_1_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_1_r;
  Go_t lizzieLet5_4QVal_Int_3QError_Int_2_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_2_r;
  QTree_Int_t lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Go_t lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_r;
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_1_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_1_r;
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_2_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_2_r;
  QTree_Int_t lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_r;
  QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_r;
  Go_t lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNone_Int_d;
  logic lizzieLet5_4QVal_Int_4QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QVal_Int_d;
  logic lizzieLet5_4QVal_Int_4QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNode_Int_d;
  logic lizzieLet5_4QVal_Int_4QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QError_Int_d;
  logic lizzieLet5_4QVal_Int_4QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet5_4QVal_Int_5QNone_Int_d;
  logic lizzieLet5_4QVal_Int_5QNone_Int_r;
  Pointer_QTree_Int_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_QTree_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  Pointer_QTree_Int_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet5_4QVal_Int_6QVal_Int_d;
  logic lizzieLet5_4QVal_Int_6QVal_Int_r;
  MyDTInt_Int_Int_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  MyDTInt_Int_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Int_t lizzieLet5_4QVal_Int_7QVal_Int_d;
  logic lizzieLet5_4QVal_Int_7QVal_Int_r;
  Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Int_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Int_t lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_d;
  logic lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QNone_Int_d;
  logic lizzieLet5_5QNone_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QVal_Int_d;
  logic lizzieLet5_5QVal_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QNode_Int_d;
  logic lizzieLet5_5QNode_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QError_Int_d;
  logic lizzieLet5_5QError_Int_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QError_Int_1_argbuf_d;
  logic lizzieLet5_5QError_Int_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QNone_Int_1_argbuf_d;
  logic lizzieLet5_5QNone_Int_1_argbuf_r;
  Pointer_QTree_Int_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_6QVal_Int_d;
  logic lizzieLet5_6QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet5_6QNode_Int_d;
  logic lizzieLet5_6QNode_Int_r;
  Pointer_QTree_Int_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_7QNone_Int_d;
  logic lizzieLet5_7QNone_Int_r;
  Pointer_QTree_Int_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_QTree_Int_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  Pointer_QTree_Int_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet5_7QNone_Int_1_argbuf_d;
  logic lizzieLet5_7QNone_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet5_8QVal_Int_d;
  logic lizzieLet5_8QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet5_8QNode_Int_d;
  logic lizzieLet5_8QNode_Int_r;
  MyDTInt_Int_Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Pointer_QTree_Int_t ma8M_1_argbuf_d;
  logic ma8M_1_argbuf_r;
  Go_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_r ;
  MyDTBool_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_r ;
  MyDTInt_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_r ;
  Pointer_QTree_Int_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_r ;
  MyDTInt_Bool_t ga8L_1_1_argbuf_d;
  logic ga8L_1_1_argbuf_r;
  Go_t go_14_1_d;
  logic go_14_1_r;
  Go_t go_14_2_d;
  logic go_14_2_r;
  MyDTBool_Bool_t isZa8K_1_1_argbuf_d;
  logic isZa8K_1_1_argbuf_r;
  Pointer_QTree_Int_t ma8M_1_1_argbuf_d;
  logic ma8M_1_1_argbuf_r;
  Pointer_QTree_Bool_t es_0_1_1_argbuf_d;
  logic es_0_1_1_argbuf_r;
  Pointer_QTree_Int_t q1a8O_3_1_argbuf_d;
  logic q1a8O_3_1_argbuf_r;
  Pointer_QTree_Int_t q1a8j_3_1_argbuf_d;
  logic q1a8j_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1a92_1_argbuf_d;
  logic q1a92_1_argbuf_r;
  Pointer_QTree_Int_t q2a8P_2_1_argbuf_d;
  logic q2a8P_2_1_argbuf_r;
  Pointer_QTree_Int_t q2a8k_2_1_argbuf_d;
  logic q2a8k_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2a93_1_1_argbuf_d;
  logic q2a93_1_1_argbuf_r;
  Pointer_QTree_Int_t q3a8Q_1_1_argbuf_d;
  logic q3a8Q_1_1_argbuf_r;
  Pointer_QTree_Int_t q3a8l_1_1_argbuf_d;
  logic q3a8l_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3a94_2_1_argbuf_d;
  logic q3a94_2_1_argbuf_r;
  Pointer_QTree_Int_t q4a8R_1_argbuf_d;
  logic q4a8R_1_argbuf_r;
  Pointer_QTree_Bool_t q4a95_3_1_argbuf_d;
  logic q4a95_3_1_argbuf_r;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r;
  CT$wmAdd_Int_t lizzieLet24_1_d;
  logic lizzieLet24_1_r;
  CT$wmAdd_Int_t lizzieLet24_2_d;
  logic lizzieLet24_2_r;
  CT$wmAdd_Int_t lizzieLet24_3_d;
  logic lizzieLet24_3_r;
  CT$wmAdd_Int_t lizzieLet24_4_d;
  logic lizzieLet24_4_r;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_r;
  CT$wnnz_t lizzieLet29_1_d;
  logic lizzieLet29_1_r;
  CT$wnnz_t lizzieLet29_2_d;
  logic lizzieLet29_2_r;
  CT$wnnz_t lizzieLet29_3_d;
  logic lizzieLet29_3_r;
  CT$wnnz_t lizzieLet29_4_d;
  logic lizzieLet29_4_r;
  \CTmain_map'_Int_Bool_t  \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_r ;
  \CTmain_map'_Int_Bool_t  lizzieLet33_1_d;
  logic lizzieLet33_1_r;
  \CTmain_map'_Int_Bool_t  lizzieLet33_2_d;
  logic lizzieLet33_2_r;
  \CTmain_map'_Int_Bool_t  lizzieLet33_3_d;
  logic lizzieLet33_3_r;
  \CTmain_map'_Int_Bool_t  lizzieLet33_4_d;
  logic lizzieLet33_4_r;
  QTree_Bool_t readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d;
  logic readPointer_QTree_BoolwslW_1_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet15_1_d;
  logic lizzieLet15_1_r;
  QTree_Bool_t lizzieLet15_2_d;
  logic lizzieLet15_2_r;
  QTree_Bool_t lizzieLet15_3_d;
  logic lizzieLet15_3_r;
  QTree_Bool_t lizzieLet15_4_d;
  logic lizzieLet15_4_r;
  QTree_Int_t readPointer_QTree_Intma8M_1_argbuf_rwb_d;
  logic readPointer_QTree_Intma8M_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet17_1_d;
  logic lizzieLet17_1_r;
  QTree_Int_t lizzieLet17_2_d;
  logic lizzieLet17_2_r;
  QTree_Int_t lizzieLet17_3_d;
  logic lizzieLet17_3_r;
  QTree_Int_t lizzieLet17_4_d;
  logic lizzieLet17_4_r;
  QTree_Int_t lizzieLet17_5_d;
  logic lizzieLet17_5_r;
  QTree_Int_t lizzieLet17_6_d;
  logic lizzieLet17_6_r;
  QTree_Int_t readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intw1slS_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet5_1_d;
  logic lizzieLet5_1_r;
  QTree_Int_t lizzieLet5_2_d;
  logic lizzieLet5_2_r;
  QTree_Int_t lizzieLet5_3_d;
  logic lizzieLet5_3_r;
  QTree_Int_t lizzieLet5_4_d;
  logic lizzieLet5_4_r;
  QTree_Int_t lizzieLet5_5_d;
  logic lizzieLet5_5_r;
  QTree_Int_t lizzieLet5_6_d;
  logic lizzieLet5_6_r;
  QTree_Int_t lizzieLet5_7_d;
  logic lizzieLet5_7_r;
  QTree_Int_t lizzieLet5_8_d;
  logic lizzieLet5_8_r;
  QTree_Int_t readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Intw2slT_1_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  Pointer_CT$wnnz_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Int_t t1a8o_3_1_argbuf_d;
  logic t1a8o_3_1_argbuf_r;
  Pointer_QTree_Int_t t2a8p_2_1_argbuf_d;
  logic t2a8p_2_1_argbuf_r;
  Pointer_QTree_Int_t t3a8q_1_1_argbuf_d;
  logic t3a8q_1_1_argbuf_r;
  Pointer_QTree_Int_t t4a8r_1_argbuf_d;
  logic t4a8r_1_argbuf_r;
  Int_t va8N_1_argbuf_d;
  logic va8N_1_argbuf_r;
  Int_t va8e_1_argbuf_d;
  logic va8e_1_argbuf_r;
  Pointer_QTree_Int_t w1slS_1_1_argbuf_d;
  logic w1slS_1_1_argbuf_r;
  Pointer_QTree_Int_t w1slS_1_1_d;
  logic w1slS_1_1_r;
  Pointer_QTree_Int_t w1slS_1_2_d;
  logic w1slS_1_2_r;
  Pointer_QTree_Int_t w2slT_1_1_argbuf_d;
  logic w2slT_1_1_argbuf_r;
  Pointer_QTree_Int_t w2slT_1_1_d;
  logic w2slT_1_1_r;
  Pointer_QTree_Int_t w2slT_1_2_d;
  logic w2slT_1_2_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_d;
  logic writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet16_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet1_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet30_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet31_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_rwb_d;
  logic writeCT$wnnzlizzieLet32_1_argbuf_rwb_r;
  Pointer_CT$wnnz_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Bool_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Bool_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Bool_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Int_Bool_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet20_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet22_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet14_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  MyDTInt_Int_Int_t wslR_2_2_argbuf_d;
  logic wslR_2_2_argbuf_r;
  MyDTInt_Int_Int_t wslR_2_1_d;
  logic wslR_2_1_r;
  MyDTInt_Int_Int_t wslR_2_2_d;
  logic wslR_2_2_r;
  MyDTInt_Int_Int_t wslR_3_2_argbuf_d;
  logic wslR_3_2_argbuf_r;
  MyDTInt_Int_Int_t wslR_3_1_d;
  logic wslR_3_1_r;
  MyDTInt_Int_Int_t wslR_3_2_d;
  logic wslR_3_2_r;
  MyDTInt_Int_Int_t wslR_4_1_argbuf_d;
  logic wslR_4_1_argbuf_r;
  Pointer_QTree_Bool_t wslW_1_1_argbuf_d;
  logic wslW_1_1_argbuf_r;
  CT$wnnz_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  CT$wnnz_t wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_d;
  logic wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_r;
  CT$wnnz_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  CT$wnnz_t wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_d;
  logic wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_r;
  \Int#_t  es_6_1ww2XmM_1_1_Add32_d;
  logic es_6_1ww2XmM_1_1_Add32_r;
  \Int#_t  wwslZ_3_1ww1XmJ_2_1_Add32_d;
  logic wwslZ_3_1ww1XmJ_2_1_Add32_r;
  MyBool_t xa88_1_argbuf_d;
  logic xa88_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(goFork,Go),
                                (goFor_2,Go),
                                (goFor_3,Go),
                                (goFor_4,Go),
                                (goFor_5,Go),
                                (goFor_6,Go),
                                (goFor_7,Go),
                                (goFor_8,Go),
                                (goFor_9,Go)] */
  logic [8:0] sourceGo_emitted;
  logic [8:0] sourceGo_done;
  assign goFork_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign goFor_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign goFor_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign goFor_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign goFor_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign goFor_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign goFor_7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign goFor_8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign goFor_9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign sourceGo_done = (sourceGo_emitted | ({goFor_9_d[0],
                                               goFor_8_d[0],
                                               goFor_7_d[0],
                                               goFor_6_d[0],
                                               goFor_5_d[0],
                                               goFor_4_d[0],
                                               goFor_3_d[0],
                                               goFor_2_d[0],
                                               goFork_d[0]} & {goFor_9_r,
                                                               goFor_8_r,
                                                               goFor_7_r,
                                                               goFor_6_r,
                                                               goFor_5_r,
                                                               goFor_4_r,
                                                               goFor_3_r,
                                                               goFor_2_r,
                                                               goFork_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 9'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 9'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_2,Go) > (initHP_CT$wmAdd_Int,Word16#) */
  assign initHP_CT$wmAdd_Int_d = {16'd0, goFor_2_d[0]};
  assign goFor_2_r = initHP_CT$wmAdd_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wmAdd_Int1,Go) > (incrHP_CT$wmAdd_Int,Word16#) */
  assign incrHP_CT$wmAdd_Int_d = {16'd1, incrHP_CT$wmAdd_Int1_d[0]};
  assign incrHP_CT$wmAdd_Int1_r = incrHP_CT$wmAdd_Int_r;
  
  /* merge (Ty Go) : [(goFor_3,Go),
                 (incrHP_CT$wmAdd_Int2,Go)] > (incrHP_mergeCT$wmAdd_Int,Go) */
  logic [1:0] incrHP_mergeCT$wmAdd_Int_selected;
  logic [1:0] incrHP_mergeCT$wmAdd_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wmAdd_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wmAdd_Int_select))
        incrHP_mergeCT$wmAdd_Int_selected = incrHP_mergeCT$wmAdd_Int_select;
      else
        if (goFor_3_d[0]) incrHP_mergeCT$wmAdd_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wmAdd_Int2_d[0])
          incrHP_mergeCT$wmAdd_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Int_select <= (incrHP_mergeCT$wmAdd_Int_r ? 2'd0 :
                                          incrHP_mergeCT$wmAdd_Int_selected);
  always_comb
    if (incrHP_mergeCT$wmAdd_Int_selected[0])
      incrHP_mergeCT$wmAdd_Int_d = goFor_3_d;
    else if (incrHP_mergeCT$wmAdd_Int_selected[1])
      incrHP_mergeCT$wmAdd_Int_d = incrHP_CT$wmAdd_Int2_d;
    else incrHP_mergeCT$wmAdd_Int_d = 1'd0;
  assign {incrHP_CT$wmAdd_Int2_r,
          goFor_3_r} = (incrHP_mergeCT$wmAdd_Int_r ? incrHP_mergeCT$wmAdd_Int_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wmAdd_Int_buf,Go) > [(incrHP_CT$wmAdd_Int1,Go),
                                                    (incrHP_CT$wmAdd_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wmAdd_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wmAdd_Int_buf_done;
  assign incrHP_CT$wmAdd_Int1_d = (incrHP_mergeCT$wmAdd_Int_buf_d[0] && (! incrHP_mergeCT$wmAdd_Int_buf_emitted[0]));
  assign incrHP_CT$wmAdd_Int2_d = (incrHP_mergeCT$wmAdd_Int_buf_d[0] && (! incrHP_mergeCT$wmAdd_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wmAdd_Int_buf_done = (incrHP_mergeCT$wmAdd_Int_buf_emitted | ({incrHP_CT$wmAdd_Int2_d[0],
                                                                                       incrHP_CT$wmAdd_Int1_d[0]} & {incrHP_CT$wmAdd_Int2_r,
                                                                                                                     incrHP_CT$wmAdd_Int1_r}));
  assign incrHP_mergeCT$wmAdd_Int_buf_r = (& incrHP_mergeCT$wmAdd_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Int_buf_emitted <= (incrHP_mergeCT$wmAdd_Int_buf_r ? 2'd0 :
                                               incrHP_mergeCT$wmAdd_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wmAdd_Int,Word16#) (forkHP1_CT$wmAdd_Int,Word16#) > (addHP_CT$wmAdd_Int,Word16#) */
  assign addHP_CT$wmAdd_Int_d = {(incrHP_CT$wmAdd_Int_d[16:1] + forkHP1_CT$wmAdd_Int_d[16:1]),
                                 (incrHP_CT$wmAdd_Int_d[0] && forkHP1_CT$wmAdd_Int_d[0])};
  assign {incrHP_CT$wmAdd_Int_r,
          forkHP1_CT$wmAdd_Int_r} = {2 {(addHP_CT$wmAdd_Int_r && addHP_CT$wmAdd_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wmAdd_Int,Word16#),
                      (addHP_CT$wmAdd_Int,Word16#)] > (mergeHP_CT$wmAdd_Int,Word16#) */
  logic [1:0] mergeHP_CT$wmAdd_Int_selected;
  logic [1:0] mergeHP_CT$wmAdd_Int_select;
  always_comb
    begin
      mergeHP_CT$wmAdd_Int_selected = 2'd0;
      if ((| mergeHP_CT$wmAdd_Int_select))
        mergeHP_CT$wmAdd_Int_selected = mergeHP_CT$wmAdd_Int_select;
      else
        if (initHP_CT$wmAdd_Int_d[0])
          mergeHP_CT$wmAdd_Int_selected[0] = 1'd1;
        else if (addHP_CT$wmAdd_Int_d[0])
          mergeHP_CT$wmAdd_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Int_select <= 2'd0;
    else
      mergeHP_CT$wmAdd_Int_select <= (mergeHP_CT$wmAdd_Int_r ? 2'd0 :
                                      mergeHP_CT$wmAdd_Int_selected);
  always_comb
    if (mergeHP_CT$wmAdd_Int_selected[0])
      mergeHP_CT$wmAdd_Int_d = initHP_CT$wmAdd_Int_d;
    else if (mergeHP_CT$wmAdd_Int_selected[1])
      mergeHP_CT$wmAdd_Int_d = addHP_CT$wmAdd_Int_d;
    else mergeHP_CT$wmAdd_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wmAdd_Int_r,
          initHP_CT$wmAdd_Int_r} = (mergeHP_CT$wmAdd_Int_r ? mergeHP_CT$wmAdd_Int_selected :
                                    2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wmAdd_Int,Go) > (incrHP_mergeCT$wmAdd_Int_buf,Go) */
  Go_t incrHP_mergeCT$wmAdd_Int_bufchan_d;
  logic incrHP_mergeCT$wmAdd_Int_bufchan_r;
  assign incrHP_mergeCT$wmAdd_Int_r = ((! incrHP_mergeCT$wmAdd_Int_bufchan_d[0]) || incrHP_mergeCT$wmAdd_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wmAdd_Int_r)
        incrHP_mergeCT$wmAdd_Int_bufchan_d <= incrHP_mergeCT$wmAdd_Int_d;
  Go_t incrHP_mergeCT$wmAdd_Int_bufchan_buf;
  assign incrHP_mergeCT$wmAdd_Int_bufchan_r = (! incrHP_mergeCT$wmAdd_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wmAdd_Int_buf_d = (incrHP_mergeCT$wmAdd_Int_bufchan_buf[0] ? incrHP_mergeCT$wmAdd_Int_bufchan_buf :
                                           incrHP_mergeCT$wmAdd_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wmAdd_Int_buf_r && incrHP_mergeCT$wmAdd_Int_bufchan_buf[0]))
        incrHP_mergeCT$wmAdd_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wmAdd_Int_buf_r) && (! incrHP_mergeCT$wmAdd_Int_bufchan_buf[0])))
        incrHP_mergeCT$wmAdd_Int_bufchan_buf <= incrHP_mergeCT$wmAdd_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wmAdd_Int,Word16#) > (mergeHP_CT$wmAdd_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wmAdd_Int_bufchan_d;
  logic mergeHP_CT$wmAdd_Int_bufchan_r;
  assign mergeHP_CT$wmAdd_Int_r = ((! mergeHP_CT$wmAdd_Int_bufchan_d[0]) || mergeHP_CT$wmAdd_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wmAdd_Int_r)
        mergeHP_CT$wmAdd_Int_bufchan_d <= mergeHP_CT$wmAdd_Int_d;
  \Word16#_t  mergeHP_CT$wmAdd_Int_bufchan_buf;
  assign mergeHP_CT$wmAdd_Int_bufchan_r = (! mergeHP_CT$wmAdd_Int_bufchan_buf[0]);
  assign mergeHP_CT$wmAdd_Int_buf_d = (mergeHP_CT$wmAdd_Int_bufchan_buf[0] ? mergeHP_CT$wmAdd_Int_bufchan_buf :
                                       mergeHP_CT$wmAdd_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wmAdd_Int_buf_r && mergeHP_CT$wmAdd_Int_bufchan_buf[0]))
        mergeHP_CT$wmAdd_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wmAdd_Int_buf_r) && (! mergeHP_CT$wmAdd_Int_bufchan_buf[0])))
        mergeHP_CT$wmAdd_Int_bufchan_buf <= mergeHP_CT$wmAdd_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wmAdd_Int_buf,Word16#) > [(forkHP1_CT$wmAdd_Int,Word16#),
                                                          (forkHP1_CT$wmAdd_In2,Word16#),
                                                          (forkHP1_CT$wmAdd_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wmAdd_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wmAdd_Int_buf_done;
  assign forkHP1_CT$wmAdd_Int_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[0]))};
  assign forkHP1_CT$wmAdd_In2_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[1]))};
  assign forkHP1_CT$wmAdd_In3_d = {mergeHP_CT$wmAdd_Int_buf_d[16:1],
                                   (mergeHP_CT$wmAdd_Int_buf_d[0] && (! mergeHP_CT$wmAdd_Int_buf_emitted[2]))};
  assign mergeHP_CT$wmAdd_Int_buf_done = (mergeHP_CT$wmAdd_Int_buf_emitted | ({forkHP1_CT$wmAdd_In3_d[0],
                                                                               forkHP1_CT$wmAdd_In2_d[0],
                                                                               forkHP1_CT$wmAdd_Int_d[0]} & {forkHP1_CT$wmAdd_In3_r,
                                                                                                             forkHP1_CT$wmAdd_In2_r,
                                                                                                             forkHP1_CT$wmAdd_Int_r}));
  assign mergeHP_CT$wmAdd_Int_buf_r = (& mergeHP_CT$wmAdd_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wmAdd_Int_buf_emitted <= (mergeHP_CT$wmAdd_Int_buf_r ? 3'd0 :
                                           mergeHP_CT$wmAdd_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wmAdd_Int) : [(dconReadIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int),
                                     (dconWriteIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int)] > (memMergeChoice_CT$wmAdd_Int,C2) (memMergeIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  logic [1:0] dconReadIn_CT$wmAdd_Int_select_d;
  assign dconReadIn_CT$wmAdd_Int_select_d = ((| dconReadIn_CT$wmAdd_Int_select_q) ? dconReadIn_CT$wmAdd_Int_select_q :
                                             (dconReadIn_CT$wmAdd_Int_d[0] ? 2'd1 :
                                              (dconWriteIn_CT$wmAdd_Int_d[0] ? 2'd2 :
                                               2'd0)));
  logic [1:0] dconReadIn_CT$wmAdd_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Int_select_q <= (dconReadIn_CT$wmAdd_Int_done ? 2'd0 :
                                           dconReadIn_CT$wmAdd_Int_select_d);
  logic [1:0] dconReadIn_CT$wmAdd_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Int_emit_q <= (dconReadIn_CT$wmAdd_Int_done ? 2'd0 :
                                         dconReadIn_CT$wmAdd_Int_emit_d);
  logic [1:0] dconReadIn_CT$wmAdd_Int_emit_d;
  assign dconReadIn_CT$wmAdd_Int_emit_d = (dconReadIn_CT$wmAdd_Int_emit_q | ({memMergeChoice_CT$wmAdd_Int_d[0],
                                                                              memMergeIn_CT$wmAdd_Int_d[0]} & {memMergeChoice_CT$wmAdd_Int_r,
                                                                                                               memMergeIn_CT$wmAdd_Int_r}));
  logic dconReadIn_CT$wmAdd_Int_done;
  assign dconReadIn_CT$wmAdd_Int_done = (& dconReadIn_CT$wmAdd_Int_emit_d);
  assign {dconWriteIn_CT$wmAdd_Int_r,
          dconReadIn_CT$wmAdd_Int_r} = (dconReadIn_CT$wmAdd_Int_done ? dconReadIn_CT$wmAdd_Int_select_d :
                                        2'd0);
  assign memMergeIn_CT$wmAdd_Int_d = ((dconReadIn_CT$wmAdd_Int_select_d[0] && (! dconReadIn_CT$wmAdd_Int_emit_q[0])) ? dconReadIn_CT$wmAdd_Int_d :
                                      ((dconReadIn_CT$wmAdd_Int_select_d[1] && (! dconReadIn_CT$wmAdd_Int_emit_q[0])) ? dconWriteIn_CT$wmAdd_Int_d :
                                       {132'd0, 1'd0}));
  assign memMergeChoice_CT$wmAdd_Int_d = ((dconReadIn_CT$wmAdd_Int_select_d[0] && (! dconReadIn_CT$wmAdd_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                          ((dconReadIn_CT$wmAdd_Int_select_d[1] && (! dconReadIn_CT$wmAdd_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                           {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wmAdd_Int,
      Ty MemOut_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int_dbuf,MemIn_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) */
  logic [114:0] memMergeIn_CT$wmAdd_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wmAdd_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wmAdd_Int_dbuf_din;
  logic [114:0] memOut_CT$wmAdd_Int_q;
  logic memOut_CT$wmAdd_Int_valid;
  logic memMergeIn_CT$wmAdd_Int_dbuf_we;
  logic memOut_CT$wmAdd_Int_we;
  assign memMergeIn_CT$wmAdd_Int_dbuf_din = memMergeIn_CT$wmAdd_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wmAdd_Int_dbuf_address = memMergeIn_CT$wmAdd_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wmAdd_Int_dbuf_we = (memMergeIn_CT$wmAdd_Int_dbuf_d[1:1] && memMergeIn_CT$wmAdd_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wmAdd_Int_we <= 1'd0;
        memOut_CT$wmAdd_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wmAdd_Int_we <= memMergeIn_CT$wmAdd_Int_dbuf_we;
        memOut_CT$wmAdd_Int_valid <= memMergeIn_CT$wmAdd_Int_dbuf_d[0];
        if (memMergeIn_CT$wmAdd_Int_dbuf_we)
          begin
            memMergeIn_CT$wmAdd_Int_dbuf_mem[memMergeIn_CT$wmAdd_Int_dbuf_address] <= memMergeIn_CT$wmAdd_Int_dbuf_din;
            memOut_CT$wmAdd_Int_q <= memMergeIn_CT$wmAdd_Int_dbuf_din;
          end
        else
          memOut_CT$wmAdd_Int_q <= memMergeIn_CT$wmAdd_Int_dbuf_mem[memMergeIn_CT$wmAdd_Int_dbuf_address];
      end
  assign memOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_q,
                                  memOut_CT$wmAdd_Int_we,
                                  memOut_CT$wmAdd_Int_valid};
  assign memMergeIn_CT$wmAdd_Int_dbuf_r = ((! memOut_CT$wmAdd_Int_valid) || memOut_CT$wmAdd_Int_r);
  logic [31:0] profiling_MemIn_CT$wmAdd_Int_read;
  logic [31:0] profiling_MemIn_CT$wmAdd_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wmAdd_Int_write <= 0;
        profiling_MemIn_CT$wmAdd_Int_read <= 0;
      end
    else
      if ((memMergeIn_CT$wmAdd_Int_dbuf_we == 1'd1))
        profiling_MemIn_CT$wmAdd_Int_write <= (profiling_MemIn_CT$wmAdd_Int_write + 1);
      else
        if ((memOut_CT$wmAdd_Int_valid == 1'd1))
          profiling_MemIn_CT$wmAdd_Int_read <= (profiling_MemIn_CT$wmAdd_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wmAdd_Int) : (memMergeChoice_CT$wmAdd_Int,C2) (memOut_CT$wmAdd_Int_dbuf,MemOut_CT$wmAdd_Int) > [(memReadOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int),
                                                                                                                    (memWriteOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int)] */
  logic [1:0] memOut_CT$wmAdd_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wmAdd_Int_d[0] && memOut_CT$wmAdd_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wmAdd_Int_d[1:1])
        1'd0: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wmAdd_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_dbuf_d[116:1],
                                      memOut_CT$wmAdd_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wmAdd_Int_d = {memOut_CT$wmAdd_Int_dbuf_d[116:1],
                                       memOut_CT$wmAdd_Int_dbuf_onehotd[1]};
  assign memOut_CT$wmAdd_Int_dbuf_r = (| (memOut_CT$wmAdd_Int_dbuf_onehotd & {memWriteOut_CT$wmAdd_Int_r,
                                                                              memReadOut_CT$wmAdd_Int_r}));
  assign memMergeChoice_CT$wmAdd_Int_r = memOut_CT$wmAdd_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int_rbuf,MemIn_CT$wmAdd_Int) > (memMergeIn_CT$wmAdd_Int_dbuf,MemIn_CT$wmAdd_Int) */
  assign memMergeIn_CT$wmAdd_Int_rbuf_r = ((! memMergeIn_CT$wmAdd_Int_dbuf_d[0]) || memMergeIn_CT$wmAdd_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wmAdd_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wmAdd_Int_rbuf_r)
        memMergeIn_CT$wmAdd_Int_dbuf_d <= memMergeIn_CT$wmAdd_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wmAdd_Int) : (memMergeIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) > (memMergeIn_CT$wmAdd_Int_rbuf,MemIn_CT$wmAdd_Int) */
  MemIn_CT$wmAdd_Int_t memMergeIn_CT$wmAdd_Int_buf;
  assign memMergeIn_CT$wmAdd_Int_r = (! memMergeIn_CT$wmAdd_Int_buf[0]);
  assign memMergeIn_CT$wmAdd_Int_rbuf_d = (memMergeIn_CT$wmAdd_Int_buf[0] ? memMergeIn_CT$wmAdd_Int_buf :
                                           memMergeIn_CT$wmAdd_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wmAdd_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wmAdd_Int_rbuf_r && memMergeIn_CT$wmAdd_Int_buf[0]))
        memMergeIn_CT$wmAdd_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wmAdd_Int_rbuf_r) && (! memMergeIn_CT$wmAdd_Int_buf[0])))
        memMergeIn_CT$wmAdd_Int_buf <= memMergeIn_CT$wmAdd_Int_d;
  
  /* dbuf (Ty MemOut_CT$wmAdd_Int) : (memOut_CT$wmAdd_Int_rbuf,MemOut_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int_dbuf,MemOut_CT$wmAdd_Int) */
  assign memOut_CT$wmAdd_Int_rbuf_r = ((! memOut_CT$wmAdd_Int_dbuf_d[0]) || memOut_CT$wmAdd_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wmAdd_Int_rbuf_r)
        memOut_CT$wmAdd_Int_dbuf_d <= memOut_CT$wmAdd_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wmAdd_Int) : (memOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) > (memOut_CT$wmAdd_Int_rbuf,MemOut_CT$wmAdd_Int) */
  MemOut_CT$wmAdd_Int_t memOut_CT$wmAdd_Int_buf;
  assign memOut_CT$wmAdd_Int_r = (! memOut_CT$wmAdd_Int_buf[0]);
  assign memOut_CT$wmAdd_Int_rbuf_d = (memOut_CT$wmAdd_Int_buf[0] ? memOut_CT$wmAdd_Int_buf :
                                       memOut_CT$wmAdd_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wmAdd_Int_rbuf_r && memOut_CT$wmAdd_Int_buf[0]))
        memOut_CT$wmAdd_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wmAdd_Int_rbuf_r) && (! memOut_CT$wmAdd_Int_buf[0])))
        memOut_CT$wmAdd_Int_buf <= memOut_CT$wmAdd_Int_d;
  
  /* destruct (Ty Pointer_CT$wmAdd_Int,
          Dcon Pointer_CT$wmAdd_Int) : (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Int) > [(destructReadIn_CT$wmAdd_Int,Word16#)] */
  assign destructReadIn_CT$wmAdd_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                          scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wmAdd_Int_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Int,
      Dcon ReadIn_CT$wmAdd_Int) : [(destructReadIn_CT$wmAdd_Int,Word16#)] > (dconReadIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  assign dconReadIn_CT$wmAdd_Int_d = ReadIn_CT$wmAdd_Int_dc((& {destructReadIn_CT$wmAdd_Int_d[0]}), destructReadIn_CT$wmAdd_Int_d);
  assign {destructReadIn_CT$wmAdd_Int_r} = {1 {(dconReadIn_CT$wmAdd_Int_r && dconReadIn_CT$wmAdd_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wmAdd_Int,
          Dcon ReadOut_CT$wmAdd_Int) : (memReadOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) > [(readPointer_CT$wmAdd_Intscfarg_0_1_argbuf,CT$wmAdd_Int)] */
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wmAdd_Int_d[116:2],
                                                        memReadOut_CT$wmAdd_Int_d[0]};
  assign memReadOut_CT$wmAdd_Int_r = readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wmAdd_Int) : [(lizzieLet0_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet12_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet25_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet26_1_argbuf,CT$wmAdd_Int),
                               (lizzieLet27_1_argbuf,CT$wmAdd_Int)] > (writeMerge_choice_CT$wmAdd_Int,C5) (writeMerge_data_CT$wmAdd_Int,CT$wmAdd_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet12_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet25_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet26_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet27_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wmAdd_Int_d[0],
                                                                      writeMerge_data_CT$wmAdd_Int_d[0]} & {writeMerge_choice_CT$wmAdd_Int_r,
                                                                                                            writeMerge_data_CT$wmAdd_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wmAdd_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet12_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                              ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                               {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wmAdd_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                 {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wmAdd_Int) : (writeMerge_choice_CT$wmAdd_Int,C5) (demuxWriteResult_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) > [(writeCT$wmAdd_IntlizzieLet0_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet12_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet25_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet26_1_argbuf,Pointer_CT$wmAdd_Int),
                                                                                                                              (writeCT$wmAdd_IntlizzieLet27_1_argbuf,Pointer_CT$wmAdd_Int)] */
  logic [4:0] demuxWriteResult_CT$wmAdd_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wmAdd_Int_d[0] && demuxWriteResult_CT$wmAdd_Int_d[0]))
      unique case (writeMerge_choice_CT$wmAdd_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wmAdd_Int_onehotd = 5'd0;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                   demuxWriteResult_CT$wmAdd_Int_onehotd[0]};
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[1]};
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[2]};
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[3]};
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Int_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Int_onehotd[4]};
  assign demuxWriteResult_CT$wmAdd_Int_r = (| (demuxWriteResult_CT$wmAdd_Int_onehotd & {writeCT$wmAdd_IntlizzieLet27_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet26_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet25_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet12_1_argbuf_r,
                                                                                        writeCT$wmAdd_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wmAdd_Int_r = demuxWriteResult_CT$wmAdd_Int_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Int,
      Dcon WriteIn_CT$wmAdd_Int) : [(forkHP1_CT$wmAdd_In2,Word16#),
                                    (writeMerge_data_CT$wmAdd_Int,CT$wmAdd_Int)] > (dconWriteIn_CT$wmAdd_Int,MemIn_CT$wmAdd_Int) */
  assign dconWriteIn_CT$wmAdd_Int_d = WriteIn_CT$wmAdd_Int_dc((& {forkHP1_CT$wmAdd_In2_d[0],
                                                                  writeMerge_data_CT$wmAdd_Int_d[0]}), forkHP1_CT$wmAdd_In2_d, writeMerge_data_CT$wmAdd_Int_d);
  assign {forkHP1_CT$wmAdd_In2_r,
          writeMerge_data_CT$wmAdd_Int_r} = {2 {(dconWriteIn_CT$wmAdd_Int_r && dconWriteIn_CT$wmAdd_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wmAdd_Int,
      Dcon Pointer_CT$wmAdd_Int) : [(forkHP1_CT$wmAdd_In3,Word16#)] > (dconPtr_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) */
  assign dconPtr_CT$wmAdd_Int_d = Pointer_CT$wmAdd_Int_dc((& {forkHP1_CT$wmAdd_In3_d[0]}), forkHP1_CT$wmAdd_In3_d);
  assign {forkHP1_CT$wmAdd_In3_r} = {1 {(dconPtr_CT$wmAdd_Int_r && dconPtr_CT$wmAdd_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wmAdd_Int,
       Ty Pointer_CT$wmAdd_Int) : (memWriteOut_CT$wmAdd_Int,MemOut_CT$wmAdd_Int) (dconPtr_CT$wmAdd_Int,Pointer_CT$wmAdd_Int) > [(_64,Pointer_CT$wmAdd_Int),
                                                                                                                                (demuxWriteResult_CT$wmAdd_Int,Pointer_CT$wmAdd_Int)] */
  logic [1:0] dconPtr_CT$wmAdd_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wmAdd_Int_d[0] && dconPtr_CT$wmAdd_Int_d[0]))
      unique case (memWriteOut_CT$wmAdd_Int_d[1:1])
        1'd0: dconPtr_CT$wmAdd_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wmAdd_Int_onehotd = 2'd2;
        default: dconPtr_CT$wmAdd_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wmAdd_Int_onehotd = 2'd0;
  assign _64_d = {dconPtr_CT$wmAdd_Int_d[16:1],
                  dconPtr_CT$wmAdd_Int_onehotd[0]};
  assign demuxWriteResult_CT$wmAdd_Int_d = {dconPtr_CT$wmAdd_Int_d[16:1],
                                            dconPtr_CT$wmAdd_Int_onehotd[1]};
  assign dconPtr_CT$wmAdd_Int_r = (| (dconPtr_CT$wmAdd_Int_onehotd & {demuxWriteResult_CT$wmAdd_Int_r,
                                                                      _64_r}));
  assign memWriteOut_CT$wmAdd_Int_r = dconPtr_CT$wmAdd_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Int) : [(ma8M_1_argbuf,Pointer_QTree_Int),
                                    (w1slS_1_1_argbuf,Pointer_QTree_Int),
                                    (w2slT_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C3) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [2:0] ma8M_1_argbuf_select_d;
  assign ma8M_1_argbuf_select_d = ((| ma8M_1_argbuf_select_q) ? ma8M_1_argbuf_select_q :
                                   (ma8M_1_argbuf_d[0] ? 3'd1 :
                                    (w1slS_1_1_argbuf_d[0] ? 3'd2 :
                                     (w2slT_1_1_argbuf_d[0] ? 3'd4 :
                                      3'd0))));
  logic [2:0] ma8M_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8M_1_argbuf_select_q <= 3'd0;
    else
      ma8M_1_argbuf_select_q <= (ma8M_1_argbuf_done ? 3'd0 :
                                 ma8M_1_argbuf_select_d);
  logic [1:0] ma8M_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8M_1_argbuf_emit_q <= 2'd0;
    else
      ma8M_1_argbuf_emit_q <= (ma8M_1_argbuf_done ? 2'd0 :
                               ma8M_1_argbuf_emit_d);
  logic [1:0] ma8M_1_argbuf_emit_d;
  assign ma8M_1_argbuf_emit_d = (ma8M_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                          readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                            readMerge_data_QTree_Int_r}));
  logic ma8M_1_argbuf_done;
  assign ma8M_1_argbuf_done = (& ma8M_1_argbuf_emit_d);
  assign {w2slT_1_1_argbuf_r,
          w1slS_1_1_argbuf_r,
          ma8M_1_argbuf_r} = (ma8M_1_argbuf_done ? ma8M_1_argbuf_select_d :
                              3'd0);
  assign readMerge_data_QTree_Int_d = ((ma8M_1_argbuf_select_d[0] && (! ma8M_1_argbuf_emit_q[0])) ? ma8M_1_argbuf_d :
                                       ((ma8M_1_argbuf_select_d[1] && (! ma8M_1_argbuf_emit_q[0])) ? w1slS_1_1_argbuf_d :
                                        ((ma8M_1_argbuf_select_d[2] && (! ma8M_1_argbuf_emit_q[0])) ? w2slT_1_1_argbuf_d :
                                         {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Int_d = ((ma8M_1_argbuf_select_d[0] && (! ma8M_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                         ((ma8M_1_argbuf_select_d[1] && (! ma8M_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                          ((ma8M_1_argbuf_select_d[2] && (! ma8M_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                           {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C3) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intma8M_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intw1slS_1_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intw2slT_1_1_argbuf,QTree_Int)] */
  logic [2:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 3'd4;
        default: destructReadOut_QTree_Int_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 3'd0;
  assign readPointer_QTree_Intma8M_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                 destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intw1slS_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                    destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_Intw2slT_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                    destructReadOut_QTree_Int_onehotd[2]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_Intw2slT_1_1_argbuf_r,
                                                                                readPointer_QTree_Intw1slS_1_1_argbuf_r,
                                                                                readPointer_QTree_Intma8M_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C8,
           Ty QTree_Int) : [(lizzieLet11_1_1_argbuf,QTree_Int),
                            (lizzieLet13_1_argbuf,QTree_Int),
                            (lizzieLet14_1_1_argbuf,QTree_Int),
                            (lizzieLet28_1_argbuf,QTree_Int),
                            (lizzieLet7_1_1_argbuf,QTree_Int),
                            (lizzieLet8_1_1_argbuf,QTree_Int),
                            (lizzieLet9_1_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C8) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [7:0] lizzieLet11_1_1_argbuf_select_d;
  assign lizzieLet11_1_1_argbuf_select_d = ((| lizzieLet11_1_1_argbuf_select_q) ? lizzieLet11_1_1_argbuf_select_q :
                                            (lizzieLet11_1_1_argbuf_d[0] ? 8'd1 :
                                             (lizzieLet13_1_argbuf_d[0] ? 8'd2 :
                                              (lizzieLet14_1_1_argbuf_d[0] ? 8'd4 :
                                               (lizzieLet28_1_argbuf_d[0] ? 8'd8 :
                                                (lizzieLet7_1_1_argbuf_d[0] ? 8'd16 :
                                                 (lizzieLet8_1_1_argbuf_d[0] ? 8'd32 :
                                                  (lizzieLet9_1_1_argbuf_d[0] ? 8'd64 :
                                                   (dummy_write_QTree_Int_d[0] ? 8'd128 :
                                                    8'd0)))))))));
  logic [7:0] lizzieLet11_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_select_q <= 8'd0;
    else
      lizzieLet11_1_1_argbuf_select_q <= (lizzieLet11_1_1_argbuf_done ? 8'd0 :
                                          lizzieLet11_1_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_1_argbuf_emit_q <= (lizzieLet11_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet11_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_d;
  assign lizzieLet11_1_1_argbuf_emit_d = (lizzieLet11_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                            writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                               writeMerge_data_QTree_Int_r}));
  logic lizzieLet11_1_1_argbuf_done;
  assign lizzieLet11_1_1_argbuf_done = (& lizzieLet11_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r,
          lizzieLet13_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r} = (lizzieLet11_1_1_argbuf_done ? lizzieLet11_1_1_argbuf_select_d :
                                       8'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                        ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_argbuf_d :
                                         ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet14_1_1_argbuf_d :
                                          ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                           ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_1_argbuf_d :
                                            ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet8_1_1_argbuf_d :
                                             ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_1_argbuf_d :
                                              ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                               {66'd0, 1'd0}))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C1_8_dc(1'd1) :
                                          ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C2_8_dc(1'd1) :
                                           ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C3_8_dc(1'd1) :
                                            ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C4_8_dc(1'd1) :
                                             ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C5_8_dc(1'd1) :
                                              ((lizzieLet11_1_1_argbuf_select_d[5] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C6_8_dc(1'd1) :
                                               ((lizzieLet11_1_1_argbuf_select_d[6] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C7_8_dc(1'd1) :
                                                ((lizzieLet11_1_1_argbuf_select_d[7] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C8_8_dc(1'd1) :
                                                 {3'd0, 1'd0}))))))));
  
  /* demux (Ty C8,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C8) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet14_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (writeQTree_IntlizzieLet9_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                  (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [7:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[3:1])
        3'd0: demuxWriteResult_QTree_Int_onehotd = 8'd1;
        3'd1: demuxWriteResult_QTree_Int_onehotd = 8'd2;
        3'd2: demuxWriteResult_QTree_Int_onehotd = 8'd4;
        3'd3: demuxWriteResult_QTree_Int_onehotd = 8'd8;
        3'd4: demuxWriteResult_QTree_Int_onehotd = 8'd16;
        3'd5: demuxWriteResult_QTree_Int_onehotd = 8'd32;
        3'd6: demuxWriteResult_QTree_Int_onehotd = 8'd64;
        3'd7: demuxWriteResult_QTree_Int_onehotd = 8'd128;
        default: demuxWriteResult_QTree_Int_onehotd = 8'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 8'd0;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet13_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet14_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet7_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                  demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet8_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                  demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet9_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                  demuxWriteResult_QTree_Int_onehotd[6]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[7]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet8_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet28_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet14_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet13_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet11_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_63,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _63_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _63_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,Lit 0) : (goFor_4,Go) > (initHP_CT$wnnz,Word16#) */
  assign initHP_CT$wnnz_d = {16'd0, goFor_4_d[0]};
  assign goFor_4_r = initHP_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz1,Go) > (incrHP_CT$wnnz,Word16#) */
  assign incrHP_CT$wnnz_d = {16'd1, incrHP_CT$wnnz1_d[0]};
  assign incrHP_CT$wnnz1_r = incrHP_CT$wnnz_r;
  
  /* merge (Ty Go) : [(goFor_5,Go),
                 (incrHP_CT$wnnz2,Go)] > (incrHP_mergeCT$wnnz,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_selected;
  logic [1:0] incrHP_mergeCT$wnnz_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_select))
        incrHP_mergeCT$wnnz_selected = incrHP_mergeCT$wnnz_select;
      else
        if (goFor_5_d[0]) incrHP_mergeCT$wnnz_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz2_d[0])
          incrHP_mergeCT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_select <= (incrHP_mergeCT$wnnz_r ? 2'd0 :
                                     incrHP_mergeCT$wnnz_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_selected[0])
      incrHP_mergeCT$wnnz_d = goFor_5_d;
    else if (incrHP_mergeCT$wnnz_selected[1])
      incrHP_mergeCT$wnnz_d = incrHP_CT$wnnz2_d;
    else incrHP_mergeCT$wnnz_d = 1'd0;
  assign {incrHP_CT$wnnz2_r,
          goFor_5_r} = (incrHP_mergeCT$wnnz_r ? incrHP_mergeCT$wnnz_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_buf,Go) > [(incrHP_CT$wnnz1,Go),
                                               (incrHP_CT$wnnz2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_buf_done;
  assign incrHP_CT$wnnz1_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[0]));
  assign incrHP_CT$wnnz2_d = (incrHP_mergeCT$wnnz_buf_d[0] && (! incrHP_mergeCT$wnnz_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_buf_done = (incrHP_mergeCT$wnnz_buf_emitted | ({incrHP_CT$wnnz2_d[0],
                                                                             incrHP_CT$wnnz1_d[0]} & {incrHP_CT$wnnz2_r,
                                                                                                      incrHP_CT$wnnz1_r}));
  assign incrHP_mergeCT$wnnz_buf_r = (& incrHP_mergeCT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_buf_emitted <= (incrHP_mergeCT$wnnz_buf_r ? 2'd0 :
                                          incrHP_mergeCT$wnnz_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz,Word16#) (forkHP1_CT$wnnz,Word16#) > (addHP_CT$wnnz,Word16#) */
  assign addHP_CT$wnnz_d = {(incrHP_CT$wnnz_d[16:1] + forkHP1_CT$wnnz_d[16:1]),
                            (incrHP_CT$wnnz_d[0] && forkHP1_CT$wnnz_d[0])};
  assign {incrHP_CT$wnnz_r,
          forkHP1_CT$wnnz_r} = {2 {(addHP_CT$wnnz_r && addHP_CT$wnnz_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz,Word16#),
                      (addHP_CT$wnnz,Word16#)] > (mergeHP_CT$wnnz,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_selected;
  logic [1:0] mergeHP_CT$wnnz_select;
  always_comb
    begin
      mergeHP_CT$wnnz_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_select))
        mergeHP_CT$wnnz_selected = mergeHP_CT$wnnz_select;
      else
        if (initHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_d[0]) mergeHP_CT$wnnz_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_select <= 2'd0;
    else
      mergeHP_CT$wnnz_select <= (mergeHP_CT$wnnz_r ? 2'd0 :
                                 mergeHP_CT$wnnz_selected);
  always_comb
    if (mergeHP_CT$wnnz_selected[0])
      mergeHP_CT$wnnz_d = initHP_CT$wnnz_d;
    else if (mergeHP_CT$wnnz_selected[1])
      mergeHP_CT$wnnz_d = addHP_CT$wnnz_d;
    else mergeHP_CT$wnnz_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_r,
          initHP_CT$wnnz_r} = (mergeHP_CT$wnnz_r ? mergeHP_CT$wnnz_selected :
                               2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz,Go) > (incrHP_mergeCT$wnnz_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_bufchan_d;
  logic incrHP_mergeCT$wnnz_bufchan_r;
  assign incrHP_mergeCT$wnnz_r = ((! incrHP_mergeCT$wnnz_bufchan_d[0]) || incrHP_mergeCT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_r)
        incrHP_mergeCT$wnnz_bufchan_d <= incrHP_mergeCT$wnnz_d;
  Go_t incrHP_mergeCT$wnnz_bufchan_buf;
  assign incrHP_mergeCT$wnnz_bufchan_r = (! incrHP_mergeCT$wnnz_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_buf_d = (incrHP_mergeCT$wnnz_bufchan_buf[0] ? incrHP_mergeCT$wnnz_bufchan_buf :
                                      incrHP_mergeCT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_buf_r && incrHP_mergeCT$wnnz_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_buf_r) && (! incrHP_mergeCT$wnnz_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_bufchan_buf <= incrHP_mergeCT$wnnz_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz,Word16#) > (mergeHP_CT$wnnz_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_bufchan_d;
  logic mergeHP_CT$wnnz_bufchan_r;
  assign mergeHP_CT$wnnz_r = ((! mergeHP_CT$wnnz_bufchan_d[0]) || mergeHP_CT$wnnz_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_r)
        mergeHP_CT$wnnz_bufchan_d <= mergeHP_CT$wnnz_d;
  \Word16#_t  mergeHP_CT$wnnz_bufchan_buf;
  assign mergeHP_CT$wnnz_bufchan_r = (! mergeHP_CT$wnnz_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_buf_d = (mergeHP_CT$wnnz_bufchan_buf[0] ? mergeHP_CT$wnnz_bufchan_buf :
                                  mergeHP_CT$wnnz_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_buf_r && mergeHP_CT$wnnz_bufchan_buf[0]))
        mergeHP_CT$wnnz_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_buf_r) && (! mergeHP_CT$wnnz_bufchan_buf[0])))
        mergeHP_CT$wnnz_bufchan_buf <= mergeHP_CT$wnnz_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_buf,Word16#) > [(forkHP1_CT$wnnz,Word16#),
                                                     (forkHP1_CT$wnn2,Word16#),
                                                     (forkHP1_CT$wnn3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_buf_done;
  assign forkHP1_CT$wnnz_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[0]))};
  assign forkHP1_CT$wnn2_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[1]))};
  assign forkHP1_CT$wnn3_d = {mergeHP_CT$wnnz_buf_d[16:1],
                              (mergeHP_CT$wnnz_buf_d[0] && (! mergeHP_CT$wnnz_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_buf_done = (mergeHP_CT$wnnz_buf_emitted | ({forkHP1_CT$wnn3_d[0],
                                                                     forkHP1_CT$wnn2_d[0],
                                                                     forkHP1_CT$wnnz_d[0]} & {forkHP1_CT$wnn3_r,
                                                                                              forkHP1_CT$wnn2_r,
                                                                                              forkHP1_CT$wnnz_r}));
  assign mergeHP_CT$wnnz_buf_r = (& mergeHP_CT$wnnz_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_buf_emitted <= (mergeHP_CT$wnnz_buf_r ? 3'd0 :
                                      mergeHP_CT$wnnz_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz) : [(dconReadIn_CT$wnnz,MemIn_CT$wnnz),
                                (dconWriteIn_CT$wnnz,MemIn_CT$wnnz)] > (memMergeChoice_CT$wnnz,C2) (memMergeIn_CT$wnnz,MemIn_CT$wnnz) */
  logic [1:0] dconReadIn_CT$wnnz_select_d;
  assign dconReadIn_CT$wnnz_select_d = ((| dconReadIn_CT$wnnz_select_q) ? dconReadIn_CT$wnnz_select_q :
                                        (dconReadIn_CT$wnnz_d[0] ? 2'd1 :
                                         (dconWriteIn_CT$wnnz_d[0] ? 2'd2 :
                                          2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_select_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                      dconReadIn_CT$wnnz_select_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_emit_q <= (dconReadIn_CT$wnnz_done ? 2'd0 :
                                    dconReadIn_CT$wnnz_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_emit_d;
  assign dconReadIn_CT$wnnz_emit_d = (dconReadIn_CT$wnnz_emit_q | ({memMergeChoice_CT$wnnz_d[0],
                                                                    memMergeIn_CT$wnnz_d[0]} & {memMergeChoice_CT$wnnz_r,
                                                                                                memMergeIn_CT$wnnz_r}));
  logic dconReadIn_CT$wnnz_done;
  assign dconReadIn_CT$wnnz_done = (& dconReadIn_CT$wnnz_emit_d);
  assign {dconWriteIn_CT$wnnz_r,
          dconReadIn_CT$wnnz_r} = (dconReadIn_CT$wnnz_done ? dconReadIn_CT$wnnz_select_d :
                                   2'd0);
  assign memMergeIn_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconReadIn_CT$wnnz_d :
                                 ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[0])) ? dconWriteIn_CT$wnnz_d :
                                  {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_d = ((dconReadIn_CT$wnnz_select_d[0] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C1_2_dc(1'd1) :
                                     ((dconReadIn_CT$wnnz_select_d[1] && (! dconReadIn_CT$wnnz_emit_q[1])) ? C2_2_dc(1'd1) :
                                      {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz,
      Ty MemOut_CT$wnnz) : (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) > (memOut_CT$wnnz,MemOut_CT$wnnz) */
  logic [114:0] memMergeIn_CT$wnnz_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_dbuf_din;
  logic [114:0] memOut_CT$wnnz_q;
  logic memOut_CT$wnnz_valid;
  logic memMergeIn_CT$wnnz_dbuf_we;
  logic memOut_CT$wnnz_we;
  assign memMergeIn_CT$wnnz_dbuf_din = memMergeIn_CT$wnnz_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_dbuf_address = memMergeIn_CT$wnnz_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_dbuf_we = (memMergeIn_CT$wnnz_dbuf_d[1:1] && memMergeIn_CT$wnnz_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_we <= 1'd0;
        memOut_CT$wnnz_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_we <= memMergeIn_CT$wnnz_dbuf_we;
        memOut_CT$wnnz_valid <= memMergeIn_CT$wnnz_dbuf_d[0];
        if (memMergeIn_CT$wnnz_dbuf_we)
          begin
            memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address] <= memMergeIn_CT$wnnz_dbuf_din;
            memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_din;
          end
        else
          memOut_CT$wnnz_q <= memMergeIn_CT$wnnz_dbuf_mem[memMergeIn_CT$wnnz_dbuf_address];
      end
  assign memOut_CT$wnnz_d = {memOut_CT$wnnz_q,
                             memOut_CT$wnnz_we,
                             memOut_CT$wnnz_valid};
  assign memMergeIn_CT$wnnz_dbuf_r = ((! memOut_CT$wnnz_valid) || memOut_CT$wnnz_r);
  logic [31:0] profiling_MemIn_CT$wnnz_read;
  logic [31:0] profiling_MemIn_CT$wnnz_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_write <= 0;
        profiling_MemIn_CT$wnnz_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_write <= (profiling_MemIn_CT$wnnz_write + 1);
      else
        if ((memOut_CT$wnnz_valid == 1'd1))
          profiling_MemIn_CT$wnnz_read <= (profiling_MemIn_CT$wnnz_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz) : (memMergeChoice_CT$wnnz,C2) (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) > [(memReadOut_CT$wnnz,MemOut_CT$wnnz),
                                                                                                (memWriteOut_CT$wnnz,MemOut_CT$wnnz)] */
  logic [1:0] memOut_CT$wnnz_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_d[0] && memOut_CT$wnnz_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_d[1:1])
        1'd0: memOut_CT$wnnz_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                 memOut_CT$wnnz_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_d = {memOut_CT$wnnz_dbuf_d[116:1],
                                  memOut_CT$wnnz_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_dbuf_r = (| (memOut_CT$wnnz_dbuf_onehotd & {memWriteOut_CT$wnnz_r,
                                                                    memReadOut_CT$wnnz_r}));
  assign memMergeChoice_CT$wnnz_r = memOut_CT$wnnz_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_dbuf,MemIn_CT$wnnz) */
  assign memMergeIn_CT$wnnz_rbuf_r = ((! memMergeIn_CT$wnnz_dbuf_d[0]) || memMergeIn_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_rbuf_r)
        memMergeIn_CT$wnnz_dbuf_d <= memMergeIn_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz) : (memMergeIn_CT$wnnz,MemIn_CT$wnnz) > (memMergeIn_CT$wnnz_rbuf,MemIn_CT$wnnz) */
  MemIn_CT$wnnz_t memMergeIn_CT$wnnz_buf;
  assign memMergeIn_CT$wnnz_r = (! memMergeIn_CT$wnnz_buf[0]);
  assign memMergeIn_CT$wnnz_rbuf_d = (memMergeIn_CT$wnnz_buf[0] ? memMergeIn_CT$wnnz_buf :
                                      memMergeIn_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_rbuf_r && memMergeIn_CT$wnnz_buf[0]))
        memMergeIn_CT$wnnz_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_rbuf_r) && (! memMergeIn_CT$wnnz_buf[0])))
        memMergeIn_CT$wnnz_buf <= memMergeIn_CT$wnnz_d;
  
  /* dbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) > (memOut_CT$wnnz_dbuf,MemOut_CT$wnnz) */
  assign memOut_CT$wnnz_rbuf_r = ((! memOut_CT$wnnz_dbuf_d[0]) || memOut_CT$wnnz_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_rbuf_r)
        memOut_CT$wnnz_dbuf_d <= memOut_CT$wnnz_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz) : (memOut_CT$wnnz,MemOut_CT$wnnz) > (memOut_CT$wnnz_rbuf,MemOut_CT$wnnz) */
  MemOut_CT$wnnz_t memOut_CT$wnnz_buf;
  assign memOut_CT$wnnz_r = (! memOut_CT$wnnz_buf[0]);
  assign memOut_CT$wnnz_rbuf_d = (memOut_CT$wnnz_buf[0] ? memOut_CT$wnnz_buf :
                                  memOut_CT$wnnz_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_rbuf_r && memOut_CT$wnnz_buf[0]))
        memOut_CT$wnnz_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_rbuf_r) && (! memOut_CT$wnnz_buf[0])))
        memOut_CT$wnnz_buf <= memOut_CT$wnnz_d;
  
  /* destruct (Ty Pointer_CT$wnnz,
          Dcon Pointer_CT$wnnz) : (scfarg_0_1_1_argbuf,Pointer_CT$wnnz) > [(destructReadIn_CT$wnnz,Word16#)] */
  assign destructReadIn_CT$wnnz_d = {scfarg_0_1_1_argbuf_d[16:1],
                                     scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon ReadIn_CT$wnnz) : [(destructReadIn_CT$wnnz,Word16#)] > (dconReadIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconReadIn_CT$wnnz_d = ReadIn_CT$wnnz_dc((& {destructReadIn_CT$wnnz_d[0]}), destructReadIn_CT$wnnz_d);
  assign {destructReadIn_CT$wnnz_r} = {1 {(dconReadIn_CT$wnnz_r && dconReadIn_CT$wnnz_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz,
          Dcon ReadOut_CT$wnnz) : (memReadOut_CT$wnnz,MemOut_CT$wnnz) > [(readPointer_CT$wnnzscfarg_0_1_1_argbuf,CT$wnnz)] */
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_d = {memReadOut_CT$wnnz_d[116:2],
                                                     memReadOut_CT$wnnz_d[0]};
  assign memReadOut_CT$wnnz_r = readPointer_CT$wnnzscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,Ty CT$wnnz) : [(lizzieLet16_1_argbuf,CT$wnnz),
                                (lizzieLet1_1_argbuf,CT$wnnz),
                                (lizzieLet30_1_argbuf,CT$wnnz),
                                (lizzieLet31_1_argbuf,CT$wnnz),
                                (lizzieLet32_1_argbuf,CT$wnnz)] > (writeMerge_choice_CT$wnnz,C5) (writeMerge_data_CT$wnnz,CT$wnnz) */
  logic [4:0] lizzieLet16_1_argbuf_select_d;
  assign lizzieLet16_1_argbuf_select_d = ((| lizzieLet16_1_argbuf_select_q) ? lizzieLet16_1_argbuf_select_q :
                                          (lizzieLet16_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet1_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet30_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet31_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet32_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet16_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet16_1_argbuf_select_q <= (lizzieLet16_1_argbuf_done ? 5'd0 :
                                        lizzieLet16_1_argbuf_select_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet16_1_argbuf_emit_q <= (lizzieLet16_1_argbuf_done ? 2'd0 :
                                      lizzieLet16_1_argbuf_emit_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_d;
  assign lizzieLet16_1_argbuf_emit_d = (lizzieLet16_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_d[0],
                                                                        writeMerge_data_CT$wnnz_d[0]} & {writeMerge_choice_CT$wnnz_r,
                                                                                                         writeMerge_data_CT$wnnz_r}));
  logic lizzieLet16_1_argbuf_done;
  assign lizzieLet16_1_argbuf_done = (& lizzieLet16_1_argbuf_emit_d);
  assign {lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet1_1_argbuf_r,
          lizzieLet16_1_argbuf_r} = (lizzieLet16_1_argbuf_done ? lizzieLet16_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CT$wnnz_d = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                      ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet1_1_argbuf_d :
                                       ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                        ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                         ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                          {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_d = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                        ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                         ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                          ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                           ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                            {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz) : (writeMerge_choice_CT$wnnz,C5) (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz) > [(writeCT$wnnzlizzieLet16_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet1_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet30_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet31_1_argbuf,Pointer_CT$wnnz),
                                                                                                          (writeCT$wnnzlizzieLet32_1_argbuf,Pointer_CT$wnnz)] */
  logic [4:0] demuxWriteResult_CT$wnnz_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_d[0] && demuxWriteResult_CT$wnnz_d[0]))
      unique case (writeMerge_choice_CT$wnnz_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_onehotd = 5'd0;
  assign writeCT$wnnzlizzieLet16_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[0]};
  assign writeCT$wnnzlizzieLet1_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                              demuxWriteResult_CT$wnnz_onehotd[1]};
  assign writeCT$wnnzlizzieLet30_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[2]};
  assign writeCT$wnnzlizzieLet31_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[3]};
  assign writeCT$wnnzlizzieLet32_1_argbuf_d = {demuxWriteResult_CT$wnnz_d[16:1],
                                               demuxWriteResult_CT$wnnz_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_r = (| (demuxWriteResult_CT$wnnz_onehotd & {writeCT$wnnzlizzieLet32_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet31_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet30_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet1_1_argbuf_r,
                                                                              writeCT$wnnzlizzieLet16_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_r = demuxWriteResult_CT$wnnz_r;
  
  /* dcon (Ty MemIn_CT$wnnz,
      Dcon WriteIn_CT$wnnz) : [(forkHP1_CT$wnn2,Word16#),
                               (writeMerge_data_CT$wnnz,CT$wnnz)] > (dconWriteIn_CT$wnnz,MemIn_CT$wnnz) */
  assign dconWriteIn_CT$wnnz_d = WriteIn_CT$wnnz_dc((& {forkHP1_CT$wnn2_d[0],
                                                        writeMerge_data_CT$wnnz_d[0]}), forkHP1_CT$wnn2_d, writeMerge_data_CT$wnnz_d);
  assign {forkHP1_CT$wnn2_r,
          writeMerge_data_CT$wnnz_r} = {2 {(dconWriteIn_CT$wnnz_r && dconWriteIn_CT$wnnz_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz,
      Dcon Pointer_CT$wnnz) : [(forkHP1_CT$wnn3,Word16#)] > (dconPtr_CT$wnnz,Pointer_CT$wnnz) */
  assign dconPtr_CT$wnnz_d = Pointer_CT$wnnz_dc((& {forkHP1_CT$wnn3_d[0]}), forkHP1_CT$wnn3_d);
  assign {forkHP1_CT$wnn3_r} = {1 {(dconPtr_CT$wnnz_r && dconPtr_CT$wnnz_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz,
       Ty Pointer_CT$wnnz) : (memWriteOut_CT$wnnz,MemOut_CT$wnnz) (dconPtr_CT$wnnz,Pointer_CT$wnnz) > [(_62,Pointer_CT$wnnz),
                                                                                                       (demuxWriteResult_CT$wnnz,Pointer_CT$wnnz)] */
  logic [1:0] dconPtr_CT$wnnz_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_d[0] && dconPtr_CT$wnnz_d[0]))
      unique case (memWriteOut_CT$wnnz_d[1:1])
        1'd0: dconPtr_CT$wnnz_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_onehotd = 2'd0;
  assign _62_d = {dconPtr_CT$wnnz_d[16:1],
                  dconPtr_CT$wnnz_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_d = {dconPtr_CT$wnnz_d[16:1],
                                       dconPtr_CT$wnnz_onehotd[1]};
  assign dconPtr_CT$wnnz_r = (| (dconPtr_CT$wnnz_onehotd & {demuxWriteResult_CT$wnnz_r,
                                                            _62_r}));
  assign memWriteOut_CT$wnnz_r = dconPtr_CT$wnnz_r;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_6,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0, goFor_6_d[0]};
  assign goFor_6_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(goFor_7,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (goFor_7_d[0]) incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = goFor_7_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          goFor_7_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Boo2,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#)] */
  logic [2:0] mergeHP_QTree_Bool_buf_emitted;
  logic [2:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Boo2_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Boo2_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Boo2_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 3'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (wslW_1_1_argbuf,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {wslW_1_1_argbuf_d[16:1],
                                        wslW_1_1_argbuf_d[0]};
  assign wslW_1_1_argbuf_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(readPointer_QTree_BoolwslW_1_1_argbuf,QTree_Bool)] */
  assign readPointer_QTree_BoolwslW_1_1_argbuf_d = {memReadOut_QTree_Bool_d[67:2],
                                                    memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = readPointer_QTree_BoolwslW_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty QTree_Bool) : [(lizzieLet18_1_argbuf,QTree_Bool),
                             (lizzieLet19_1_argbuf,QTree_Bool),
                             (lizzieLet20_1_argbuf,QTree_Bool),
                             (lizzieLet22_1_argbuf,QTree_Bool),
                             (lizzieLet37_1_argbuf,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C5) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [4:0] lizzieLet18_1_argbuf_select_d;
  assign lizzieLet18_1_argbuf_select_d = ((| lizzieLet18_1_argbuf_select_q) ? lizzieLet18_1_argbuf_select_q :
                                          (lizzieLet18_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet19_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet20_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet22_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet37_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet18_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet18_1_argbuf_select_q <= (lizzieLet18_1_argbuf_done ? 5'd0 :
                                        lizzieLet18_1_argbuf_select_d);
  logic [1:0] lizzieLet18_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet18_1_argbuf_emit_q <= (lizzieLet18_1_argbuf_done ? 2'd0 :
                                      lizzieLet18_1_argbuf_emit_d);
  logic [1:0] lizzieLet18_1_argbuf_emit_d;
  assign lizzieLet18_1_argbuf_emit_d = (lizzieLet18_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                        writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                            writeMerge_data_QTree_Bool_r}));
  logic lizzieLet18_1_argbuf_done;
  assign lizzieLet18_1_argbuf_done = (& lizzieLet18_1_argbuf_emit_d);
  assign {lizzieLet37_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet19_1_argbuf_r,
          lizzieLet18_1_argbuf_r} = (lizzieLet18_1_argbuf_done ? lizzieLet18_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet18_1_argbuf_select_d[0] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                         ((lizzieLet18_1_argbuf_select_d[1] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet19_1_argbuf_d :
                                          ((lizzieLet18_1_argbuf_select_d[2] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                           ((lizzieLet18_1_argbuf_select_d[3] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                            ((lizzieLet18_1_argbuf_select_d[4] && (! lizzieLet18_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                             {66'd0, 1'd0})))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet18_1_argbuf_select_d[0] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                           ((lizzieLet18_1_argbuf_select_d[1] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                            ((lizzieLet18_1_argbuf_select_d[2] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                             ((lizzieLet18_1_argbuf_select_d[3] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                              ((lizzieLet18_1_argbuf_select_d[4] && (! lizzieLet18_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                               {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C5) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet18_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet19_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet20_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet22_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool)] */
  logic [4:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[3:1])
        3'd0: demuxWriteResult_QTree_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_QTree_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_QTree_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_QTree_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_QTree_Bool_onehotd = 5'd16;
        default: demuxWriteResult_QTree_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 5'd0;
  assign writeQTree_BoollizzieLet18_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet19_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet20_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet22_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet37_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {writeQTree_BoollizzieLet37_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet22_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet20_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet19_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet18_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo2,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo2_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo2_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo2_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0]}), forkHP1_QTree_Boo3_d);
  assign {forkHP1_QTree_Boo3_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_61,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _61_d = {dconPtr_QTree_Bool_d[16:1],
                  dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _61_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (goFor_8,Go) > (initHP_CTmain_map'_Int_Bool,Word16#) */
  assign \initHP_CTmain_map'_Int_Bool_d  = {16'd0, goFor_8_d[0]};
  assign goFor_8_r = \initHP_CTmain_map'_Int_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_map'_Int_Bool1,Go) > (incrHP_CTmain_map'_Int_Bool,Word16#) */
  assign \incrHP_CTmain_map'_Int_Bool_d  = {16'd1,
                                            \incrHP_CTmain_map'_Int_Bool1_d [0]};
  assign \incrHP_CTmain_map'_Int_Bool1_r  = \incrHP_CTmain_map'_Int_Bool_r ;
  
  /* merge (Ty Go) : [(goFor_9,Go),
                 (incrHP_CTmain_map'_Int_Bool2,Go)] > (incrHP_mergeCTmain_map'_Int_Bool,Go) */
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Bool_selected ;
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Bool_select ;
  always_comb
    begin
      \incrHP_mergeCTmain_map'_Int_Bool_selected  = 2'd0;
      if ((| \incrHP_mergeCTmain_map'_Int_Bool_select ))
        \incrHP_mergeCTmain_map'_Int_Bool_selected  = \incrHP_mergeCTmain_map'_Int_Bool_select ;
      else
        if (goFor_9_d[0])
          \incrHP_mergeCTmain_map'_Int_Bool_selected [0] = 1'd1;
        else if (\incrHP_CTmain_map'_Int_Bool2_d [0])
          \incrHP_mergeCTmain_map'_Int_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Bool_select  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Int_Bool_select  <= (\incrHP_mergeCTmain_map'_Int_Bool_r  ? 2'd0 :
                                                    \incrHP_mergeCTmain_map'_Int_Bool_selected );
  always_comb
    if (\incrHP_mergeCTmain_map'_Int_Bool_selected [0])
      \incrHP_mergeCTmain_map'_Int_Bool_d  = goFor_9_d;
    else if (\incrHP_mergeCTmain_map'_Int_Bool_selected [1])
      \incrHP_mergeCTmain_map'_Int_Bool_d  = \incrHP_CTmain_map'_Int_Bool2_d ;
    else \incrHP_mergeCTmain_map'_Int_Bool_d  = 1'd0;
  assign {\incrHP_CTmain_map'_Int_Bool2_r ,
          goFor_9_r} = (\incrHP_mergeCTmain_map'_Int_Bool_r  ? \incrHP_mergeCTmain_map'_Int_Bool_selected  :
                        2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_map'_Int_Bool_buf,Go) > [(incrHP_CTmain_map'_Int_Bool1,Go),
                                                            (incrHP_CTmain_map'_Int_Bool2,Go)] */
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Bool_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmain_map'_Int_Bool_buf_done ;
  assign \incrHP_CTmain_map'_Int_Bool1_d  = (\incrHP_mergeCTmain_map'_Int_Bool_buf_d [0] && (! \incrHP_mergeCTmain_map'_Int_Bool_buf_emitted [0]));
  assign \incrHP_CTmain_map'_Int_Bool2_d  = (\incrHP_mergeCTmain_map'_Int_Bool_buf_d [0] && (! \incrHP_mergeCTmain_map'_Int_Bool_buf_emitted [1]));
  assign \incrHP_mergeCTmain_map'_Int_Bool_buf_done  = (\incrHP_mergeCTmain_map'_Int_Bool_buf_emitted  | ({\incrHP_CTmain_map'_Int_Bool2_d [0],
                                                                                                           \incrHP_CTmain_map'_Int_Bool1_d [0]} & {\incrHP_CTmain_map'_Int_Bool2_r ,
                                                                                                                                                   \incrHP_CTmain_map'_Int_Bool1_r }));
  assign \incrHP_mergeCTmain_map'_Int_Bool_buf_r  = (& \incrHP_mergeCTmain_map'_Int_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Bool_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Int_Bool_buf_emitted  <= (\incrHP_mergeCTmain_map'_Int_Bool_buf_r  ? 2'd0 :
                                                         \incrHP_mergeCTmain_map'_Int_Bool_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_map'_Int_Bool,Word16#) (forkHP1_CTmain_map'_Int_Bool,Word16#) > (addHP_CTmain_map'_Int_Bool,Word16#) */
  assign \addHP_CTmain_map'_Int_Bool_d  = {(\incrHP_CTmain_map'_Int_Bool_d [16:1] + \forkHP1_CTmain_map'_Int_Bool_d [16:1]),
                                           (\incrHP_CTmain_map'_Int_Bool_d [0] && \forkHP1_CTmain_map'_Int_Bool_d [0])};
  assign {\incrHP_CTmain_map'_Int_Bool_r ,
          \forkHP1_CTmain_map'_Int_Bool_r } = {2 {(\addHP_CTmain_map'_Int_Bool_r  && \addHP_CTmain_map'_Int_Bool_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_map'_Int_Bool,Word16#),
                      (addHP_CTmain_map'_Int_Bool,Word16#)] > (mergeHP_CTmain_map'_Int_Bool,Word16#) */
  logic [1:0] \mergeHP_CTmain_map'_Int_Bool_selected ;
  logic [1:0] \mergeHP_CTmain_map'_Int_Bool_select ;
  always_comb
    begin
      \mergeHP_CTmain_map'_Int_Bool_selected  = 2'd0;
      if ((| \mergeHP_CTmain_map'_Int_Bool_select ))
        \mergeHP_CTmain_map'_Int_Bool_selected  = \mergeHP_CTmain_map'_Int_Bool_select ;
      else
        if (\initHP_CTmain_map'_Int_Bool_d [0])
          \mergeHP_CTmain_map'_Int_Bool_selected [0] = 1'd1;
        else if (\addHP_CTmain_map'_Int_Bool_d [0])
          \mergeHP_CTmain_map'_Int_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTmain_map'_Int_Bool_select  <= 2'd0;
    else
      \mergeHP_CTmain_map'_Int_Bool_select  <= (\mergeHP_CTmain_map'_Int_Bool_r  ? 2'd0 :
                                                \mergeHP_CTmain_map'_Int_Bool_selected );
  always_comb
    if (\mergeHP_CTmain_map'_Int_Bool_selected [0])
      \mergeHP_CTmain_map'_Int_Bool_d  = \initHP_CTmain_map'_Int_Bool_d ;
    else if (\mergeHP_CTmain_map'_Int_Bool_selected [1])
      \mergeHP_CTmain_map'_Int_Bool_d  = \addHP_CTmain_map'_Int_Bool_d ;
    else \mergeHP_CTmain_map'_Int_Bool_d  = {16'd0, 1'd0};
  assign {\addHP_CTmain_map'_Int_Bool_r ,
          \initHP_CTmain_map'_Int_Bool_r } = (\mergeHP_CTmain_map'_Int_Bool_r  ? \mergeHP_CTmain_map'_Int_Bool_selected  :
                                              2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_map'_Int_Bool,Go) > (incrHP_mergeCTmain_map'_Int_Bool_buf,Go) */
  Go_t \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d ;
  logic \incrHP_mergeCTmain_map'_Int_Bool_bufchan_r ;
  assign \incrHP_mergeCTmain_map'_Int_Bool_r  = ((! \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d [0]) || \incrHP_mergeCTmain_map'_Int_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmain_map'_Int_Bool_r )
        \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d  <= \incrHP_mergeCTmain_map'_Int_Bool_d ;
  Go_t \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf ;
  assign \incrHP_mergeCTmain_map'_Int_Bool_bufchan_r  = (! \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf [0]);
  assign \incrHP_mergeCTmain_map'_Int_Bool_buf_d  = (\incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf [0] ? \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf  :
                                                     \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmain_map'_Int_Bool_buf_r  && \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf [0]))
        \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmain_map'_Int_Bool_buf_r ) && (! \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf [0])))
        \incrHP_mergeCTmain_map'_Int_Bool_bufchan_buf  <= \incrHP_mergeCTmain_map'_Int_Bool_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_map'_Int_Bool,Word16#) > (mergeHP_CTmain_map'_Int_Bool_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmain_map'_Int_Bool_bufchan_d ;
  logic \mergeHP_CTmain_map'_Int_Bool_bufchan_r ;
  assign \mergeHP_CTmain_map'_Int_Bool_r  = ((! \mergeHP_CTmain_map'_Int_Bool_bufchan_d [0]) || \mergeHP_CTmain_map'_Int_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Bool_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmain_map'_Int_Bool_r )
        \mergeHP_CTmain_map'_Int_Bool_bufchan_d  <= \mergeHP_CTmain_map'_Int_Bool_d ;
  \Word16#_t  \mergeHP_CTmain_map'_Int_Bool_bufchan_buf ;
  assign \mergeHP_CTmain_map'_Int_Bool_bufchan_r  = (! \mergeHP_CTmain_map'_Int_Bool_bufchan_buf [0]);
  assign \mergeHP_CTmain_map'_Int_Bool_buf_d  = (\mergeHP_CTmain_map'_Int_Bool_bufchan_buf [0] ? \mergeHP_CTmain_map'_Int_Bool_bufchan_buf  :
                                                 \mergeHP_CTmain_map'_Int_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Bool_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTmain_map'_Int_Bool_buf_r  && \mergeHP_CTmain_map'_Int_Bool_bufchan_buf [0]))
        \mergeHP_CTmain_map'_Int_Bool_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTmain_map'_Int_Bool_buf_r ) && (! \mergeHP_CTmain_map'_Int_Bool_bufchan_buf [0])))
        \mergeHP_CTmain_map'_Int_Bool_bufchan_buf  <= \mergeHP_CTmain_map'_Int_Bool_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_map'_Int_Bool_buf,Word16#) > [(forkHP1_CTmain_map'_Int_Bool,Word16#),
                                                                  (forkHP1_CTmain_map'_Int_Boo2,Word16#),
                                                                  (forkHP1_CTmain_map'_Int_Boo3,Word16#)] */
  logic [2:0] \mergeHP_CTmain_map'_Int_Bool_buf_emitted ;
  logic [2:0] \mergeHP_CTmain_map'_Int_Bool_buf_done ;
  assign \forkHP1_CTmain_map'_Int_Bool_d  = {\mergeHP_CTmain_map'_Int_Bool_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Int_Bool_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Bool_buf_emitted [0]))};
  assign \forkHP1_CTmain_map'_Int_Boo2_d  = {\mergeHP_CTmain_map'_Int_Bool_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Int_Bool_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Bool_buf_emitted [1]))};
  assign \forkHP1_CTmain_map'_Int_Boo3_d  = {\mergeHP_CTmain_map'_Int_Bool_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Int_Bool_buf_d [0] && (! \mergeHP_CTmain_map'_Int_Bool_buf_emitted [2]))};
  assign \mergeHP_CTmain_map'_Int_Bool_buf_done  = (\mergeHP_CTmain_map'_Int_Bool_buf_emitted  | ({\forkHP1_CTmain_map'_Int_Boo3_d [0],
                                                                                                   \forkHP1_CTmain_map'_Int_Boo2_d [0],
                                                                                                   \forkHP1_CTmain_map'_Int_Bool_d [0]} & {\forkHP1_CTmain_map'_Int_Boo3_r ,
                                                                                                                                           \forkHP1_CTmain_map'_Int_Boo2_r ,
                                                                                                                                           \forkHP1_CTmain_map'_Int_Bool_r }));
  assign \mergeHP_CTmain_map'_Int_Bool_buf_r  = (& \mergeHP_CTmain_map'_Int_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Int_Bool_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmain_map'_Int_Bool_buf_emitted  <= (\mergeHP_CTmain_map'_Int_Bool_buf_r  ? 3'd0 :
                                                     \mergeHP_CTmain_map'_Int_Bool_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_map'_Int_Bool) : [(dconReadIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool),
                                             (dconWriteIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool)] > (memMergeChoice_CTmain_map'_Int_Bool,C2) (memMergeIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool) */
  logic [1:0] \dconReadIn_CTmain_map'_Int_Bool_select_d ;
  assign \dconReadIn_CTmain_map'_Int_Bool_select_d  = ((| \dconReadIn_CTmain_map'_Int_Bool_select_q ) ? \dconReadIn_CTmain_map'_Int_Bool_select_q  :
                                                       (\dconReadIn_CTmain_map'_Int_Bool_d [0] ? 2'd1 :
                                                        (\dconWriteIn_CTmain_map'_Int_Bool_d [0] ? 2'd2 :
                                                         2'd0)));
  logic [1:0] \dconReadIn_CTmain_map'_Int_Bool_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Int_Bool_select_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Int_Bool_select_q  <= (\dconReadIn_CTmain_map'_Int_Bool_done  ? 2'd0 :
                                                     \dconReadIn_CTmain_map'_Int_Bool_select_d );
  logic [1:0] \dconReadIn_CTmain_map'_Int_Bool_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Int_Bool_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Int_Bool_emit_q  <= (\dconReadIn_CTmain_map'_Int_Bool_done  ? 2'd0 :
                                                   \dconReadIn_CTmain_map'_Int_Bool_emit_d );
  logic [1:0] \dconReadIn_CTmain_map'_Int_Bool_emit_d ;
  assign \dconReadIn_CTmain_map'_Int_Bool_emit_d  = (\dconReadIn_CTmain_map'_Int_Bool_emit_q  | ({\memMergeChoice_CTmain_map'_Int_Bool_d [0],
                                                                                                  \memMergeIn_CTmain_map'_Int_Bool_d [0]} & {\memMergeChoice_CTmain_map'_Int_Bool_r ,
                                                                                                                                             \memMergeIn_CTmain_map'_Int_Bool_r }));
  logic \dconReadIn_CTmain_map'_Int_Bool_done ;
  assign \dconReadIn_CTmain_map'_Int_Bool_done  = (& \dconReadIn_CTmain_map'_Int_Bool_emit_d );
  assign {\dconWriteIn_CTmain_map'_Int_Bool_r ,
          \dconReadIn_CTmain_map'_Int_Bool_r } = (\dconReadIn_CTmain_map'_Int_Bool_done  ? \dconReadIn_CTmain_map'_Int_Bool_select_d  :
                                                  2'd0);
  assign \memMergeIn_CTmain_map'_Int_Bool_d  = ((\dconReadIn_CTmain_map'_Int_Bool_select_d [0] && (! \dconReadIn_CTmain_map'_Int_Bool_emit_q [0])) ? \dconReadIn_CTmain_map'_Int_Bool_d  :
                                                ((\dconReadIn_CTmain_map'_Int_Bool_select_d [1] && (! \dconReadIn_CTmain_map'_Int_Bool_emit_q [0])) ? \dconWriteIn_CTmain_map'_Int_Bool_d  :
                                                 {84'd0, 1'd0}));
  assign \memMergeChoice_CTmain_map'_Int_Bool_d  = ((\dconReadIn_CTmain_map'_Int_Bool_select_d [0] && (! \dconReadIn_CTmain_map'_Int_Bool_emit_q [1])) ? C1_2_dc(1'd1) :
                                                    ((\dconReadIn_CTmain_map'_Int_Bool_select_d [1] && (! \dconReadIn_CTmain_map'_Int_Bool_emit_q [1])) ? C2_2_dc(1'd1) :
                                                     {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_map'_Int_Bool,
      Ty MemOut_CTmain_map'_Int_Bool) : (memMergeIn_CTmain_map'_Int_Bool_dbuf,MemIn_CTmain_map'_Int_Bool) > (memOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool) */
  logic [66:0] \memMergeIn_CTmain_map'_Int_Bool_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmain_map'_Int_Bool_dbuf_address ;
  logic [66:0] \memMergeIn_CTmain_map'_Int_Bool_dbuf_din ;
  logic [66:0] \memOut_CTmain_map'_Int_Bool_q ;
  logic \memOut_CTmain_map'_Int_Bool_valid ;
  logic \memMergeIn_CTmain_map'_Int_Bool_dbuf_we ;
  logic \memOut_CTmain_map'_Int_Bool_we ;
  assign \memMergeIn_CTmain_map'_Int_Bool_dbuf_din  = \memMergeIn_CTmain_map'_Int_Bool_dbuf_d [84:18];
  assign \memMergeIn_CTmain_map'_Int_Bool_dbuf_address  = \memMergeIn_CTmain_map'_Int_Bool_dbuf_d [17:2];
  assign \memMergeIn_CTmain_map'_Int_Bool_dbuf_we  = (\memMergeIn_CTmain_map'_Int_Bool_dbuf_d [1:1] && \memMergeIn_CTmain_map'_Int_Bool_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmain_map'_Int_Bool_we  <= 1'd0;
        \memOut_CTmain_map'_Int_Bool_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmain_map'_Int_Bool_we  <= \memMergeIn_CTmain_map'_Int_Bool_dbuf_we ;
        \memOut_CTmain_map'_Int_Bool_valid  <= \memMergeIn_CTmain_map'_Int_Bool_dbuf_d [0];
        if (\memMergeIn_CTmain_map'_Int_Bool_dbuf_we )
          begin
            \memMergeIn_CTmain_map'_Int_Bool_dbuf_mem [\memMergeIn_CTmain_map'_Int_Bool_dbuf_address ] <= \memMergeIn_CTmain_map'_Int_Bool_dbuf_din ;
            \memOut_CTmain_map'_Int_Bool_q  <= \memMergeIn_CTmain_map'_Int_Bool_dbuf_din ;
          end
        else
          \memOut_CTmain_map'_Int_Bool_q  <= \memMergeIn_CTmain_map'_Int_Bool_dbuf_mem [\memMergeIn_CTmain_map'_Int_Bool_dbuf_address ];
      end
  assign \memOut_CTmain_map'_Int_Bool_d  = {\memOut_CTmain_map'_Int_Bool_q ,
                                            \memOut_CTmain_map'_Int_Bool_we ,
                                            \memOut_CTmain_map'_Int_Bool_valid };
  assign \memMergeIn_CTmain_map'_Int_Bool_dbuf_r  = ((! \memOut_CTmain_map'_Int_Bool_valid ) || \memOut_CTmain_map'_Int_Bool_r );
  logic [31:0] \profiling_MemIn_CTmain_map'_Int_Bool_read ;
  logic [31:0] \profiling_MemIn_CTmain_map'_Int_Bool_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTmain_map'_Int_Bool_write  <= 0;
        \profiling_MemIn_CTmain_map'_Int_Bool_read  <= 0;
      end
    else
      if ((\memMergeIn_CTmain_map'_Int_Bool_dbuf_we  == 1'd1))
        \profiling_MemIn_CTmain_map'_Int_Bool_write  <= (\profiling_MemIn_CTmain_map'_Int_Bool_write  + 1);
      else
        if ((\memOut_CTmain_map'_Int_Bool_valid  == 1'd1))
          \profiling_MemIn_CTmain_map'_Int_Bool_read  <= (\profiling_MemIn_CTmain_map'_Int_Bool_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_map'_Int_Bool) : (memMergeChoice_CTmain_map'_Int_Bool,C2) (memOut_CTmain_map'_Int_Bool_dbuf,MemOut_CTmain_map'_Int_Bool) > [(memReadOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool),
                                                                                                                                                    (memWriteOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool)] */
  logic [1:0] \memOut_CTmain_map'_Int_Bool_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmain_map'_Int_Bool_d [0] && \memOut_CTmain_map'_Int_Bool_dbuf_d [0]))
      unique case (\memMergeChoice_CTmain_map'_Int_Bool_d [1:1])
        1'd0: \memOut_CTmain_map'_Int_Bool_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmain_map'_Int_Bool_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmain_map'_Int_Bool_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmain_map'_Int_Bool_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmain_map'_Int_Bool_d  = {\memOut_CTmain_map'_Int_Bool_dbuf_d [68:1],
                                                \memOut_CTmain_map'_Int_Bool_dbuf_onehotd [0]};
  assign \memWriteOut_CTmain_map'_Int_Bool_d  = {\memOut_CTmain_map'_Int_Bool_dbuf_d [68:1],
                                                 \memOut_CTmain_map'_Int_Bool_dbuf_onehotd [1]};
  assign \memOut_CTmain_map'_Int_Bool_dbuf_r  = (| (\memOut_CTmain_map'_Int_Bool_dbuf_onehotd  & {\memWriteOut_CTmain_map'_Int_Bool_r ,
                                                                                                  \memReadOut_CTmain_map'_Int_Bool_r }));
  assign \memMergeChoice_CTmain_map'_Int_Bool_r  = \memOut_CTmain_map'_Int_Bool_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmain_map'_Int_Bool) : (memMergeIn_CTmain_map'_Int_Bool_rbuf,MemIn_CTmain_map'_Int_Bool) > (memMergeIn_CTmain_map'_Int_Bool_dbuf,MemIn_CTmain_map'_Int_Bool) */
  assign \memMergeIn_CTmain_map'_Int_Bool_rbuf_r  = ((! \memMergeIn_CTmain_map'_Int_Bool_dbuf_d [0]) || \memMergeIn_CTmain_map'_Int_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Int_Bool_dbuf_d  <= {84'd0, 1'd0};
    else
      if (\memMergeIn_CTmain_map'_Int_Bool_rbuf_r )
        \memMergeIn_CTmain_map'_Int_Bool_dbuf_d  <= \memMergeIn_CTmain_map'_Int_Bool_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmain_map'_Int_Bool) : (memMergeIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool) > (memMergeIn_CTmain_map'_Int_Bool_rbuf,MemIn_CTmain_map'_Int_Bool) */
  \MemIn_CTmain_map'_Int_Bool_t  \memMergeIn_CTmain_map'_Int_Bool_buf ;
  assign \memMergeIn_CTmain_map'_Int_Bool_r  = (! \memMergeIn_CTmain_map'_Int_Bool_buf [0]);
  assign \memMergeIn_CTmain_map'_Int_Bool_rbuf_d  = (\memMergeIn_CTmain_map'_Int_Bool_buf [0] ? \memMergeIn_CTmain_map'_Int_Bool_buf  :
                                                     \memMergeIn_CTmain_map'_Int_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Int_Bool_buf  <= {84'd0, 1'd0};
    else
      if ((\memMergeIn_CTmain_map'_Int_Bool_rbuf_r  && \memMergeIn_CTmain_map'_Int_Bool_buf [0]))
        \memMergeIn_CTmain_map'_Int_Bool_buf  <= {84'd0, 1'd0};
      else if (((! \memMergeIn_CTmain_map'_Int_Bool_rbuf_r ) && (! \memMergeIn_CTmain_map'_Int_Bool_buf [0])))
        \memMergeIn_CTmain_map'_Int_Bool_buf  <= \memMergeIn_CTmain_map'_Int_Bool_d ;
  
  /* dbuf (Ty MemOut_CTmain_map'_Int_Bool) : (memOut_CTmain_map'_Int_Bool_rbuf,MemOut_CTmain_map'_Int_Bool) > (memOut_CTmain_map'_Int_Bool_dbuf,MemOut_CTmain_map'_Int_Bool) */
  assign \memOut_CTmain_map'_Int_Bool_rbuf_r  = ((! \memOut_CTmain_map'_Int_Bool_dbuf_d [0]) || \memOut_CTmain_map'_Int_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Int_Bool_dbuf_d  <= {68'd0, 1'd0};
    else
      if (\memOut_CTmain_map'_Int_Bool_rbuf_r )
        \memOut_CTmain_map'_Int_Bool_dbuf_d  <= \memOut_CTmain_map'_Int_Bool_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmain_map'_Int_Bool) : (memOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool) > (memOut_CTmain_map'_Int_Bool_rbuf,MemOut_CTmain_map'_Int_Bool) */
  \MemOut_CTmain_map'_Int_Bool_t  \memOut_CTmain_map'_Int_Bool_buf ;
  assign \memOut_CTmain_map'_Int_Bool_r  = (! \memOut_CTmain_map'_Int_Bool_buf [0]);
  assign \memOut_CTmain_map'_Int_Bool_rbuf_d  = (\memOut_CTmain_map'_Int_Bool_buf [0] ? \memOut_CTmain_map'_Int_Bool_buf  :
                                                 \memOut_CTmain_map'_Int_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Int_Bool_buf  <= {68'd0, 1'd0};
    else
      if ((\memOut_CTmain_map'_Int_Bool_rbuf_r  && \memOut_CTmain_map'_Int_Bool_buf [0]))
        \memOut_CTmain_map'_Int_Bool_buf  <= {68'd0, 1'd0};
      else if (((! \memOut_CTmain_map'_Int_Bool_rbuf_r ) && (! \memOut_CTmain_map'_Int_Bool_buf [0])))
        \memOut_CTmain_map'_Int_Bool_buf  <= \memOut_CTmain_map'_Int_Bool_d ;
  
  /* destruct (Ty Pointer_CTmain_map'_Int_Bool,
          Dcon Pointer_CTmain_map'_Int_Bool) : (scfarg_0_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) > [(destructReadIn_CTmain_map'_Int_Bool,Word16#)] */
  assign \destructReadIn_CTmain_map'_Int_Bool_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                                    scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTmain_map'_Int_Bool_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Int_Bool,
      Dcon ReadIn_CTmain_map'_Int_Bool) : [(destructReadIn_CTmain_map'_Int_Bool,Word16#)] > (dconReadIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool) */
  assign \dconReadIn_CTmain_map'_Int_Bool_d  = \ReadIn_CTmain_map'_Int_Bool_dc ((& {\destructReadIn_CTmain_map'_Int_Bool_d [0]}), \destructReadIn_CTmain_map'_Int_Bool_d );
  assign {\destructReadIn_CTmain_map'_Int_Bool_r } = {1 {(\dconReadIn_CTmain_map'_Int_Bool_r  && \dconReadIn_CTmain_map'_Int_Bool_d [0])}};
  
  /* destruct (Ty MemOut_CTmain_map'_Int_Bool,
          Dcon ReadOut_CTmain_map'_Int_Bool) : (memReadOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool) > [(readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf,CTmain_map'_Int_Bool)] */
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_d  = {\memReadOut_CTmain_map'_Int_Bool_d [68:2],
                                                                    \memReadOut_CTmain_map'_Int_Bool_d [0]};
  assign \memReadOut_CTmain_map'_Int_Bool_r  = \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmain_map'_Int_Bool) : [(lizzieLet21_1_argbuf,CTmain_map'_Int_Bool),
                                       (lizzieLet23_1_argbuf,CTmain_map'_Int_Bool),
                                       (lizzieLet34_1_argbuf,CTmain_map'_Int_Bool),
                                       (lizzieLet35_1_argbuf,CTmain_map'_Int_Bool),
                                       (lizzieLet36_1_argbuf,CTmain_map'_Int_Bool)] > (writeMerge_choice_CTmain_map'_Int_Bool,C5) (writeMerge_data_CTmain_map'_Int_Bool,CTmain_map'_Int_Bool) */
  logic [4:0] lizzieLet21_1_argbuf_select_d;
  assign lizzieLet21_1_argbuf_select_d = ((| lizzieLet21_1_argbuf_select_q) ? lizzieLet21_1_argbuf_select_q :
                                          (lizzieLet21_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet23_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet34_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet35_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet36_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet21_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet21_1_argbuf_select_q <= (lizzieLet21_1_argbuf_done ? 5'd0 :
                                        lizzieLet21_1_argbuf_select_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet21_1_argbuf_emit_q <= (lizzieLet21_1_argbuf_done ? 2'd0 :
                                      lizzieLet21_1_argbuf_emit_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_d;
  assign lizzieLet21_1_argbuf_emit_d = (lizzieLet21_1_argbuf_emit_q | ({\writeMerge_choice_CTmain_map'_Int_Bool_d [0],
                                                                        \writeMerge_data_CTmain_map'_Int_Bool_d [0]} & {\writeMerge_choice_CTmain_map'_Int_Bool_r ,
                                                                                                                        \writeMerge_data_CTmain_map'_Int_Bool_r }));
  logic lizzieLet21_1_argbuf_done;
  assign lizzieLet21_1_argbuf_done = (& lizzieLet21_1_argbuf_emit_d);
  assign {lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet34_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet21_1_argbuf_r} = (lizzieLet21_1_argbuf_done ? lizzieLet21_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmain_map'_Int_Bool_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                                     ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                      ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet34_1_argbuf_d :
                                                       ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                        ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                         {67'd0, 1'd0})))));
  assign \writeMerge_choice_CTmain_map'_Int_Bool_d  = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                       ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                        ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                         ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                          ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                           {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_map'_Int_Bool) : (writeMerge_choice_CTmain_map'_Int_Bool,C5) (demuxWriteResult_CTmain_map'_Int_Bool,Pointer_CTmain_map'_Int_Bool) > [(writeCTmain_map'_Int_BoollizzieLet21_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                                                                                                              (writeCTmain_map'_Int_BoollizzieLet23_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                                                                                                              (writeCTmain_map'_Int_BoollizzieLet34_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                                                                                                              (writeCTmain_map'_Int_BoollizzieLet35_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                                                                                                              (writeCTmain_map'_Int_BoollizzieLet36_1_argbuf,Pointer_CTmain_map'_Int_Bool)] */
  logic [4:0] \demuxWriteResult_CTmain_map'_Int_Bool_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmain_map'_Int_Bool_d [0] && \demuxWriteResult_CTmain_map'_Int_Bool_d [0]))
      unique case (\writeMerge_choice_CTmain_map'_Int_Bool_d [3:1])
        3'd0: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd16;
        default: \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTmain_map'_Int_Bool_onehotd  = 5'd0;
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Bool_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Int_Bool_onehotd [0]};
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Bool_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Int_Bool_onehotd [1]};
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Bool_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Int_Bool_onehotd [2]};
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Bool_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Int_Bool_onehotd [3]};
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Int_Bool_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Int_Bool_onehotd [4]};
  assign \demuxWriteResult_CTmain_map'_Int_Bool_r  = (| (\demuxWriteResult_CTmain_map'_Int_Bool_onehotd  & {\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_r }));
  assign \writeMerge_choice_CTmain_map'_Int_Bool_r  = \demuxWriteResult_CTmain_map'_Int_Bool_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Int_Bool,
      Dcon WriteIn_CTmain_map'_Int_Bool) : [(forkHP1_CTmain_map'_Int_Boo2,Word16#),
                                            (writeMerge_data_CTmain_map'_Int_Bool,CTmain_map'_Int_Bool)] > (dconWriteIn_CTmain_map'_Int_Bool,MemIn_CTmain_map'_Int_Bool) */
  assign \dconWriteIn_CTmain_map'_Int_Bool_d  = \WriteIn_CTmain_map'_Int_Bool_dc ((& {\forkHP1_CTmain_map'_Int_Boo2_d [0],
                                                                                      \writeMerge_data_CTmain_map'_Int_Bool_d [0]}), \forkHP1_CTmain_map'_Int_Boo2_d , \writeMerge_data_CTmain_map'_Int_Bool_d );
  assign {\forkHP1_CTmain_map'_Int_Boo2_r ,
          \writeMerge_data_CTmain_map'_Int_Bool_r } = {2 {(\dconWriteIn_CTmain_map'_Int_Bool_r  && \dconWriteIn_CTmain_map'_Int_Bool_d [0])}};
  
  /* dcon (Ty Pointer_CTmain_map'_Int_Bool,
      Dcon Pointer_CTmain_map'_Int_Bool) : [(forkHP1_CTmain_map'_Int_Boo3,Word16#)] > (dconPtr_CTmain_map'_Int_Bool,Pointer_CTmain_map'_Int_Bool) */
  assign \dconPtr_CTmain_map'_Int_Bool_d  = \Pointer_CTmain_map'_Int_Bool_dc ((& {\forkHP1_CTmain_map'_Int_Boo3_d [0]}), \forkHP1_CTmain_map'_Int_Boo3_d );
  assign {\forkHP1_CTmain_map'_Int_Boo3_r } = {1 {(\dconPtr_CTmain_map'_Int_Bool_r  && \dconPtr_CTmain_map'_Int_Bool_d [0])}};
  
  /* demux (Ty MemOut_CTmain_map'_Int_Bool,
       Ty Pointer_CTmain_map'_Int_Bool) : (memWriteOut_CTmain_map'_Int_Bool,MemOut_CTmain_map'_Int_Bool) (dconPtr_CTmain_map'_Int_Bool,Pointer_CTmain_map'_Int_Bool) > [(_60,Pointer_CTmain_map'_Int_Bool),
                                                                                                                                                                        (demuxWriteResult_CTmain_map'_Int_Bool,Pointer_CTmain_map'_Int_Bool)] */
  logic [1:0] \dconPtr_CTmain_map'_Int_Bool_onehotd ;
  always_comb
    if ((\memWriteOut_CTmain_map'_Int_Bool_d [0] && \dconPtr_CTmain_map'_Int_Bool_d [0]))
      unique case (\memWriteOut_CTmain_map'_Int_Bool_d [1:1])
        1'd0: \dconPtr_CTmain_map'_Int_Bool_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmain_map'_Int_Bool_onehotd  = 2'd2;
        default: \dconPtr_CTmain_map'_Int_Bool_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmain_map'_Int_Bool_onehotd  = 2'd0;
  assign _60_d = {\dconPtr_CTmain_map'_Int_Bool_d [16:1],
                  \dconPtr_CTmain_map'_Int_Bool_onehotd [0]};
  assign \demuxWriteResult_CTmain_map'_Int_Bool_d  = {\dconPtr_CTmain_map'_Int_Bool_d [16:1],
                                                      \dconPtr_CTmain_map'_Int_Bool_onehotd [1]};
  assign \dconPtr_CTmain_map'_Int_Bool_r  = (| (\dconPtr_CTmain_map'_Int_Bool_onehotd  & {\demuxWriteResult_CTmain_map'_Int_Bool_r ,
                                                                                          _60_r}));
  assign \memWriteOut_CTmain_map'_Int_Bool_r  = \dconPtr_CTmain_map'_Int_Bool_r ;
  
  /* buf (Ty Go) : (goFork,Go) > (go_1_argbuf,Go) */
  Go_t goFork_bufchan_d;
  logic goFork_bufchan_r;
  assign goFork_r = ((! goFork_bufchan_d[0]) || goFork_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_d <= 1'd0;
    else if (goFork_r) goFork_bufchan_d <= goFork_d;
  Go_t goFork_bufchan_buf;
  assign goFork_bufchan_r = (! goFork_bufchan_buf[0]);
  assign go_1_argbuf_d = (goFork_bufchan_buf[0] ? goFork_bufchan_buf :
                          goFork_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) goFork_bufchan_buf <= 1'd0;
    else
      if ((go_1_argbuf_r && goFork_bufchan_buf[0]))
        goFork_bufchan_buf <= 1'd0;
      else if (((! go_1_argbuf_r) && (! goFork_bufchan_buf[0])))
        goFork_bufchan_buf <= goFork_bufchan_d;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (w1sm4_1_1,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (wsm3_1_0,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) > [($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6,Go),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR,MyDTInt_Int_Int),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS,Pointer_QTree_Int),
                                                                                                                                                                                                                                   ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT,Pointer_QTree_Int)] */
  logic [3:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted ;
  logic [3:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_d  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [0]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_d  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [1]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_d  = {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [16:1],
                                                                                               (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [2]))};
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_d  = {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [32:17],
                                                                                               (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [3]))};
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  | ({\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_d [0],
                                                                                                                                                                                         \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_d [0]} & {\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_r ,
                                                                                                                                                                                                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_r }));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  = (& \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= 4'd0;
    else
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  ? 4'd0 :
                                                                                                \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6,Go) > [(go_6_1,Go),
                                                                                                     (go_6_2,Go)] */
  logic [1:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted ;
  logic [1:0] \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_done ;
  assign go_6_1_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted [0]));
  assign go_6_2_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_d [0] && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted [1]));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_done  = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted  | ({go_6_2_d[0],
                                                                                                                                                                                             go_6_1_d[0]} & {go_6_2_r,
                                                                                                                                                                                                             go_6_1_r}));
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_r  = (& \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted  <= 2'd0;
    else
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_emitted  <= (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_r  ? 2'd0 :
                                                                                                  \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intgo_6_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS,Pointer_QTree_Int) > (w1slS_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d  <= {16'd0,
                                                                                                     1'd0};
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_d ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf [0]);
  assign w1slS_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf  :
                             \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf  <= {16'd0,
                                                                                                       1'd0};
    else
      if ((w1slS_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
      else if (((! w1slS_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw1slS_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT,Pointer_QTree_Int) > (w2slT_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d  <= {16'd0,
                                                                                                     1'd0};
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_d ;
  Pointer_QTree_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf [0]);
  assign w2slT_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf  :
                             \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf  <= {16'd0,
                                                                                                       1'd0};
    else
      if ((w2slT_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
      else if (((! w2slT_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Intw2slT_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int_Int) : ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR,MyDTInt_Int_Int) > (wslR_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d ;
  logic \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_r ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_r  = ((! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d [0]) || \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d  <= 1'd0;
    else
      if (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_r )
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_d ;
  MyDTInt_Int_Int_t \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf ;
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_r  = (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf [0]);
  assign wslR_1_argbuf_d = (\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf [0] ? \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf  :
                            \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf  <= 1'd0;
    else
      if ((wslR_1_argbuf_r && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf [0]))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf  <= 1'd0;
      else if (((! wslR_1_argbuf_r) && (! \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf [0])))
        \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_buf  <= \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_IntwslR_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmAdd_Int_resbuf,Pointer_QTree_Int) > (es_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_bufchan_d ;
  logic \$wmAdd_Int_resbuf_bufchan_r ;
  assign \$wmAdd_Int_resbuf_r  = ((! \$wmAdd_Int_resbuf_bufchan_d [0]) || \$wmAdd_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wmAdd_Int_resbuf_r )
        \$wmAdd_Int_resbuf_bufchan_d  <= \$wmAdd_Int_resbuf_d ;
  Pointer_QTree_Int_t \$wmAdd_Int_resbuf_bufchan_buf ;
  assign \$wmAdd_Int_resbuf_bufchan_r  = (! \$wmAdd_Int_resbuf_bufchan_buf [0]);
  assign es_3_1_argbuf_d = (\$wmAdd_Int_resbuf_bufchan_buf [0] ? \$wmAdd_Int_resbuf_bufchan_buf  :
                            \$wmAdd_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((es_3_1_argbuf_r && \$wmAdd_Int_resbuf_bufchan_buf [0]))
        \$wmAdd_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! es_3_1_argbuf_r) && (! \$wmAdd_Int_resbuf_bufchan_buf [0])))
        \$wmAdd_Int_resbuf_bufchan_buf  <= \$wmAdd_Int_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) > [($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7,Go),
                                                                                                                                                                         ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3,Pointer_QTree_Int),
                                                                                                                                                                         ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4,Pointer_QTree_Int)] */
  logic [2:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted ;
  logic [2:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [0]));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_d  = {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [16:1],
                                                                        (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_d  = {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [32:17],
                                                                         (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted [2]))};
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  | ({\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_d [0],
                                                                                                                                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_d [0],
                                                                                                                                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0]} & {\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_r ,
                                                                                                                                                                                                                \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_r ,
                                                                                                                                                                                                                \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r }));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  = (& \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= 3'd0;
    else
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_emitted  <= (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  ? 3'd0 :
                                                                          \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7,Go) > [(go_7_1,Go),
                                                                               (go_7_2,Go),
                                                                               (go_7_3,Go),
                                                                               (go_7_4,Go),
                                                                               (go_7_5,Go),
                                                                               (go_7_6,Go)] */
  logic [5:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted ;
  logic [5:0] \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done ;
  assign go_7_1_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [0]));
  assign go_7_2_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [1]));
  assign go_7_3_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [2]));
  assign go_7_4_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [3]));
  assign go_7_5_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [4]));
  assign go_7_6_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_d [0] && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted [5]));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done  = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  | ({go_7_6_d[0],
                                                                                                                                                 go_7_5_d[0],
                                                                                                                                                 go_7_4_d[0],
                                                                                                                                                 go_7_3_d[0],
                                                                                                                                                 go_7_2_d[0],
                                                                                                                                                 go_7_1_d[0]} & {go_7_6_r,
                                                                                                                                                                 go_7_5_r,
                                                                                                                                                                 go_7_4_r,
                                                                                                                                                                 go_7_3_r,
                                                                                                                                                                 go_7_2_r,
                                                                                                                                                                 go_7_1_r}));
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r  = (& \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  <= 6'd0;
    else
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_emitted  <= (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_r  ? 6'd0 :
                                                                            \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intgo_7_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4,Pointer_QTree_Int) > (w1sm4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_r ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_r  = ((! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d [0]) || \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d  <= {16'd0,
                                                                               1'd0};
    else
      if (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_r )
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_d ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_r  = (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf [0]);
  assign w1sm4_1_argbuf_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf [0] ? \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf  :
                             \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
    else
      if ((w1sm4_1_argbuf_r && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf [0]))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf  <= {16'd0,
                                                                                   1'd0};
      else if (((! w1sm4_1_argbuf_r) && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf [0])))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_buf  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intw1sm4_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3,Pointer_QTree_Int) > (wsm3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d ;
  logic \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_r ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_r  = ((! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d [0]) || \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d  <= {16'd0,
                                                                              1'd0};
    else
      if (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_r )
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_d ;
  Pointer_QTree_Int_t \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf ;
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_r  = (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf [0]);
  assign wsm3_1_argbuf_d = (\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf [0] ? \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf  :
                            \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf  <= {16'd0,
                                                                                1'd0};
    else
      if ((wsm3_1_argbuf_r && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf [0]))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
      else if (((! wsm3_1_argbuf_r) && (! \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf [0])))
        \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_buf  <= \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Intwsm3_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wmain_resbuf,Int#)] > (es_0_1I#,Int) */
  assign \es_0_1I#_d  = \I#_dc ((& {\$wmain_resbuf_d [0]}), \$wmain_resbuf_d );
  assign {\$wmain_resbuf_r } = {1 {(\es_0_1I#_r  && \es_0_1I#_d [0])}};
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool,
          Dcon TupGo___Pointer_QTree_Bool) : ($wnnzTupGo___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool) > [($wnnzTupGo___Pointer_QTree_Boolgo_8,Go),
                                                                                                               ($wnnzTupGo___Pointer_QTree_BoolwslW,Pointer_QTree_Bool)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Bool_1_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Bool_1_done ;
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_8_d  = (\$wnnzTupGo___Pointer_QTree_Bool_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Bool_1_emitted [0]));
  assign \$wnnzTupGo___Pointer_QTree_BoolwslW_d  = {\$wnnzTupGo___Pointer_QTree_Bool_1_d [16:1],
                                                    (\$wnnzTupGo___Pointer_QTree_Bool_1_d [0] && (! \$wnnzTupGo___Pointer_QTree_Bool_1_emitted [1]))};
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_done  = (\$wnnzTupGo___Pointer_QTree_Bool_1_emitted  | ({\$wnnzTupGo___Pointer_QTree_BoolwslW_d [0],
                                                                                                     \$wnnzTupGo___Pointer_QTree_Boolgo_8_d [0]} & {\$wnnzTupGo___Pointer_QTree_BoolwslW_r ,
                                                                                                                                                    \$wnnzTupGo___Pointer_QTree_Boolgo_8_r }));
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_r  = (& \$wnnzTupGo___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Bool_1_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Bool_1_emitted  <= (\$wnnzTupGo___Pointer_QTree_Bool_1_r  ? 2'd0 :
                                                      \$wnnzTupGo___Pointer_QTree_Bool_1_done );
  
  /* fork (Ty Go) : ($wnnzTupGo___Pointer_QTree_Boolgo_8,Go) > [(go_8_1,Go),
                                                           (go_8_2,Go)] */
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted ;
  logic [1:0] \$wnnzTupGo___Pointer_QTree_Boolgo_8_done ;
  assign go_8_1_d = (\$wnnzTupGo___Pointer_QTree_Boolgo_8_d [0] && (! \$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted [0]));
  assign go_8_2_d = (\$wnnzTupGo___Pointer_QTree_Boolgo_8_d [0] && (! \$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted [1]));
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_8_done  = (\$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted  | ({go_8_2_d[0],
                                                                                                         go_8_1_d[0]} & {go_8_2_r,
                                                                                                                         go_8_1_r}));
  assign \$wnnzTupGo___Pointer_QTree_Boolgo_8_r  = (& \$wnnzTupGo___Pointer_QTree_Boolgo_8_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted  <= 2'd0;
    else
      \$wnnzTupGo___Pointer_QTree_Boolgo_8_emitted  <= (\$wnnzTupGo___Pointer_QTree_Boolgo_8_r  ? 2'd0 :
                                                        \$wnnzTupGo___Pointer_QTree_Boolgo_8_done );
  
  /* buf (Ty Pointer_QTree_Bool) : ($wnnzTupGo___Pointer_QTree_BoolwslW,Pointer_QTree_Bool) > (wslW_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d ;
  logic \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_r ;
  assign \$wnnzTupGo___Pointer_QTree_BoolwslW_r  = ((! \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d [0]) || \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wnnzTupGo___Pointer_QTree_BoolwslW_r )
        \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d  <= \$wnnzTupGo___Pointer_QTree_BoolwslW_d ;
  Pointer_QTree_Bool_t \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf ;
  assign \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_r  = (! \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf [0]);
  assign wslW_1_argbuf_d = (\$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf [0] ? \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf  :
                            \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((wslW_1_argbuf_r && \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf [0]))
        \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! wslW_1_argbuf_r) && (! \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf [0])))
        \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_buf  <= \$wnnzTupGo___Pointer_QTree_BoolwslW_bufchan_d ;
  
  /* buf (Ty Int#) : ($wnnz_resbuf,Int#) > ($wmain_resbuf,Int#) */
  \Int#_t  \$wnnz_resbuf_bufchan_d ;
  logic \$wnnz_resbuf_bufchan_r ;
  assign \$wnnz_resbuf_r  = ((! \$wnnz_resbuf_bufchan_d [0]) || \$wnnz_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \$wnnz_resbuf_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\$wnnz_resbuf_r ) \$wnnz_resbuf_bufchan_d  <= \$wnnz_resbuf_d ;
  \Int#_t  \$wnnz_resbuf_bufchan_buf ;
  assign \$wnnz_resbuf_bufchan_r  = (! \$wnnz_resbuf_bufchan_buf [0]);
  assign \$wmain_resbuf_d  = (\$wnnz_resbuf_bufchan_buf [0] ? \$wnnz_resbuf_bufchan_buf  :
                              \$wnnz_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \$wnnz_resbuf_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\$wmain_resbuf_r  && \$wnnz_resbuf_bufchan_buf [0]))
        \$wnnz_resbuf_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \$wmain_resbuf_r ) && (! \$wnnz_resbuf_bufchan_buf [0])))
        \$wnnz_resbuf_bufchan_buf  <= \$wnnz_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyBool,
          Dcon TupGo___MyDTBool_Bool___MyBool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) > [(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9,Go),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done;
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[1:1],
                                                                   (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted | ({applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d[0]} & {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r ? 3'd0 :
                                                                     applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool) > [(arg0_1,MyDTBool_Bool),
                                                                                                  (arg0_2,MyDTBool_Bool),
                                                                                                  (arg0_3,MyDTBool_Bool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done;
  assign arg0_1_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[0]));
  assign arg0_2_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[1]));
  assign arg0_3_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[2]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted | ({arg0_3_d[0],
                                                                                                                                       arg0_2_d[0],
                                                                                                                                       arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                                       arg0_2_r,
                                                                                                                                                       arg0_1_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r ? 3'd0 :
                                                                       applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  
  /* fork (Ty MyBool) : (applyfnBool_Bool_5_resbuf,MyBool) > [(es_0_4_1,MyBool),
                                                         (es_0_4_2,MyBool),
                                                         (es_0_4_3,MyBool)] */
  logic [2:0] applyfnBool_Bool_5_resbuf_emitted;
  logic [2:0] applyfnBool_Bool_5_resbuf_done;
  assign es_0_4_1_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[0]))};
  assign es_0_4_2_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[1]))};
  assign es_0_4_3_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[2]))};
  assign applyfnBool_Bool_5_resbuf_done = (applyfnBool_Bool_5_resbuf_emitted | ({es_0_4_3_d[0],
                                                                                 es_0_4_2_d[0],
                                                                                 es_0_4_1_d[0]} & {es_0_4_3_r,
                                                                                                   es_0_4_2_r,
                                                                                                   es_0_4_1_r}));
  assign applyfnBool_Bool_5_resbuf_r = (& applyfnBool_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnBool_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnBool_Bool_5_resbuf_emitted <= (applyfnBool_Bool_5_resbuf_r ? 3'd0 :
                                            applyfnBool_Bool_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10,Go),
                                                                                                                           (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2,MyDTInt_Bool),
                                                                                                                           (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[32:1],
                                                                (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted[2]))};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d[0],
                                                                                                                         applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d[0],
                                                                                                                         applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_r,
                                                                                                                                                                                   applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_r,
                                                                                                                                                                                   applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r ? 3'd0 :
                                                                applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done);
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2,MyDTInt_Bool) > [(arg0_2_1,MyDTInt_Bool),
                                                                                             (arg0_2_2,MyDTInt_Bool),
                                                                                             (arg0_2_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                                 arg0_2_2_d[0],
                                                                                                                                 arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                                   arg0_2_2_r,
                                                                                                                                                   arg0_2_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_r ? 3'd0 :
                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_2_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(xa88_1,MyBool),
                                                        (xa88_2,MyBool)] */
  logic [1:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [1:0] applyfnInt_Bool_5_resbuf_done;
  assign xa88_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign xa88_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({xa88_2_d[0],
                                                                               xa88_1_d[0]} & {xa88_2_r,
                                                                                               xa88_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 2'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 2'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[32:1],
                                                                     (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[64:33],
                                                                       (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted[2]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                                                                         applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r ? 3'd0 :
                                                                       applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done);
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int) > [(arg0_4_1,MyDTInt_Int_Int),
                                                                                                          (arg0_4_2,MyDTInt_Int_Int),
                                                                                                          (arg0_4_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done;
  assign arg0_4_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[0]));
  assign arg0_4_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[1]));
  assign arg0_4_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted | ({arg0_4_3_d[0],
                                                                                                                                               arg0_4_2_d[0],
                                                                                                                                               arg0_4_1_d[0]} & {arg0_4_3_r,
                                                                                                                                                                 arg0_4_2_r,
                                                                                                                                                                 arg0_4_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_Int_5_resbuf,Int)] > (es_0_3_1QVal_Int,QTree_Int) */
  assign es_0_3_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_Int_5_resbuf_d[0]}), applyfnInt_Int_Int_5_resbuf_d);
  assign {applyfnInt_Int_Int_5_resbuf_r} = {1 {(es_0_3_1QVal_Int_r && es_0_3_1QVal_Int_d[0])}};
  
  /* demux (Ty MyDTBool_Bool,
       Ty MyBool) : (arg0_1,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool) > [(arg0_1Dcon_main2,MyBool)] */
  assign arg0_1Dcon_main2_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[1:1],
                               (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0])};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r = (arg0_1Dcon_main2_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_main2_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  
  /* fork (Ty MyBool) : (arg0_1Dcon_main2,MyBool) > [(arg0_1Dcon_main2_1,MyBool),
                                                (arg0_1Dcon_main2_2,MyBool)] */
  logic [1:0] arg0_1Dcon_main2_emitted;
  logic [1:0] arg0_1Dcon_main2_done;
  assign arg0_1Dcon_main2_1_d = {arg0_1Dcon_main2_d[1:1],
                                 (arg0_1Dcon_main2_d[0] && (! arg0_1Dcon_main2_emitted[0]))};
  assign arg0_1Dcon_main2_2_d = {arg0_1Dcon_main2_d[1:1],
                                 (arg0_1Dcon_main2_d[0] && (! arg0_1Dcon_main2_emitted[1]))};
  assign arg0_1Dcon_main2_done = (arg0_1Dcon_main2_emitted | ({arg0_1Dcon_main2_2_d[0],
                                                               arg0_1Dcon_main2_1_d[0]} & {arg0_1Dcon_main2_2_r,
                                                                                           arg0_1Dcon_main2_1_r}));
  assign arg0_1Dcon_main2_r = (& arg0_1Dcon_main2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_main2_emitted <= 2'd0;
    else
      arg0_1Dcon_main2_emitted <= (arg0_1Dcon_main2_r ? 2'd0 :
                                   arg0_1Dcon_main2_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_1Dcon_main2_1,MyBool) (arg0_2Dcon_main2,Go) > [(arg0_1Dcon_main2_1MyFalse,Go),
                                                                     (arg0_1Dcon_main2_1MyTrue,Go)] */
  logic [1:0] arg0_2Dcon_main2_onehotd;
  always_comb
    if ((arg0_1Dcon_main2_1_d[0] && arg0_2Dcon_main2_d[0]))
      unique case (arg0_1Dcon_main2_1_d[1:1])
        1'd0: arg0_2Dcon_main2_onehotd = 2'd1;
        1'd1: arg0_2Dcon_main2_onehotd = 2'd2;
        default: arg0_2Dcon_main2_onehotd = 2'd0;
      endcase
    else arg0_2Dcon_main2_onehotd = 2'd0;
  assign arg0_1Dcon_main2_1MyFalse_d = arg0_2Dcon_main2_onehotd[0];
  assign arg0_1Dcon_main2_1MyTrue_d = arg0_2Dcon_main2_onehotd[1];
  assign arg0_2Dcon_main2_r = (| (arg0_2Dcon_main2_onehotd & {arg0_1Dcon_main2_1MyTrue_r,
                                                              arg0_1Dcon_main2_1MyFalse_r}));
  assign arg0_1Dcon_main2_1_r = arg0_2Dcon_main2_r;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(arg0_1Dcon_main2_1MyFalse,Go)] > (arg0_1Dcon_main2_1MyFalse_1MyTrue,MyBool) */
  assign arg0_1Dcon_main2_1MyFalse_1MyTrue_d = MyTrue_dc((& {arg0_1Dcon_main2_1MyFalse_d[0]}), arg0_1Dcon_main2_1MyFalse_d);
  assign {arg0_1Dcon_main2_1MyFalse_r} = {1 {(arg0_1Dcon_main2_1MyFalse_1MyTrue_r && arg0_1Dcon_main2_1MyFalse_1MyTrue_d[0])}};
  
  /* buf (Ty MyBool) : (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux,MyBool) > (applyfnBool_Bool_5_resbuf,MyBool) */
  MyBool_t arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  logic arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_r;
  assign arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_r = ((! arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d[0]) || arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d <= {1'd0,
                                                                                               1'd0};
    else
      if (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_r)
        arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d <= arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_d;
  MyBool_t arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf;
  assign arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_r = (! arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]);
  assign applyfnBool_Bool_5_resbuf_d = (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0] ? arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf :
                                        arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                 1'd0};
    else
      if ((applyfnBool_Bool_5_resbuf_r && arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]))
        arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                   1'd0};
      else if (((! applyfnBool_Bool_5_resbuf_r) && (! arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0])))
        arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(arg0_1Dcon_main2_1MyTrue,Go)] > (arg0_1Dcon_main2_1MyTrue_1MyFalse,MyBool) */
  assign arg0_1Dcon_main2_1MyTrue_1MyFalse_d = MyFalse_dc((& {arg0_1Dcon_main2_1MyTrue_d[0]}), arg0_1Dcon_main2_1MyTrue_d);
  assign {arg0_1Dcon_main2_1MyTrue_r} = {1 {(arg0_1Dcon_main2_1MyTrue_1MyFalse_r && arg0_1Dcon_main2_1MyTrue_1MyFalse_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_1Dcon_main2_2,MyBool) [(arg0_1Dcon_main2_1MyFalse_1MyTrue,MyBool),
                                               (arg0_1Dcon_main2_1MyTrue_1MyFalse,MyBool)] > (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux,MyBool) */
  logic [1:0] arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux;
  logic [1:0] arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_onehot;
  always_comb
    unique case (arg0_1Dcon_main2_2_d[1:1])
      1'd0:
        {arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux} = {2'd1,
                                                                                        arg0_1Dcon_main2_1MyFalse_1MyTrue_d};
      1'd1:
        {arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux} = {2'd2,
                                                                                        arg0_1Dcon_main2_1MyTrue_1MyFalse_d};
      default:
        {arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux} = {2'd0,
                                                                                        {1'd0,
                                                                                         1'd0}};
    endcase
  assign arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d = {arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux[1:1],
                                                                                     (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux[0] && arg0_1Dcon_main2_2_d[0])};
  assign arg0_1Dcon_main2_2_r = (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d[0] && arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_r);
  assign {arg0_1Dcon_main2_1MyTrue_1MyFalse_r,
          arg0_1Dcon_main2_1MyFalse_1MyTrue_r} = (arg0_1Dcon_main2_2_r ? arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_onehot :
                                                  2'd0);
  
  /* demux (Ty MyDTBool_Bool,
       Ty Go) : (arg0_2,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9,Go) > [(arg0_2Dcon_main2,Go)] */
  assign arg0_2Dcon_main2_d = (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d[0]);
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_r = (arg0_2Dcon_main2_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d[0]));
  assign arg0_2_r = (arg0_2Dcon_main2_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_9_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_2_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1,Int) > [(arg0_2_1Dcon_main1,Int)] */
  assign arg0_2_1Dcon_main1_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d[32:1],
                                 (arg0_2_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d[0]));
  assign arg0_2_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_1_d[0]));
  
  /* fork (Ty Int) : (arg0_2_1Dcon_main1,Int) > [(arg0_2_1Dcon_main1_1,Int),
                                            (arg0_2_1Dcon_main1_2,Int),
                                            (arg0_2_1Dcon_main1_3,Int),
                                            (arg0_2_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_2_1Dcon_main1_emitted;
  logic [3:0] arg0_2_1Dcon_main1_done;
  assign arg0_2_1Dcon_main1_1_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[0]))};
  assign arg0_2_1Dcon_main1_2_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[1]))};
  assign arg0_2_1Dcon_main1_3_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[2]))};
  assign arg0_2_1Dcon_main1_4_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[3]))};
  assign arg0_2_1Dcon_main1_done = (arg0_2_1Dcon_main1_emitted | ({arg0_2_1Dcon_main1_4_d[0],
                                                                   arg0_2_1Dcon_main1_3_d[0],
                                                                   arg0_2_1Dcon_main1_2_d[0],
                                                                   arg0_2_1Dcon_main1_1_d[0]} & {arg0_2_1Dcon_main1_4_r,
                                                                                                 arg0_2_1Dcon_main1_3_r,
                                                                                                 arg0_2_1Dcon_main1_2_r,
                                                                                                 arg0_2_1Dcon_main1_1_r}));
  assign arg0_2_1Dcon_main1_r = (& arg0_2_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_2_1Dcon_main1_emitted <= (arg0_2_1Dcon_main1_r ? 4'd0 :
                                     arg0_2_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_1Dcon_main1_1I#,Int) > [(x1ajF_destruct,Int#)] */
  assign x1ajF_destruct_d = {\arg0_2_1Dcon_main1_1I#_d [32:1],
                             \arg0_2_1Dcon_main1_1I#_d [0]};
  assign \arg0_2_1Dcon_main1_1I#_r  = x1ajF_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_1Dcon_main1_2,Int) (arg0_2_1Dcon_main1_1,Int) > [(arg0_2_1Dcon_main1_1I#,Int)] */
  assign \arg0_2_1Dcon_main1_1I#_d  = {arg0_2_1Dcon_main1_1_d[32:1],
                                       (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0])};
  assign arg0_2_1Dcon_main1_1_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  assign arg0_2_1Dcon_main1_2_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_2_1Dcon_main1_3,Int) (arg0_2_2Dcon_main1,Go) > [(arg0_2_1Dcon_main1_3I#,Go)] */
  assign \arg0_2_1Dcon_main1_3I#_d  = (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]);
  assign arg0_2_2Dcon_main1_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  assign arg0_2_1Dcon_main1_3_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  
  /* fork (Ty Go) : (arg0_2_1Dcon_main1_3I#,Go) > [(arg0_2_1Dcon_main1_3I#_1,Go),
                                              (arg0_2_1Dcon_main1_3I#_2,Go),
                                              (arg0_2_1Dcon_main1_3I#_3,Go)] */
  logic [2:0] \arg0_2_1Dcon_main1_3I#_emitted ;
  logic [2:0] \arg0_2_1Dcon_main1_3I#_done ;
  assign \arg0_2_1Dcon_main1_3I#_1_d  = (\arg0_2_1Dcon_main1_3I#_d [0] && (! \arg0_2_1Dcon_main1_3I#_emitted [0]));
  assign \arg0_2_1Dcon_main1_3I#_2_d  = (\arg0_2_1Dcon_main1_3I#_d [0] && (! \arg0_2_1Dcon_main1_3I#_emitted [1]));
  assign \arg0_2_1Dcon_main1_3I#_3_d  = (\arg0_2_1Dcon_main1_3I#_d [0] && (! \arg0_2_1Dcon_main1_3I#_emitted [2]));
  assign \arg0_2_1Dcon_main1_3I#_done  = (\arg0_2_1Dcon_main1_3I#_emitted  | ({\arg0_2_1Dcon_main1_3I#_3_d [0],
                                                                               \arg0_2_1Dcon_main1_3I#_2_d [0],
                                                                               \arg0_2_1Dcon_main1_3I#_1_d [0]} & {\arg0_2_1Dcon_main1_3I#_3_r ,
                                                                                                                   \arg0_2_1Dcon_main1_3I#_2_r ,
                                                                                                                   \arg0_2_1Dcon_main1_3I#_1_r }));
  assign \arg0_2_1Dcon_main1_3I#_r  = (& \arg0_2_1Dcon_main1_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_emitted  <= 3'd0;
    else
      \arg0_2_1Dcon_main1_3I#_emitted  <= (\arg0_2_1Dcon_main1_3I#_r  ? 3'd0 :
                                           \arg0_2_1Dcon_main1_3I#_done );
  
  /* buf (Ty Go) : (arg0_2_1Dcon_main1_3I#_1,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_2_1Dcon_main1_3I#_1_bufchan_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_bufchan_r ;
  assign \arg0_2_1Dcon_main1_3I#_1_r  = ((! \arg0_2_1Dcon_main1_3I#_1_bufchan_d [0]) || \arg0_2_1Dcon_main1_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_2_1Dcon_main1_3I#_1_r )
        \arg0_2_1Dcon_main1_3I#_1_bufchan_d  <= \arg0_2_1Dcon_main1_3I#_1_d ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_bufchan_buf ;
  assign \arg0_2_1Dcon_main1_3I#_1_bufchan_r  = (! \arg0_2_1Dcon_main1_3I#_1_bufchan_buf [0]);
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_2_1Dcon_main1_3I#_1_bufchan_buf [0] ? \arg0_2_1Dcon_main1_3I#_1_bufchan_buf  :
                                                \arg0_2_1Dcon_main1_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_2_1Dcon_main1_3I#_1_argbuf_r  && \arg0_2_1Dcon_main1_3I#_1_bufchan_buf [0]))
        \arg0_2_1Dcon_main1_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_2_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_2_1Dcon_main1_3I#_1_bufchan_buf [0])))
        \arg0_2_1Dcon_main1_3I#_1_bufchan_buf  <= \arg0_2_1Dcon_main1_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf_0,Int#) */
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_0_d  = {32'd0,
                                                  \arg0_2_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_r  = \arg0_2_1Dcon_main1_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_2_1Dcon_main1_3I#_1_argbuf_0,Int#) (x1ajF_destruct,Int#) > (lizzieLet2_1wild1XF_1_Eq,Bool) */
  assign lizzieLet2_1wild1XF_1_Eq_d = {(\arg0_2_1Dcon_main1_3I#_1_argbuf_0_d [32:1] == x1ajF_destruct_d[32:1]),
                                       (\arg0_2_1Dcon_main1_3I#_1_argbuf_0_d [0] && x1ajF_destruct_d[0])};
  assign {\arg0_2_1Dcon_main1_3I#_1_argbuf_0_r ,
          x1ajF_destruct_r} = {2 {(lizzieLet2_1wild1XF_1_Eq_r && lizzieLet2_1wild1XF_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_2_1Dcon_main1_3I#_2,Go) > (arg0_2_1Dcon_main1_3I#_2_argbuf,Go) */
  Go_t \arg0_2_1Dcon_main1_3I#_2_bufchan_d ;
  logic \arg0_2_1Dcon_main1_3I#_2_bufchan_r ;
  assign \arg0_2_1Dcon_main1_3I#_2_r  = ((! \arg0_2_1Dcon_main1_3I#_2_bufchan_d [0]) || \arg0_2_1Dcon_main1_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_2_1Dcon_main1_3I#_2_r )
        \arg0_2_1Dcon_main1_3I#_2_bufchan_d  <= \arg0_2_1Dcon_main1_3I#_2_d ;
  Go_t \arg0_2_1Dcon_main1_3I#_2_bufchan_buf ;
  assign \arg0_2_1Dcon_main1_3I#_2_bufchan_r  = (! \arg0_2_1Dcon_main1_3I#_2_bufchan_buf [0]);
  assign \arg0_2_1Dcon_main1_3I#_2_argbuf_d  = (\arg0_2_1Dcon_main1_3I#_2_bufchan_buf [0] ? \arg0_2_1Dcon_main1_3I#_2_bufchan_buf  :
                                                \arg0_2_1Dcon_main1_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_2_1Dcon_main1_3I#_2_argbuf_r  && \arg0_2_1Dcon_main1_3I#_2_bufchan_buf [0]))
        \arg0_2_1Dcon_main1_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_2_1Dcon_main1_3I#_2_argbuf_r ) && (! \arg0_2_1Dcon_main1_3I#_2_bufchan_buf [0])))
        \arg0_2_1Dcon_main1_3I#_2_bufchan_buf  <= \arg0_2_1Dcon_main1_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_2_1Dcon_main1_3I#_2_argbuf,Go),
                            (lizzieLet3_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_2_1Dcon_main1_3I#_2_argbuf_d [0],
                                                             lizzieLet3_1_argbuf_d[0]}), \arg0_2_1Dcon_main1_3I#_2_argbuf_d , lizzieLet3_1_argbuf_d);
  assign {\arg0_2_1Dcon_main1_3I#_2_argbuf_r ,
          lizzieLet3_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_2_1Dcon_main1_4,Int) [(lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux,MyBool)] > (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux,MyBool) */
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d = {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d[1:1],
                                                                             (arg0_2_1Dcon_main1_4_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d[0])};
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_r = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_r && (arg0_2_1Dcon_main1_4_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d[0]));
  assign arg0_2_1Dcon_main1_4_r = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_r && (arg0_2_1Dcon_main1_4_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10,Go) > [(arg0_2_2Dcon_main1,Go)] */
  assign arg0_2_2Dcon_main1_d = (arg0_2_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d[0]));
  assign arg0_2_2_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_10_d[0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_2_3,MyDTInt_Bool) [(lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux,MyBool)] > (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux,MyBool) */
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_d = {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d[1:1],
                                                                                 (arg0_2_3_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d[0])};
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_r = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_r && (arg0_2_3_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d[0]));
  assign arg0_2_3_r = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_r && (arg0_2_3_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_d[0]));
  
  /* mux (Ty MyDTBool_Bool,
     Ty MyBool) : (arg0_3,MyDTBool_Bool) [(arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux,MyBool)] > (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux,MyBool) */
  assign arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_d = {arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d[1:1],
                                                                                         (arg0_3_d[0] && arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d[0])};
  assign arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_r = (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d[0]));
  assign arg0_3_r = (arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main2_1MyFalse_1MyTruearg0_1Dcon_main2_1MyTrue_1MyFalse_mux_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int) > [(arg0_4_1Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_4_1Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[32:1],
                                          (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r = (\arg0_4_1Dcon_$fNumInt_$c+_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  assign arg0_4_1_r = (\arg0_4_1Dcon_$fNumInt_$c+_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_4_2Dcon_$fNumInt_$c+,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                          (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_4_2Dcon_$fNumInt_$c+_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_4_2_r = (\arg0_4_2Dcon_$fNumInt_$c+_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_1,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_2,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_3,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c+_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_done ;
  assign \arg0_4_2Dcon_$fNumInt_$c+_1_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_2_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_4_d  = {\arg0_4_2Dcon_$fNumInt_$c+_d [32:1],
                                            (\arg0_4_2Dcon_$fNumInt_$c+_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_done  = (\arg0_4_2Dcon_$fNumInt_$c+_emitted  | ({\arg0_4_2Dcon_$fNumInt_$c+_4_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_3_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_2_d [0],
                                                                                     \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$c+_4_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_3_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_2_r ,
                                                                                                                            \arg0_4_2Dcon_$fNumInt_$c+_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$c+_r  = (& \arg0_4_2Dcon_$fNumInt_$c+_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_4_2Dcon_$fNumInt_$c+_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$c+_emitted  <= (\arg0_4_2Dcon_$fNumInt_$c+_r  ? 4'd0 :
                                              \arg0_4_2Dcon_$fNumInt_$c+_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c+_1I#,Int) > [(xa1lV_destruct,Int#)] */
  assign xa1lV_destruct_d = {\arg0_4_2Dcon_$fNumInt_$c+_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$c+_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$c+_1I#_r  = xa1lV_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_2,Int) (arg0_4_2Dcon_$fNumInt_$c+_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$c+_1_d [32:1],
                                              (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$c+_1_r  = (\arg0_4_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_2_r  = (\arg0_4_2Dcon_$fNumInt_$c+_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3,Int) (arg0_4_1Dcon_$fNumInt_$c+,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_d  = {\arg0_4_1Dcon_$fNumInt_$c+_d [32:1],
                                              (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0])};
  assign \arg0_4_1Dcon_$fNumInt_$c+_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3_d [0] && \arg0_4_1Dcon_$fNumInt_$c+_d [0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_1,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_2,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_3,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c+_3I#_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$c+_3I#_done ;
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$c+_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_done  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  | ({\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_r  = (& \arg0_4_2Dcon_$fNumInt_$c+_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$c+_3I#_emitted  <= (\arg0_4_2Dcon_$fNumInt_$c+_3I#_r  ? 4'd0 :
                                                  \arg0_4_2Dcon_$fNumInt_$c+_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#,Int) > [(ya1lW_destruct,Int#)] */
  assign ya1lW_destruct_d = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  = ya1lW_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_2,Int) (arg0_4_2Dcon_$fNumInt_$c+_3I#_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_2_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$c+_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_3,Int) (xa1lV_destruct,Int#) > [(arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#,Int#)] */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d  = {xa1lV_destruct_d[32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0])};
  assign xa1lV_destruct_r = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3_r  = (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3_d [0] && xa1lV_destruct_d[0]));
  
  /* op_add (Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#,Int#) (ya1lW_destruct,Int#) > (arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#) */
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d  = {(\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d [32:1] + ya1lW_destruct_d[32:1]),
                                                                 (\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_d [0] && ya1lW_destruct_d[0])};
  assign {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_r ,
          ya1lW_destruct_r} = {2 {(\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r  && \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32,Int#)] > (es_0_2_1I#,Int) */
  assign \es_0_2_1I#_d  = \I#_dc ((& {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d [0]}), \arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_d );
  assign {\arg0_4_2Dcon_$fNumInt_$c+_3I#_3I#_1ya1lW_1_Add32_r } = {1 {(\es_0_2_1I#_r  && \es_0_2_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_3I#_4,Int) [(es_0_2_1I#,Int)] > (es_0_2_1I#_mux,Int) */
  assign \es_0_2_1I#_mux_d  = {\es_0_2_1I#_d [32:1],
                               (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0])};
  assign \es_0_2_1I#_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_3I#_4_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c+_4,Int) [(es_0_2_1I#_mux,Int)] > (es_0_2_1I#_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_d  = {\es_0_2_1I#_mux_d [32:1],
                                   (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0])};
  assign \es_0_2_1I#_mux_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$c+_4_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$c+_4_d [0] && \es_0_2_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_4_3,MyDTInt_Int_Int) [(es_0_2_1I#_mux_mux,Int)] > (es_0_2_1I#_mux_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_mux_d  = {\es_0_2_1I#_mux_mux_d [32:1],
                                       (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0])};
  assign \es_0_2_1I#_mux_mux_r  = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  assign arg0_4_3_r = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet4_1,MyBool),
                                                    (lizzieLet4_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet4_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet4_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet4_2_d[0],
                                                                       lizzieLet4_1_d[0]} & {lizzieLet4_2_r,
                                                                                             lizzieLet4_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int,
          Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) : (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) > [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11,Go),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                             (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0,Pointer_CT$wmAdd_Int)] */
  logic [4:0] call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted;
  logic [4:0] call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done;
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[0]));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[1]));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[16:1],
                                                                                                                           (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[2]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[32:17],
                                                                                                                           (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[3]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[48:33],
                                                                                                                        (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0] && (! call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted[4]))};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done = (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted | ({call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d[0],
                                                                                                                                                                                                                                             call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d[0]} & {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r,
                                                                                                                                                                                                                                                                                                                                                                 call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_r,
                                                                                                                                                                                                                                                                                                                                                                 call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_r,
                                                                                                                                                                                                                                                                                                                                                                 call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_r,
                                                                                                                                                                                                                                                                                                                                                                 call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_r}));
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r = (& call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted <= 5'd0;
    else
      call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_emitted <= (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r ? 5'd0 :
                                                                                                                          call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wmAdd_Int_goConst,Go) > (call_$wmAdd_Int_initBufi,Go) */
  Go_t call_$wmAdd_Int_goConst_buf;
  assign call_$wmAdd_Int_goConst_r = (! call_$wmAdd_Int_goConst_buf[0]);
  assign call_$wmAdd_Int_initBufi_d = (call_$wmAdd_Int_goConst_buf[0] ? call_$wmAdd_Int_goConst_buf :
                                       call_$wmAdd_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wmAdd_Int_initBufi_r && call_$wmAdd_Int_goConst_buf[0]))
        call_$wmAdd_Int_goConst_buf <= 1'd0;
      else if (((! call_$wmAdd_Int_initBufi_r) && (! call_$wmAdd_Int_goConst_buf[0])))
        call_$wmAdd_Int_goConst_buf <= call_$wmAdd_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wmAdd_Int_goMux1,Go),
                           (lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf,Go),
                           (lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf,Go),
                           (lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf,Go),
                           (lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] call_$wmAdd_Int_goMux1_select_d;
  assign call_$wmAdd_Int_goMux1_select_d = ((| call_$wmAdd_Int_goMux1_select_q) ? call_$wmAdd_Int_goMux1_select_q :
                                            (call_$wmAdd_Int_goMux1_d[0] ? 5'd1 :
                                             (lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] call_$wmAdd_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goMux1_select_q <= 5'd0;
    else
      call_$wmAdd_Int_goMux1_select_q <= (call_$wmAdd_Int_goMux1_done ? 5'd0 :
                                          call_$wmAdd_Int_goMux1_select_d);
  logic [1:0] call_$wmAdd_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wmAdd_Int_goMux1_emit_q <= (call_$wmAdd_Int_goMux1_done ? 2'd0 :
                                        call_$wmAdd_Int_goMux1_emit_d);
  logic [1:0] call_$wmAdd_Int_goMux1_emit_d;
  assign call_$wmAdd_Int_goMux1_emit_d = (call_$wmAdd_Int_goMux1_emit_q | ({go_11_goMux_choice_d[0],
                                                                            go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                      go_11_goMux_data_r}));
  logic call_$wmAdd_Int_goMux1_done;
  assign call_$wmAdd_Int_goMux1_done = (& call_$wmAdd_Int_goMux1_emit_d);
  assign {lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_r,
          lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_r,
          lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_r,
          lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_r,
          call_$wmAdd_Int_goMux1_r} = (call_$wmAdd_Int_goMux1_done ? call_$wmAdd_Int_goMux1_select_d :
                                       5'd0);
  assign go_11_goMux_data_d = ((call_$wmAdd_Int_goMux1_select_d[0] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? call_$wmAdd_Int_goMux1_d :
                               ((call_$wmAdd_Int_goMux1_select_d[1] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_d :
                                ((call_$wmAdd_Int_goMux1_select_d[2] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_d :
                                 ((call_$wmAdd_Int_goMux1_select_d[3] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_d :
                                  ((call_$wmAdd_Int_goMux1_select_d[4] && (! call_$wmAdd_Int_goMux1_emit_q[0])) ? lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((call_$wmAdd_Int_goMux1_select_d[0] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wmAdd_Int_goMux1_select_d[1] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wmAdd_Int_goMux1_select_d[2] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wmAdd_Int_goMux1_select_d[3] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wmAdd_Int_goMux1_select_d[4] && (! call_$wmAdd_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wmAdd_Int_initBuf,Go) > [(call_$wmAdd_Int_unlockFork1,Go),
                                               (call_$wmAdd_Int_unlockFork2,Go),
                                               (call_$wmAdd_Int_unlockFork3,Go),
                                               (call_$wmAdd_Int_unlockFork4,Go),
                                               (call_$wmAdd_Int_unlockFork5,Go)] */
  logic [4:0] call_$wmAdd_Int_initBuf_emitted;
  logic [4:0] call_$wmAdd_Int_initBuf_done;
  assign call_$wmAdd_Int_unlockFork1_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[0]));
  assign call_$wmAdd_Int_unlockFork2_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[1]));
  assign call_$wmAdd_Int_unlockFork3_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[2]));
  assign call_$wmAdd_Int_unlockFork4_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[3]));
  assign call_$wmAdd_Int_unlockFork5_d = (call_$wmAdd_Int_initBuf_d[0] && (! call_$wmAdd_Int_initBuf_emitted[4]));
  assign call_$wmAdd_Int_initBuf_done = (call_$wmAdd_Int_initBuf_emitted | ({call_$wmAdd_Int_unlockFork5_d[0],
                                                                             call_$wmAdd_Int_unlockFork4_d[0],
                                                                             call_$wmAdd_Int_unlockFork3_d[0],
                                                                             call_$wmAdd_Int_unlockFork2_d[0],
                                                                             call_$wmAdd_Int_unlockFork1_d[0]} & {call_$wmAdd_Int_unlockFork5_r,
                                                                                                                  call_$wmAdd_Int_unlockFork4_r,
                                                                                                                  call_$wmAdd_Int_unlockFork3_r,
                                                                                                                  call_$wmAdd_Int_unlockFork2_r,
                                                                                                                  call_$wmAdd_Int_unlockFork1_r}));
  assign call_$wmAdd_Int_initBuf_r = (& call_$wmAdd_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_initBuf_emitted <= 5'd0;
    else
      call_$wmAdd_Int_initBuf_emitted <= (call_$wmAdd_Int_initBuf_r ? 5'd0 :
                                          call_$wmAdd_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wmAdd_Int_initBufi,Go) > (call_$wmAdd_Int_initBuf,Go) */
  assign call_$wmAdd_Int_initBufi_r = ((! call_$wmAdd_Int_initBuf_d[0]) || call_$wmAdd_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wmAdd_Int_initBufi_r)
        call_$wmAdd_Int_initBuf_d <= call_$wmAdd_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wmAdd_Int_unlockFork1,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11,Go)] > (call_$wmAdd_Int_goMux1,Go) */
  assign call_$wmAdd_Int_goMux1_d = (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d[0]);
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_r = (call_$wmAdd_Int_goMux1_r && (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d[0]));
  assign call_$wmAdd_Int_unlockFork1_r = (call_$wmAdd_Int_goMux1_r && (call_$wmAdd_Int_unlockFork1_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intgo_11_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_$wmAdd_Int_unlockFork2,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1,MyDTInt_Int_Int)] > (call_$wmAdd_Int_goMux2,MyDTInt_Int_Int) */
  assign call_$wmAdd_Int_goMux2_d = (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d[0]);
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_r = (call_$wmAdd_Int_goMux2_r && (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d[0]));
  assign call_$wmAdd_Int_unlockFork2_r = (call_$wmAdd_Int_goMux2_r && (call_$wmAdd_Int_unlockFork2_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_IntwslR_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wmAdd_Int_unlockFork3,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1,Pointer_QTree_Int)] > (call_$wmAdd_Int_goMux3,Pointer_QTree_Int) */
  assign call_$wmAdd_Int_goMux3_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d[16:1],
                                     (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_r = (call_$wmAdd_Int_goMux3_r && (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d[0]));
  assign call_$wmAdd_Int_unlockFork3_r = (call_$wmAdd_Int_goMux3_r && (call_$wmAdd_Int_unlockFork3_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw1slS_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wmAdd_Int_unlockFork4,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1,Pointer_QTree_Int)] > (call_$wmAdd_Int_goMux4,Pointer_QTree_Int) */
  assign call_$wmAdd_Int_goMux4_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d[16:1],
                                     (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_r = (call_$wmAdd_Int_goMux4_r && (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d[0]));
  assign call_$wmAdd_Int_unlockFork4_r = (call_$wmAdd_Int_goMux4_r && (call_$wmAdd_Int_unlockFork4_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intw2slT_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wmAdd_Int) : (call_$wmAdd_Int_unlockFork5,Go) [(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0,Pointer_CT$wmAdd_Int)] > (call_$wmAdd_Int_goMux5,Pointer_CT$wmAdd_Int) */
  assign call_$wmAdd_Int_goMux5_d = {call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[16:1],
                                     (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0])};
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_r = (call_$wmAdd_Int_goMux5_r && (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0]));
  assign call_$wmAdd_Int_unlockFork5_r = (call_$wmAdd_Int_goMux5_r && (call_$wmAdd_Int_unlockFork5_d[0] && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) : (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) > [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12,Go),
                                                                                                                                                                          (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1,Pointer_QTree_Bool),
                                                                                                                                                                          (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1,Pointer_CT$wnnz)] */
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted;
  logic [2:0] call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done;
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d = (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[0]));
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[16:1],
                                                                           (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[1]))};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[32:17],
                                                                           (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0] && (! call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted[2]))};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done = (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted | ({call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d[0],
                                                                                                                                               call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d[0],
                                                                                                                                               call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d[0]} & {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_r,
                                                                                                                                                                                                                    call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_r,
                                                                                                                                                                                                                    call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_r}));
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r = (& call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted <= 3'd0;
    else
      call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_emitted <= (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r ? 3'd0 :
                                                                           call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_goConst,Go) > (call_$wnnz_initBufi,Go) */
  Go_t call_$wnnz_goConst_buf;
  assign call_$wnnz_goConst_r = (! call_$wnnz_goConst_buf[0]);
  assign call_$wnnz_initBufi_d = (call_$wnnz_goConst_buf[0] ? call_$wnnz_goConst_buf :
                                  call_$wnnz_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_initBufi_r && call_$wnnz_goConst_buf[0]))
        call_$wnnz_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_initBufi_r) && (! call_$wnnz_goConst_buf[0])))
        call_$wnnz_goConst_buf <= call_$wnnz_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_goMux1,Go),
                           (lizzieLet29_3Lcall_$wnnz3_1_argbuf,Go),
                           (lizzieLet29_3Lcall_$wnnz2_1_argbuf,Go),
                           (lizzieLet29_3Lcall_$wnnz1_1_argbuf,Go),
                           (lizzieLet15_3QNode_Bool_1_argbuf,Go)] > (go_12_goMux_choice,C5) (go_12_goMux_data,Go) */
  logic [4:0] call_$wnnz_goMux1_select_d;
  assign call_$wnnz_goMux1_select_d = ((| call_$wnnz_goMux1_select_q) ? call_$wnnz_goMux1_select_q :
                                       (call_$wnnz_goMux1_d[0] ? 5'd1 :
                                        (lizzieLet29_3Lcall_$wnnz3_1_argbuf_d[0] ? 5'd2 :
                                         (lizzieLet29_3Lcall_$wnnz2_1_argbuf_d[0] ? 5'd4 :
                                          (lizzieLet29_3Lcall_$wnnz1_1_argbuf_d[0] ? 5'd8 :
                                           (lizzieLet15_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                            5'd0))))));
  logic [4:0] call_$wnnz_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_goMux1_select_q <= (call_$wnnz_goMux1_done ? 5'd0 :
                                     call_$wnnz_goMux1_select_d);
  logic [1:0] call_$wnnz_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_goMux1_emit_q <= (call_$wnnz_goMux1_done ? 2'd0 :
                                   call_$wnnz_goMux1_emit_d);
  logic [1:0] call_$wnnz_goMux1_emit_d;
  assign call_$wnnz_goMux1_emit_d = (call_$wnnz_goMux1_emit_q | ({go_12_goMux_choice_d[0],
                                                                  go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                            go_12_goMux_data_r}));
  logic call_$wnnz_goMux1_done;
  assign call_$wnnz_goMux1_done = (& call_$wnnz_goMux1_emit_d);
  assign {lizzieLet15_3QNode_Bool_1_argbuf_r,
          lizzieLet29_3Lcall_$wnnz1_1_argbuf_r,
          lizzieLet29_3Lcall_$wnnz2_1_argbuf_r,
          lizzieLet29_3Lcall_$wnnz3_1_argbuf_r,
          call_$wnnz_goMux1_r} = (call_$wnnz_goMux1_done ? call_$wnnz_goMux1_select_d :
                                  5'd0);
  assign go_12_goMux_data_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[0])) ? call_$wnnz_goMux1_d :
                               ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_$wnnz3_1_argbuf_d :
                                ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_$wnnz2_1_argbuf_d :
                                 ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet29_3Lcall_$wnnz1_1_argbuf_d :
                                  ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[0])) ? lizzieLet15_3QNode_Bool_1_argbuf_d :
                                   1'd0)))));
  assign go_12_goMux_choice_d = ((call_$wnnz_goMux1_select_d[0] && (! call_$wnnz_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wnnz_goMux1_select_d[1] && (! call_$wnnz_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wnnz_goMux1_select_d[2] && (! call_$wnnz_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wnnz_goMux1_select_d[3] && (! call_$wnnz_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wnnz_goMux1_select_d[4] && (! call_$wnnz_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_initBuf,Go) > [(call_$wnnz_unlockFork1,Go),
                                          (call_$wnnz_unlockFork2,Go),
                                          (call_$wnnz_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_initBuf_emitted;
  logic [2:0] call_$wnnz_initBuf_done;
  assign call_$wnnz_unlockFork1_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[0]));
  assign call_$wnnz_unlockFork2_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[1]));
  assign call_$wnnz_unlockFork3_d = (call_$wnnz_initBuf_d[0] && (! call_$wnnz_initBuf_emitted[2]));
  assign call_$wnnz_initBuf_done = (call_$wnnz_initBuf_emitted | ({call_$wnnz_unlockFork3_d[0],
                                                                   call_$wnnz_unlockFork2_d[0],
                                                                   call_$wnnz_unlockFork1_d[0]} & {call_$wnnz_unlockFork3_r,
                                                                                                   call_$wnnz_unlockFork2_r,
                                                                                                   call_$wnnz_unlockFork1_r}));
  assign call_$wnnz_initBuf_r = (& call_$wnnz_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_initBuf_emitted <= (call_$wnnz_initBuf_r ? 3'd0 :
                                     call_$wnnz_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_initBufi,Go) > (call_$wnnz_initBuf,Go) */
  assign call_$wnnz_initBufi_r = ((! call_$wnnz_initBuf_d[0]) || call_$wnnz_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_initBufi_r)
        call_$wnnz_initBuf_d <= call_$wnnz_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_unlockFork1,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12,Go)] > (call_$wnnz_goMux1,Go) */
  assign call_$wnnz_goMux1_d = (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d[0]);
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d[0]));
  assign call_$wnnz_unlockFork1_r = (call_$wnnz_goMux1_r && (call_$wnnz_unlockFork1_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzgo_12_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_$wnnz_unlockFork2,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1,Pointer_QTree_Bool)] > (call_$wnnz_goMux2,Pointer_QTree_Bool) */
  assign call_$wnnz_goMux2_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d[16:1],
                                (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d[0]));
  assign call_$wnnz_unlockFork2_r = (call_$wnnz_goMux2_r && (call_$wnnz_unlockFork2_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzwslW_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz) : (call_$wnnz_unlockFork3,Go) [(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1,Pointer_CT$wnnz)] > (call_$wnnz_goMux3,Pointer_CT$wnnz) */
  assign call_$wnnz_goMux3_d = {call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d[16:1],
                                (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d[0])};
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d[0]));
  assign call_$wnnz_unlockFork3_r = (call_$wnnz_goMux3_r && (call_$wnnz_unlockFork3_d[0] && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnzsc_0_1_d[0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool) : (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1,TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool) > [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13,Go),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2,Pointer_CTmain_map'_Int_Bool)] */
  logic [4:0] \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted ;
  logic [4:0] \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_done ;
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d  = (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0] && (! \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted [0]));
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d  = (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0] && (! \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted [1]));
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d  = (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0] && (! \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted [2]));
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d  = {\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [16:1],
                                                                                                                                   (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0] && (! \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted [3]))};
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d  = {\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [32:17],
                                                                                                                                     (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0] && (! \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted [4]))};
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_done  = (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted  | ({\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d [0]} & {\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                                  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_r ,
                                                                                                                                                                                                                                                                                                                                                                                                  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_r ,
                                                                                                                                                                                                                                                                                                                                                                                                  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_r ,
                                                                                                                                                                                                                                                                                                                                                                                                  \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_r }));
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_r  = (& \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted  <= 5'd0;
    else
      \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_emitted  <= (\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_r  ? 5'd0 :
                                                                                                                                     \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_done );
  
  /* rbuf (Ty Go) : (call_main_map'_Int_Bool_goConst,Go) > (call_main_map'_Int_Bool_initBufi,Go) */
  Go_t \call_main_map'_Int_Bool_goConst_buf ;
  assign \call_main_map'_Int_Bool_goConst_r  = (! \call_main_map'_Int_Bool_goConst_buf [0]);
  assign \call_main_map'_Int_Bool_initBufi_d  = (\call_main_map'_Int_Bool_goConst_buf [0] ? \call_main_map'_Int_Bool_goConst_buf  :
                                                 \call_main_map'_Int_Bool_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_main_map'_Int_Bool_goConst_buf  <= 1'd0;
    else
      if ((\call_main_map'_Int_Bool_initBufi_r  && \call_main_map'_Int_Bool_goConst_buf [0]))
        \call_main_map'_Int_Bool_goConst_buf  <= 1'd0;
      else if (((! \call_main_map'_Int_Bool_initBufi_r ) && (! \call_main_map'_Int_Bool_goConst_buf [0])))
        \call_main_map'_Int_Bool_goConst_buf  <= \call_main_map'_Int_Bool_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_map'_Int_Bool_goMux1,Go),
                           (lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf,Go),
                           (lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf,Go),
                           (lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf,Go),
                           (lizzieLet17_4QNode_Int_1_argbuf,Go)] > (go_13_goMux_choice,C5) (go_13_goMux_data,Go) */
  logic [4:0] \call_main_map'_Int_Bool_goMux1_select_d ;
  assign \call_main_map'_Int_Bool_goMux1_select_d  = ((| \call_main_map'_Int_Bool_goMux1_select_q ) ? \call_main_map'_Int_Bool_goMux1_select_q  :
                                                      (\call_main_map'_Int_Bool_goMux1_d [0] ? 5'd1 :
                                                       (\lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_d [0] ? 5'd2 :
                                                        (\lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_d [0] ? 5'd4 :
                                                         (\lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_d [0] ? 5'd8 :
                                                          (lizzieLet17_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                           5'd0))))));
  logic [4:0] \call_main_map'_Int_Bool_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Bool_goMux1_select_q  <= 5'd0;
    else
      \call_main_map'_Int_Bool_goMux1_select_q  <= (\call_main_map'_Int_Bool_goMux1_done  ? 5'd0 :
                                                    \call_main_map'_Int_Bool_goMux1_select_d );
  logic [1:0] \call_main_map'_Int_Bool_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Bool_goMux1_emit_q  <= 2'd0;
    else
      \call_main_map'_Int_Bool_goMux1_emit_q  <= (\call_main_map'_Int_Bool_goMux1_done  ? 2'd0 :
                                                  \call_main_map'_Int_Bool_goMux1_emit_d );
  logic [1:0] \call_main_map'_Int_Bool_goMux1_emit_d ;
  assign \call_main_map'_Int_Bool_goMux1_emit_d  = (\call_main_map'_Int_Bool_goMux1_emit_q  | ({go_13_goMux_choice_d[0],
                                                                                                go_13_goMux_data_d[0]} & {go_13_goMux_choice_r,
                                                                                                                          go_13_goMux_data_r}));
  logic \call_main_map'_Int_Bool_goMux1_done ;
  assign \call_main_map'_Int_Bool_goMux1_done  = (& \call_main_map'_Int_Bool_goMux1_emit_d );
  assign {lizzieLet17_4QNode_Int_1_argbuf_r,
          \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_r ,
          \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_r ,
          \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_r ,
          \call_main_map'_Int_Bool_goMux1_r } = (\call_main_map'_Int_Bool_goMux1_done  ? \call_main_map'_Int_Bool_goMux1_select_d  :
                                                 5'd0);
  assign go_13_goMux_data_d = ((\call_main_map'_Int_Bool_goMux1_select_d [0] && (! \call_main_map'_Int_Bool_goMux1_emit_q [0])) ? \call_main_map'_Int_Bool_goMux1_d  :
                               ((\call_main_map'_Int_Bool_goMux1_select_d [1] && (! \call_main_map'_Int_Bool_goMux1_emit_q [0])) ? \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_d  :
                                ((\call_main_map'_Int_Bool_goMux1_select_d [2] && (! \call_main_map'_Int_Bool_goMux1_emit_q [0])) ? \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_d  :
                                 ((\call_main_map'_Int_Bool_goMux1_select_d [3] && (! \call_main_map'_Int_Bool_goMux1_emit_q [0])) ? \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_d  :
                                  ((\call_main_map'_Int_Bool_goMux1_select_d [4] && (! \call_main_map'_Int_Bool_goMux1_emit_q [0])) ? lizzieLet17_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_13_goMux_choice_d = ((\call_main_map'_Int_Bool_goMux1_select_d [0] && (! \call_main_map'_Int_Bool_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_main_map'_Int_Bool_goMux1_select_d [1] && (! \call_main_map'_Int_Bool_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_main_map'_Int_Bool_goMux1_select_d [2] && (! \call_main_map'_Int_Bool_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_main_map'_Int_Bool_goMux1_select_d [3] && (! \call_main_map'_Int_Bool_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_main_map'_Int_Bool_goMux1_select_d [4] && (! \call_main_map'_Int_Bool_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_map'_Int_Bool_initBuf,Go) > [(call_main_map'_Int_Bool_unlockFork1,Go),
                                                       (call_main_map'_Int_Bool_unlockFork2,Go),
                                                       (call_main_map'_Int_Bool_unlockFork3,Go),
                                                       (call_main_map'_Int_Bool_unlockFork4,Go),
                                                       (call_main_map'_Int_Bool_unlockFork5,Go)] */
  logic [4:0] \call_main_map'_Int_Bool_initBuf_emitted ;
  logic [4:0] \call_main_map'_Int_Bool_initBuf_done ;
  assign \call_main_map'_Int_Bool_unlockFork1_d  = (\call_main_map'_Int_Bool_initBuf_d [0] && (! \call_main_map'_Int_Bool_initBuf_emitted [0]));
  assign \call_main_map'_Int_Bool_unlockFork2_d  = (\call_main_map'_Int_Bool_initBuf_d [0] && (! \call_main_map'_Int_Bool_initBuf_emitted [1]));
  assign \call_main_map'_Int_Bool_unlockFork3_d  = (\call_main_map'_Int_Bool_initBuf_d [0] && (! \call_main_map'_Int_Bool_initBuf_emitted [2]));
  assign \call_main_map'_Int_Bool_unlockFork4_d  = (\call_main_map'_Int_Bool_initBuf_d [0] && (! \call_main_map'_Int_Bool_initBuf_emitted [3]));
  assign \call_main_map'_Int_Bool_unlockFork5_d  = (\call_main_map'_Int_Bool_initBuf_d [0] && (! \call_main_map'_Int_Bool_initBuf_emitted [4]));
  assign \call_main_map'_Int_Bool_initBuf_done  = (\call_main_map'_Int_Bool_initBuf_emitted  | ({\call_main_map'_Int_Bool_unlockFork5_d [0],
                                                                                                 \call_main_map'_Int_Bool_unlockFork4_d [0],
                                                                                                 \call_main_map'_Int_Bool_unlockFork3_d [0],
                                                                                                 \call_main_map'_Int_Bool_unlockFork2_d [0],
                                                                                                 \call_main_map'_Int_Bool_unlockFork1_d [0]} & {\call_main_map'_Int_Bool_unlockFork5_r ,
                                                                                                                                                \call_main_map'_Int_Bool_unlockFork4_r ,
                                                                                                                                                \call_main_map'_Int_Bool_unlockFork3_r ,
                                                                                                                                                \call_main_map'_Int_Bool_unlockFork2_r ,
                                                                                                                                                \call_main_map'_Int_Bool_unlockFork1_r }));
  assign \call_main_map'_Int_Bool_initBuf_r  = (& \call_main_map'_Int_Bool_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Bool_initBuf_emitted  <= 5'd0;
    else
      \call_main_map'_Int_Bool_initBuf_emitted  <= (\call_main_map'_Int_Bool_initBuf_r  ? 5'd0 :
                                                    \call_main_map'_Int_Bool_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_map'_Int_Bool_initBufi,Go) > (call_main_map'_Int_Bool_initBuf,Go) */
  assign \call_main_map'_Int_Bool_initBufi_r  = ((! \call_main_map'_Int_Bool_initBuf_d [0]) || \call_main_map'_Int_Bool_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Int_Bool_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_main_map'_Int_Bool_initBufi_r )
        \call_main_map'_Int_Bool_initBuf_d  <= \call_main_map'_Int_Bool_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_map'_Int_Bool_unlockFork1,Go) [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13,Go)] > (call_main_map'_Int_Bool_goMux1,Go) */
  assign \call_main_map'_Int_Bool_goMux1_d  = (\call_main_map'_Int_Bool_unlockFork1_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d [0]);
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_r  = (\call_main_map'_Int_Bool_goMux1_r  && (\call_main_map'_Int_Bool_unlockFork1_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d [0]));
  assign \call_main_map'_Int_Bool_unlockFork1_r  = (\call_main_map'_Int_Bool_goMux1_r  && (\call_main_map'_Int_Bool_unlockFork1_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolgo_13_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool) : (call_main_map'_Int_Bool_unlockFork2,Go) [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K,MyDTBool_Bool)] > (call_main_map'_Int_Bool_goMux2,MyDTBool_Bool) */
  assign \call_main_map'_Int_Bool_goMux2_d  = (\call_main_map'_Int_Bool_unlockFork2_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d [0]);
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_r  = (\call_main_map'_Int_Bool_goMux2_r  && (\call_main_map'_Int_Bool_unlockFork2_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d [0]));
  assign \call_main_map'_Int_Bool_unlockFork2_r  = (\call_main_map'_Int_Bool_goMux2_r  && (\call_main_map'_Int_Bool_unlockFork2_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_BoolisZa8K_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_main_map'_Int_Bool_unlockFork3,Go) [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L,MyDTInt_Bool)] > (call_main_map'_Int_Bool_goMux3,MyDTInt_Bool) */
  assign \call_main_map'_Int_Bool_goMux3_d  = (\call_main_map'_Int_Bool_unlockFork3_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d [0]);
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_r  = (\call_main_map'_Int_Bool_goMux3_r  && (\call_main_map'_Int_Bool_unlockFork3_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d [0]));
  assign \call_main_map'_Int_Bool_unlockFork3_r  = (\call_main_map'_Int_Bool_goMux3_r  && (\call_main_map'_Int_Bool_unlockFork3_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolga8L_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_main_map'_Int_Bool_unlockFork4,Go) [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M,Pointer_QTree_Int)] > (call_main_map'_Int_Bool_goMux4,Pointer_QTree_Int) */
  assign \call_main_map'_Int_Bool_goMux4_d  = {\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d [16:1],
                                               (\call_main_map'_Int_Bool_unlockFork4_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d [0])};
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_r  = (\call_main_map'_Int_Bool_goMux4_r  && (\call_main_map'_Int_Bool_unlockFork4_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d [0]));
  assign \call_main_map'_Int_Bool_unlockFork4_r  = (\call_main_map'_Int_Bool_goMux4_r  && (\call_main_map'_Int_Bool_unlockFork4_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolma8M_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_map'_Int_Bool) : (call_main_map'_Int_Bool_unlockFork5,Go) [(call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2,Pointer_CTmain_map'_Int_Bool)] > (call_main_map'_Int_Bool_goMux5,Pointer_CTmain_map'_Int_Bool) */
  assign \call_main_map'_Int_Bool_goMux5_d  = {\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d [16:1],
                                               (\call_main_map'_Int_Bool_unlockFork5_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d [0])};
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_r  = (\call_main_map'_Int_Bool_goMux5_r  && (\call_main_map'_Int_Bool_unlockFork5_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d [0]));
  assign \call_main_map'_Int_Bool_unlockFork5_r  = (\call_main_map'_Int_Bool_goMux5_r  && (\call_main_map'_Int_Bool_unlockFork5_d [0] && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Boolsc_0_2_d [0]));
  
  /* sink (Ty Int) : (es_0_1I#,Int) > */
  assign {\es_0_1I#_r , \es_0_1I#_dout } = {\es_0_1I#_rout ,
                                            \es_0_1I#_d };
  
  /* buf (Ty Int) : (es_0_2_1I#_mux_mux_mux,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t \es_0_2_1I#_mux_mux_mux_bufchan_d ;
  logic \es_0_2_1I#_mux_mux_mux_bufchan_r ;
  assign \es_0_2_1I#_mux_mux_mux_r  = ((! \es_0_2_1I#_mux_mux_mux_bufchan_d [0]) || \es_0_2_1I#_mux_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_2_1I#_mux_mux_mux_bufchan_d  <= {32'd0, 1'd0};
    else
      if (\es_0_2_1I#_mux_mux_mux_r )
        \es_0_2_1I#_mux_mux_mux_bufchan_d  <= \es_0_2_1I#_mux_mux_mux_d ;
  Int_t \es_0_2_1I#_mux_mux_mux_bufchan_buf ;
  assign \es_0_2_1I#_mux_mux_mux_bufchan_r  = (! \es_0_2_1I#_mux_mux_mux_bufchan_buf [0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (\es_0_2_1I#_mux_mux_mux_bufchan_buf [0] ? \es_0_2_1I#_mux_mux_mux_bufchan_buf  :
                                          \es_0_2_1I#_mux_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \es_0_2_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && \es_0_2_1I#_mux_mux_mux_bufchan_buf [0]))
        \es_0_2_1I#_mux_mux_mux_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! \es_0_2_1I#_mux_mux_mux_bufchan_buf [0])))
        \es_0_2_1I#_mux_mux_mux_bufchan_buf  <= \es_0_2_1I#_mux_mux_mux_bufchan_d ;
  
  /* buf (Ty QTree_Int) : (es_0_3_1QVal_Int,QTree_Int) > (lizzieLet7_1_1_argbuf,QTree_Int) */
  QTree_Int_t es_0_3_1QVal_Int_bufchan_d;
  logic es_0_3_1QVal_Int_bufchan_r;
  assign es_0_3_1QVal_Int_r = ((! es_0_3_1QVal_Int_bufchan_d[0]) || es_0_3_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_3_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_3_1QVal_Int_r)
        es_0_3_1QVal_Int_bufchan_d <= es_0_3_1QVal_Int_d;
  QTree_Int_t es_0_3_1QVal_Int_bufchan_buf;
  assign es_0_3_1QVal_Int_bufchan_r = (! es_0_3_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (es_0_3_1QVal_Int_bufchan_buf[0] ? es_0_3_1QVal_Int_bufchan_buf :
                                    es_0_3_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && es_0_3_1QVal_Int_bufchan_buf[0]))
        es_0_3_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! es_0_3_1QVal_Int_bufchan_buf[0])))
        es_0_3_1QVal_Int_bufchan_buf <= es_0_3_1QVal_Int_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_4_1,MyBool) (lizzieLet17_4QVal_Int_3,Go) > [(es_0_4_1MyFalse,Go),
                                                                  (es_0_4_1MyTrue,Go)] */
  logic [1:0] lizzieLet17_4QVal_Int_3_onehotd;
  always_comb
    if ((es_0_4_1_d[0] && lizzieLet17_4QVal_Int_3_d[0]))
      unique case (es_0_4_1_d[1:1])
        1'd0: lizzieLet17_4QVal_Int_3_onehotd = 2'd1;
        1'd1: lizzieLet17_4QVal_Int_3_onehotd = 2'd2;
        default: lizzieLet17_4QVal_Int_3_onehotd = 2'd0;
      endcase
    else lizzieLet17_4QVal_Int_3_onehotd = 2'd0;
  assign es_0_4_1MyFalse_d = lizzieLet17_4QVal_Int_3_onehotd[0];
  assign es_0_4_1MyTrue_d = lizzieLet17_4QVal_Int_3_onehotd[1];
  assign lizzieLet17_4QVal_Int_3_r = (| (lizzieLet17_4QVal_Int_3_onehotd & {es_0_4_1MyTrue_r,
                                                                            es_0_4_1MyFalse_r}));
  assign es_0_4_1_r = lizzieLet17_4QVal_Int_3_r;
  
  /* buf (Ty Go) : (es_0_4_1MyFalse,Go) > (es_0_4_1MyFalse_1_argbuf,Go) */
  Go_t es_0_4_1MyFalse_bufchan_d;
  logic es_0_4_1MyFalse_bufchan_r;
  assign es_0_4_1MyFalse_r = ((! es_0_4_1MyFalse_bufchan_d[0]) || es_0_4_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_4_1MyFalse_r)
        es_0_4_1MyFalse_bufchan_d <= es_0_4_1MyFalse_d;
  Go_t es_0_4_1MyFalse_bufchan_buf;
  assign es_0_4_1MyFalse_bufchan_r = (! es_0_4_1MyFalse_bufchan_buf[0]);
  assign es_0_4_1MyFalse_1_argbuf_d = (es_0_4_1MyFalse_bufchan_buf[0] ? es_0_4_1MyFalse_bufchan_buf :
                                       es_0_4_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_4_1MyFalse_1_argbuf_r && es_0_4_1MyFalse_bufchan_buf[0]))
        es_0_4_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_4_1MyFalse_1_argbuf_r) && (! es_0_4_1MyFalse_bufchan_buf[0])))
        es_0_4_1MyFalse_bufchan_buf <= es_0_4_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_4_1MyTrue,Go) > [(es_0_4_1MyTrue_1,Go),
                                      (es_0_4_1MyTrue_2,Go)] */
  logic [1:0] es_0_4_1MyTrue_emitted;
  logic [1:0] es_0_4_1MyTrue_done;
  assign es_0_4_1MyTrue_1_d = (es_0_4_1MyTrue_d[0] && (! es_0_4_1MyTrue_emitted[0]));
  assign es_0_4_1MyTrue_2_d = (es_0_4_1MyTrue_d[0] && (! es_0_4_1MyTrue_emitted[1]));
  assign es_0_4_1MyTrue_done = (es_0_4_1MyTrue_emitted | ({es_0_4_1MyTrue_2_d[0],
                                                           es_0_4_1MyTrue_1_d[0]} & {es_0_4_1MyTrue_2_r,
                                                                                     es_0_4_1MyTrue_1_r}));
  assign es_0_4_1MyTrue_r = (& es_0_4_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_emitted <= 2'd0;
    else
      es_0_4_1MyTrue_emitted <= (es_0_4_1MyTrue_r ? 2'd0 :
                                 es_0_4_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(es_0_4_1MyTrue_1,Go)] > (es_0_4_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign es_0_4_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {es_0_4_1MyTrue_1_d[0]}), es_0_4_1MyTrue_1_d);
  assign {es_0_4_1MyTrue_1_r} = {1 {(es_0_4_1MyTrue_1QNone_Bool_r && es_0_4_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_4_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet20_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_4_1MyTrue_1QNone_Bool_bufchan_d;
  logic es_0_4_1MyTrue_1QNone_Bool_bufchan_r;
  assign es_0_4_1MyTrue_1QNone_Bool_r = ((! es_0_4_1MyTrue_1QNone_Bool_bufchan_d[0]) || es_0_4_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_4_1MyTrue_1QNone_Bool_r)
        es_0_4_1MyTrue_1QNone_Bool_bufchan_d <= es_0_4_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t es_0_4_1MyTrue_1QNone_Bool_bufchan_buf;
  assign es_0_4_1MyTrue_1QNone_Bool_bufchan_r = (! es_0_4_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (es_0_4_1MyTrue_1QNone_Bool_bufchan_buf[0] ? es_0_4_1MyTrue_1QNone_Bool_bufchan_buf :
                                   es_0_4_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && es_0_4_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        es_0_4_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! es_0_4_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        es_0_4_1MyTrue_1QNone_Bool_bufchan_buf <= es_0_4_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (es_0_4_1MyTrue_2,Go) > (es_0_4_1MyTrue_2_argbuf,Go) */
  Go_t es_0_4_1MyTrue_2_bufchan_d;
  logic es_0_4_1MyTrue_2_bufchan_r;
  assign es_0_4_1MyTrue_2_r = ((! es_0_4_1MyTrue_2_bufchan_d[0]) || es_0_4_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_4_1MyTrue_2_r)
        es_0_4_1MyTrue_2_bufchan_d <= es_0_4_1MyTrue_2_d;
  Go_t es_0_4_1MyTrue_2_bufchan_buf;
  assign es_0_4_1MyTrue_2_bufchan_r = (! es_0_4_1MyTrue_2_bufchan_buf[0]);
  assign es_0_4_1MyTrue_2_argbuf_d = (es_0_4_1MyTrue_2_bufchan_buf[0] ? es_0_4_1MyTrue_2_bufchan_buf :
                                      es_0_4_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_4_1MyTrue_2_argbuf_r && es_0_4_1MyTrue_2_bufchan_buf[0]))
        es_0_4_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_4_1MyTrue_2_argbuf_r) && (! es_0_4_1MyTrue_2_bufchan_buf[0])))
        es_0_4_1MyTrue_2_bufchan_buf <= es_0_4_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmain_map'_Int_Bool) : (es_0_4_2,MyBool) (lizzieLet17_6QVal_Int,Pointer_CTmain_map'_Int_Bool) > [(es_0_4_2MyFalse,Pointer_CTmain_map'_Int_Bool),
                                                                                                                    (es_0_4_2MyTrue,Pointer_CTmain_map'_Int_Bool)] */
  logic [1:0] lizzieLet17_6QVal_Int_onehotd;
  always_comb
    if ((es_0_4_2_d[0] && lizzieLet17_6QVal_Int_d[0]))
      unique case (es_0_4_2_d[1:1])
        1'd0: lizzieLet17_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet17_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet17_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet17_6QVal_Int_onehotd = 2'd0;
  assign es_0_4_2MyFalse_d = {lizzieLet17_6QVal_Int_d[16:1],
                              lizzieLet17_6QVal_Int_onehotd[0]};
  assign es_0_4_2MyTrue_d = {lizzieLet17_6QVal_Int_d[16:1],
                             lizzieLet17_6QVal_Int_onehotd[1]};
  assign lizzieLet17_6QVal_Int_r = (| (lizzieLet17_6QVal_Int_onehotd & {es_0_4_2MyTrue_r,
                                                                        es_0_4_2MyFalse_r}));
  assign es_0_4_2_r = lizzieLet17_6QVal_Int_r;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (es_0_4_2MyFalse,Pointer_CTmain_map'_Int_Bool) > (es_0_4_2MyFalse_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyFalse_bufchan_d;
  logic es_0_4_2MyFalse_bufchan_r;
  assign es_0_4_2MyFalse_r = ((! es_0_4_2MyFalse_bufchan_d[0]) || es_0_4_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_4_2MyFalse_r)
        es_0_4_2MyFalse_bufchan_d <= es_0_4_2MyFalse_d;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyFalse_bufchan_buf;
  assign es_0_4_2MyFalse_bufchan_r = (! es_0_4_2MyFalse_bufchan_buf[0]);
  assign es_0_4_2MyFalse_1_argbuf_d = (es_0_4_2MyFalse_bufchan_buf[0] ? es_0_4_2MyFalse_bufchan_buf :
                                       es_0_4_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_4_2MyFalse_1_argbuf_r && es_0_4_2MyFalse_bufchan_buf[0]))
        es_0_4_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_4_2MyFalse_1_argbuf_r) && (! es_0_4_2MyFalse_bufchan_buf[0])))
        es_0_4_2MyFalse_bufchan_buf <= es_0_4_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (es_0_4_2MyTrue,Pointer_CTmain_map'_Int_Bool) > (es_0_4_2MyTrue_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyTrue_bufchan_d;
  logic es_0_4_2MyTrue_bufchan_r;
  assign es_0_4_2MyTrue_r = ((! es_0_4_2MyTrue_bufchan_d[0]) || es_0_4_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_4_2MyTrue_r) es_0_4_2MyTrue_bufchan_d <= es_0_4_2MyTrue_d;
  \Pointer_CTmain_map'_Int_Bool_t  es_0_4_2MyTrue_bufchan_buf;
  assign es_0_4_2MyTrue_bufchan_r = (! es_0_4_2MyTrue_bufchan_buf[0]);
  assign es_0_4_2MyTrue_1_argbuf_d = (es_0_4_2MyTrue_bufchan_buf[0] ? es_0_4_2MyTrue_bufchan_buf :
                                      es_0_4_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_4_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_4_2MyTrue_1_argbuf_r && es_0_4_2MyTrue_bufchan_buf[0]))
        es_0_4_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_4_2MyTrue_1_argbuf_r) && (! es_0_4_2MyTrue_bufchan_buf[0])))
        es_0_4_2MyTrue_bufchan_buf <= es_0_4_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (es_0_4_3,MyBool) (xa88_2,MyBool) > [(es_0_4_3MyFalse,MyBool),
                                                         (_59,MyBool)] */
  logic [1:0] xa88_2_onehotd;
  always_comb
    if ((es_0_4_3_d[0] && xa88_2_d[0]))
      unique case (es_0_4_3_d[1:1])
        1'd0: xa88_2_onehotd = 2'd1;
        1'd1: xa88_2_onehotd = 2'd2;
        default: xa88_2_onehotd = 2'd0;
      endcase
    else xa88_2_onehotd = 2'd0;
  assign es_0_4_3MyFalse_d = {xa88_2_d[1:1], xa88_2_onehotd[0]};
  assign _59_d = {xa88_2_d[1:1], xa88_2_onehotd[1]};
  assign xa88_2_r = (| (xa88_2_onehotd & {_59_r,
                                          es_0_4_3MyFalse_r}));
  assign es_0_4_3_r = xa88_2_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(es_0_4_3MyFalse,MyBool)] > (es_0_4_3MyFalse_1QVal_Bool,QTree_Bool) */
  assign es_0_4_3MyFalse_1QVal_Bool_d = QVal_Bool_dc((& {es_0_4_3MyFalse_d[0]}), es_0_4_3MyFalse_d);
  assign {es_0_4_3MyFalse_r} = {1 {(es_0_4_3MyFalse_1QVal_Bool_r && es_0_4_3MyFalse_1QVal_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_4_3MyFalse_1QVal_Bool,QTree_Bool) > (lizzieLet19_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_4_3MyFalse_1QVal_Bool_bufchan_d;
  logic es_0_4_3MyFalse_1QVal_Bool_bufchan_r;
  assign es_0_4_3MyFalse_1QVal_Bool_r = ((! es_0_4_3MyFalse_1QVal_Bool_bufchan_d[0]) || es_0_4_3MyFalse_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_3MyFalse_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_4_3MyFalse_1QVal_Bool_r)
        es_0_4_3MyFalse_1QVal_Bool_bufchan_d <= es_0_4_3MyFalse_1QVal_Bool_d;
  QTree_Bool_t es_0_4_3MyFalse_1QVal_Bool_bufchan_buf;
  assign es_0_4_3MyFalse_1QVal_Bool_bufchan_r = (! es_0_4_3MyFalse_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet19_1_argbuf_d = (es_0_4_3MyFalse_1QVal_Bool_bufchan_buf[0] ? es_0_4_3MyFalse_1QVal_Bool_bufchan_buf :
                                   es_0_4_3MyFalse_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_4_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet19_1_argbuf_r && es_0_4_3MyFalse_1QVal_Bool_bufchan_buf[0]))
        es_0_4_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet19_1_argbuf_r) && (! es_0_4_3MyFalse_1QVal_Bool_bufchan_buf[0])))
        es_0_4_3MyFalse_1QVal_Bool_bufchan_buf <= es_0_4_3MyFalse_1QVal_Bool_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32,Int#) > (contRet_0_1_1_argbuf,Int#) */
  \Int#_t  es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d;
  logic es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_r;
  assign es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_r = ((! es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d[0]) || es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d <= {32'd0,
                                                              1'd0};
    else
      if (es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_r)
        es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d <= es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_d;
  \Int#_t  es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf;
  assign es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_r = (! es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf[0] ? es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf :
                                   es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf[0]))
        es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf <= {32'd0,
                                                                  1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf[0])))
        es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_buf <= es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_1ww2XmM_1_1_Add32,Int#) (lizzieLet29_4Lcall_$wnnz0,Int#) > (es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32,Int#) */
  assign es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_d = {(es_6_1ww2XmM_1_1_Add32_d[32:1] + lizzieLet29_4Lcall_$wnnz0_d[32:1]),
                                                        (es_6_1ww2XmM_1_1_Add32_d[0] && lizzieLet29_4Lcall_$wnnz0_d[0])};
  assign {es_6_1ww2XmM_1_1_Add32_r,
          lizzieLet29_4Lcall_$wnnz0_r} = {2 {(es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_r && es_4_4_1lizzieLet29_4Lcall_$wnnz0_1_Add32_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (ga8L_2_2,MyDTInt_Bool) > (ga8L_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t ga8L_2_2_bufchan_d;
  logic ga8L_2_2_bufchan_r;
  assign ga8L_2_2_r = ((! ga8L_2_2_bufchan_d[0]) || ga8L_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_2_2_bufchan_d <= 1'd0;
    else if (ga8L_2_2_r) ga8L_2_2_bufchan_d <= ga8L_2_2_d;
  MyDTInt_Bool_t ga8L_2_2_bufchan_buf;
  assign ga8L_2_2_bufchan_r = (! ga8L_2_2_bufchan_buf[0]);
  assign ga8L_2_2_argbuf_d = (ga8L_2_2_bufchan_buf[0] ? ga8L_2_2_bufchan_buf :
                              ga8L_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_2_2_bufchan_buf <= 1'd0;
    else
      if ((ga8L_2_2_argbuf_r && ga8L_2_2_bufchan_buf[0]))
        ga8L_2_2_bufchan_buf <= 1'd0;
      else if (((! ga8L_2_2_argbuf_r) && (! ga8L_2_2_bufchan_buf[0])))
        ga8L_2_2_bufchan_buf <= ga8L_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (ga8L_2_destruct,MyDTInt_Bool) > [(ga8L_2_1,MyDTInt_Bool),
                                                           (ga8L_2_2,MyDTInt_Bool)] */
  logic [1:0] ga8L_2_destruct_emitted;
  logic [1:0] ga8L_2_destruct_done;
  assign ga8L_2_1_d = (ga8L_2_destruct_d[0] && (! ga8L_2_destruct_emitted[0]));
  assign ga8L_2_2_d = (ga8L_2_destruct_d[0] && (! ga8L_2_destruct_emitted[1]));
  assign ga8L_2_destruct_done = (ga8L_2_destruct_emitted | ({ga8L_2_2_d[0],
                                                             ga8L_2_1_d[0]} & {ga8L_2_2_r,
                                                                               ga8L_2_1_r}));
  assign ga8L_2_destruct_r = (& ga8L_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_2_destruct_emitted <= 2'd0;
    else
      ga8L_2_destruct_emitted <= (ga8L_2_destruct_r ? 2'd0 :
                                  ga8L_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (ga8L_3_2,MyDTInt_Bool) > (ga8L_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t ga8L_3_2_bufchan_d;
  logic ga8L_3_2_bufchan_r;
  assign ga8L_3_2_r = ((! ga8L_3_2_bufchan_d[0]) || ga8L_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_3_2_bufchan_d <= 1'd0;
    else if (ga8L_3_2_r) ga8L_3_2_bufchan_d <= ga8L_3_2_d;
  MyDTInt_Bool_t ga8L_3_2_bufchan_buf;
  assign ga8L_3_2_bufchan_r = (! ga8L_3_2_bufchan_buf[0]);
  assign ga8L_3_2_argbuf_d = (ga8L_3_2_bufchan_buf[0] ? ga8L_3_2_bufchan_buf :
                              ga8L_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_3_2_bufchan_buf <= 1'd0;
    else
      if ((ga8L_3_2_argbuf_r && ga8L_3_2_bufchan_buf[0]))
        ga8L_3_2_bufchan_buf <= 1'd0;
      else if (((! ga8L_3_2_argbuf_r) && (! ga8L_3_2_bufchan_buf[0])))
        ga8L_3_2_bufchan_buf <= ga8L_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (ga8L_3_destruct,MyDTInt_Bool) > [(ga8L_3_1,MyDTInt_Bool),
                                                           (ga8L_3_2,MyDTInt_Bool)] */
  logic [1:0] ga8L_3_destruct_emitted;
  logic [1:0] ga8L_3_destruct_done;
  assign ga8L_3_1_d = (ga8L_3_destruct_d[0] && (! ga8L_3_destruct_emitted[0]));
  assign ga8L_3_2_d = (ga8L_3_destruct_d[0] && (! ga8L_3_destruct_emitted[1]));
  assign ga8L_3_destruct_done = (ga8L_3_destruct_emitted | ({ga8L_3_2_d[0],
                                                             ga8L_3_1_d[0]} & {ga8L_3_2_r,
                                                                               ga8L_3_1_r}));
  assign ga8L_3_destruct_r = (& ga8L_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_3_destruct_emitted <= 2'd0;
    else
      ga8L_3_destruct_emitted <= (ga8L_3_destruct_r ? 2'd0 :
                                  ga8L_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (ga8L_4_destruct,MyDTInt_Bool) > (ga8L_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t ga8L_4_destruct_bufchan_d;
  logic ga8L_4_destruct_bufchan_r;
  assign ga8L_4_destruct_r = ((! ga8L_4_destruct_bufchan_d[0]) || ga8L_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_4_destruct_bufchan_d <= 1'd0;
    else
      if (ga8L_4_destruct_r)
        ga8L_4_destruct_bufchan_d <= ga8L_4_destruct_d;
  MyDTInt_Bool_t ga8L_4_destruct_bufchan_buf;
  assign ga8L_4_destruct_bufchan_r = (! ga8L_4_destruct_bufchan_buf[0]);
  assign ga8L_4_1_argbuf_d = (ga8L_4_destruct_bufchan_buf[0] ? ga8L_4_destruct_bufchan_buf :
                              ga8L_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ga8L_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((ga8L_4_1_argbuf_r && ga8L_4_destruct_bufchan_buf[0]))
        ga8L_4_destruct_bufchan_buf <= 1'd0;
      else if (((! ga8L_4_1_argbuf_r) && (! ga8L_4_destruct_bufchan_buf[0])))
        ga8L_4_destruct_bufchan_buf <= ga8L_4_destruct_bufchan_d;
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5),
                                          (go_11_goMux_choice_3,C5),
                                          (go_11_goMux_choice_4,C5)] */
  logic [3:0] go_11_goMux_choice_emitted;
  logic [3:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_3_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[2]))};
  assign go_11_goMux_choice_4_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[3]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_4_d[0],
                                                                   go_11_goMux_choice_3_d[0],
                                                                   go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_4_r,
                                                                                                 go_11_goMux_choice_3_r,
                                                                                                 go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 4'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 4'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_11_goMux_choice_1,C5) [(call_$wmAdd_Int_goMux2,MyDTInt_Int_Int),
                                                      (wslR_2_2_argbuf,MyDTInt_Int_Int),
                                                      (wslR_3_2_argbuf,MyDTInt_Int_Int),
                                                      (wslR_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (wslR_1_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] wslR_1_goMux_mux_mux;
  logic [4:0] wslR_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd1,
                                                           call_$wmAdd_Int_goMux2_d};
      3'd1:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd2,
                                                           wslR_2_2_argbuf_d};
      3'd2:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd4,
                                                           wslR_3_2_argbuf_d};
      3'd3:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd8,
                                                           wslR_4_1_argbuf_d};
      3'd4:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd16,
                                                           lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_d};
      default:
        {wslR_1_goMux_mux_onehot, wslR_1_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign wslR_1_goMux_mux_d = (wslR_1_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0]);
  assign go_11_goMux_choice_1_r = (wslR_1_goMux_mux_d[0] && wslR_1_goMux_mux_r);
  assign {lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_r,
          wslR_4_1_argbuf_r,
          wslR_3_2_argbuf_r,
          wslR_2_2_argbuf_r,
          call_$wmAdd_Int_goMux2_r} = (go_11_goMux_choice_1_r ? wslR_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_2,C5) [(call_$wmAdd_Int_goMux3,Pointer_QTree_Int),
                                                        (q3a8l_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2a8k_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1a8j_3_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int)] > (w1slS_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] w1slS_1_goMux_mux_mux;
  logic [4:0] w1slS_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Int_goMux3_d};
      3'd1:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd2,
                                                             q3a8l_1_1_argbuf_d};
      3'd2:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd4,
                                                             q2a8k_2_1_argbuf_d};
      3'd3:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd8,
                                                             q1a8j_3_1_argbuf_d};
      3'd4:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd16,
                                                             lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_d};
      default:
        {w1slS_1_goMux_mux_onehot, w1slS_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w1slS_1_goMux_mux_d = {w1slS_1_goMux_mux_mux[16:1],
                                (w1slS_1_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0])};
  assign go_11_goMux_choice_2_r = (w1slS_1_goMux_mux_d[0] && w1slS_1_goMux_mux_r);
  assign {lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_r,
          q1a8j_3_1_argbuf_r,
          q2a8k_2_1_argbuf_r,
          q3a8l_1_1_argbuf_r,
          call_$wmAdd_Int_goMux3_r} = (go_11_goMux_choice_2_r ? w1slS_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_3,C5) [(call_$wmAdd_Int_goMux4,Pointer_QTree_Int),
                                                        (t3a8q_1_1_argbuf,Pointer_QTree_Int),
                                                        (t2a8p_2_1_argbuf,Pointer_QTree_Int),
                                                        (t1a8o_3_1_argbuf,Pointer_QTree_Int),
                                                        (t4a8r_1_argbuf,Pointer_QTree_Int)] > (w2slT_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] w2slT_1_goMux_mux_mux;
  logic [4:0] w2slT_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_3_d[3:1])
      3'd0:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Int_goMux4_d};
      3'd1:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd2,
                                                             t3a8q_1_1_argbuf_d};
      3'd2:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd4,
                                                             t2a8p_2_1_argbuf_d};
      3'd3:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd8,
                                                             t1a8o_3_1_argbuf_d};
      3'd4:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd16,
                                                             t4a8r_1_argbuf_d};
      default:
        {w2slT_1_goMux_mux_onehot, w2slT_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w2slT_1_goMux_mux_d = {w2slT_1_goMux_mux_mux[16:1],
                                (w2slT_1_goMux_mux_mux[0] && go_11_goMux_choice_3_d[0])};
  assign go_11_goMux_choice_3_r = (w2slT_1_goMux_mux_d[0] && w2slT_1_goMux_mux_r);
  assign {t4a8r_1_argbuf_r,
          t1a8o_3_1_argbuf_r,
          t2a8p_2_1_argbuf_r,
          t3a8q_1_1_argbuf_r,
          call_$wmAdd_Int_goMux4_r} = (go_11_goMux_choice_3_r ? w2slT_1_goMux_mux_onehot :
                                       5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wmAdd_Int) : (go_11_goMux_choice_4,C5) [(call_$wmAdd_Int_goMux5,Pointer_CT$wmAdd_Int),
                                                           (sca2_1_argbuf,Pointer_CT$wmAdd_Int),
                                                           (sca1_1_argbuf,Pointer_CT$wmAdd_Int),
                                                           (sca0_1_argbuf,Pointer_CT$wmAdd_Int),
                                                           (sca3_1_argbuf,Pointer_CT$wmAdd_Int)] > (sc_0_goMux_mux,Pointer_CT$wmAdd_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wmAdd_Int_goMux5_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_11_goMux_choice_4_d[0])};
  assign go_11_goMux_choice_4_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wmAdd_Int_goMux5_r} = (go_11_goMux_choice_4_r ? sc_0_goMux_mux_onehot :
                                       5'd0);
  
  /* fork (Ty C5) : (go_12_goMux_choice,C5) > [(go_12_goMux_choice_1,C5),
                                          (go_12_goMux_choice_2,C5)] */
  logic [1:0] go_12_goMux_choice_emitted;
  logic [1:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 2'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 2'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_12_goMux_choice_1,C5) [(call_$wnnz_goMux2,Pointer_QTree_Bool),
                                                         (q2a93_1_1_argbuf,Pointer_QTree_Bool),
                                                         (q3a94_2_1_argbuf,Pointer_QTree_Bool),
                                                         (q4a95_3_1_argbuf,Pointer_QTree_Bool),
                                                         (q1a92_1_argbuf,Pointer_QTree_Bool)] > (wslW_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] wslW_1_goMux_mux_mux;
  logic [4:0] wslW_1_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_goMux2_d};
      3'd1:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd2,
                                                           q2a93_1_1_argbuf_d};
      3'd2:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd4,
                                                           q3a94_2_1_argbuf_d};
      3'd3:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd8,
                                                           q4a95_3_1_argbuf_d};
      3'd4:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd16,
                                                           q1a92_1_argbuf_d};
      default:
        {wslW_1_goMux_mux_onehot, wslW_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wslW_1_goMux_mux_d = {wslW_1_goMux_mux_mux[16:1],
                               (wslW_1_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0])};
  assign go_12_goMux_choice_1_r = (wslW_1_goMux_mux_d[0] && wslW_1_goMux_mux_r);
  assign {q1a92_1_argbuf_r,
          q4a95_3_1_argbuf_r,
          q3a94_2_1_argbuf_r,
          q2a93_1_1_argbuf_r,
          call_$wnnz_goMux2_r} = (go_12_goMux_choice_1_r ? wslW_1_goMux_mux_onehot :
                                  5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz) : (go_12_goMux_choice_2,C5) [(call_$wnnz_goMux3,Pointer_CT$wnnz),
                                                      (sca2_1_1_argbuf,Pointer_CT$wnnz),
                                                      (sca1_1_1_argbuf,Pointer_CT$wnnz),
                                                      (sca0_1_1_argbuf,Pointer_CT$wnnz),
                                                      (sca3_1_1_argbuf,Pointer_CT$wnnz)] > (sc_0_1_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_goMux3_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0])};
  assign go_12_goMux_choice_2_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_$wnnz_goMux3_r} = (go_12_goMux_choice_2_r ? sc_0_1_goMux_mux_onehot :
                                  5'd0);
  
  /* fork (Ty C5) : (go_13_goMux_choice,C5) > [(go_13_goMux_choice_1,C5),
                                          (go_13_goMux_choice_2,C5),
                                          (go_13_goMux_choice_3,C5),
                                          (go_13_goMux_choice_4,C5)] */
  logic [3:0] go_13_goMux_choice_emitted;
  logic [3:0] go_13_goMux_choice_done;
  assign go_13_goMux_choice_1_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[0]))};
  assign go_13_goMux_choice_2_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[1]))};
  assign go_13_goMux_choice_3_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[2]))};
  assign go_13_goMux_choice_4_d = {go_13_goMux_choice_d[3:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[3]))};
  assign go_13_goMux_choice_done = (go_13_goMux_choice_emitted | ({go_13_goMux_choice_4_d[0],
                                                                   go_13_goMux_choice_3_d[0],
                                                                   go_13_goMux_choice_2_d[0],
                                                                   go_13_goMux_choice_1_d[0]} & {go_13_goMux_choice_4_r,
                                                                                                 go_13_goMux_choice_3_r,
                                                                                                 go_13_goMux_choice_2_r,
                                                                                                 go_13_goMux_choice_1_r}));
  assign go_13_goMux_choice_r = (& go_13_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_goMux_choice_emitted <= 4'd0;
    else
      go_13_goMux_choice_emitted <= (go_13_goMux_choice_r ? 4'd0 :
                                     go_13_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool) : (go_13_goMux_choice_1,C5) [(call_main_map'_Int_Bool_goMux2,MyDTBool_Bool),
                                                    (isZa8K_2_2_argbuf,MyDTBool_Bool),
                                                    (isZa8K_3_2_argbuf,MyDTBool_Bool),
                                                    (isZa8K_4_1_argbuf,MyDTBool_Bool),
                                                    (lizzieLet17_5QNode_Int_2_argbuf,MyDTBool_Bool)] > (isZa8K_goMux_mux,MyDTBool_Bool) */
  logic [0:0] isZa8K_goMux_mux_mux;
  logic [4:0] isZa8K_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_1_d[3:1])
      3'd0:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Int_Bool_goMux2_d };
      3'd1:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd2,
                                                           isZa8K_2_2_argbuf_d};
      3'd2:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd4,
                                                           isZa8K_3_2_argbuf_d};
      3'd3:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd8,
                                                           isZa8K_4_1_argbuf_d};
      3'd4:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd16,
                                                           lizzieLet17_5QNode_Int_2_argbuf_d};
      default:
        {isZa8K_goMux_mux_onehot, isZa8K_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZa8K_goMux_mux_d = (isZa8K_goMux_mux_mux[0] && go_13_goMux_choice_1_d[0]);
  assign go_13_goMux_choice_1_r = (isZa8K_goMux_mux_d[0] && isZa8K_goMux_mux_r);
  assign {lizzieLet17_5QNode_Int_2_argbuf_r,
          isZa8K_4_1_argbuf_r,
          isZa8K_3_2_argbuf_r,
          isZa8K_2_2_argbuf_r,
          \call_main_map'_Int_Bool_goMux2_r } = (go_13_goMux_choice_1_r ? isZa8K_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_13_goMux_choice_2,C5) [(call_main_map'_Int_Bool_goMux3,MyDTInt_Bool),
                                                   (ga8L_2_2_argbuf,MyDTInt_Bool),
                                                   (ga8L_3_2_argbuf,MyDTInt_Bool),
                                                   (ga8L_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet17_3QNode_Int_2_argbuf,MyDTInt_Bool)] > (ga8L_goMux_mux,MyDTInt_Bool) */
  logic [0:0] ga8L_goMux_mux_mux;
  logic [4:0] ga8L_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_2_d[3:1])
      3'd0:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Int_Bool_goMux3_d };
      3'd1:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd2,
                                                       ga8L_2_2_argbuf_d};
      3'd2:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd4,
                                                       ga8L_3_2_argbuf_d};
      3'd3:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd8,
                                                       ga8L_4_1_argbuf_d};
      3'd4:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd16,
                                                       lizzieLet17_3QNode_Int_2_argbuf_d};
      default:
        {ga8L_goMux_mux_onehot, ga8L_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign ga8L_goMux_mux_d = (ga8L_goMux_mux_mux[0] && go_13_goMux_choice_2_d[0]);
  assign go_13_goMux_choice_2_r = (ga8L_goMux_mux_d[0] && ga8L_goMux_mux_r);
  assign {lizzieLet17_3QNode_Int_2_argbuf_r,
          ga8L_4_1_argbuf_r,
          ga8L_3_2_argbuf_r,
          ga8L_2_2_argbuf_r,
          \call_main_map'_Int_Bool_goMux3_r } = (go_13_goMux_choice_2_r ? ga8L_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_13_goMux_choice_3,C5) [(call_main_map'_Int_Bool_goMux4,Pointer_QTree_Int),
                                                        (q3a8Q_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2a8P_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1a8O_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4a8R_1_argbuf,Pointer_QTree_Int)] > (ma8M_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] ma8M_goMux_mux_mux;
  logic [4:0] ma8M_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_3_d[3:1])
      3'd0:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Int_Bool_goMux4_d };
      3'd1:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd2,
                                                       q3a8Q_1_1_argbuf_d};
      3'd2:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd4,
                                                       q2a8P_2_1_argbuf_d};
      3'd3:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd8,
                                                       q1a8O_3_1_argbuf_d};
      3'd4:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd16,
                                                       q4a8R_1_argbuf_d};
      default:
        {ma8M_goMux_mux_onehot, ma8M_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign ma8M_goMux_mux_d = {ma8M_goMux_mux_mux[16:1],
                             (ma8M_goMux_mux_mux[0] && go_13_goMux_choice_3_d[0])};
  assign go_13_goMux_choice_3_r = (ma8M_goMux_mux_d[0] && ma8M_goMux_mux_r);
  assign {q4a8R_1_argbuf_r,
          q1a8O_3_1_argbuf_r,
          q2a8P_2_1_argbuf_r,
          q3a8Q_1_1_argbuf_r,
          \call_main_map'_Int_Bool_goMux4_r } = (go_13_goMux_choice_3_r ? ma8M_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Int_Bool) : (go_13_goMux_choice_4,C5) [(call_main_map'_Int_Bool_goMux5,Pointer_CTmain_map'_Int_Bool),
                                                                   (sca2_2_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (sca1_2_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (sca0_2_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (sca3_2_1_argbuf,Pointer_CTmain_map'_Int_Bool)] > (sc_0_2_goMux_mux,Pointer_CTmain_map'_Int_Bool) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Int_Bool_goMux5_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_13_goMux_choice_4_d[0])};
  assign go_13_goMux_choice_4_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_main_map'_Int_Bool_goMux5_r } = (go_13_goMux_choice_4_r ? sc_0_2_goMux_mux_onehot :
                                                 5'd0);
  
  /* dcon (Ty CTmain_map'_Int_Bool,
      Dcon Lmain_map'_Int_Boolsbos) : [(go_14_1,Go)] > (go_14_1Lmain_map'_Int_Boolsbos,CTmain_map'_Int_Bool) */
  assign \go_14_1Lmain_map'_Int_Boolsbos_d  = \Lmain_map'_Int_Boolsbos_dc ((& {go_14_1_d[0]}), go_14_1_d);
  assign {go_14_1_r} = {1 {(\go_14_1Lmain_map'_Int_Boolsbos_r  && \go_14_1Lmain_map'_Int_Boolsbos_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Bool) : (go_14_1Lmain_map'_Int_Boolsbos,CTmain_map'_Int_Bool) > (lizzieLet23_1_argbuf,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d ;
  logic \go_14_1Lmain_map'_Int_Boolsbos_bufchan_r ;
  assign \go_14_1Lmain_map'_Int_Boolsbos_r  = ((! \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d [0]) || \go_14_1Lmain_map'_Int_Boolsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d  <= {67'd0, 1'd0};
    else
      if (\go_14_1Lmain_map'_Int_Boolsbos_r )
        \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d  <= \go_14_1Lmain_map'_Int_Boolsbos_d ;
  \CTmain_map'_Int_Bool_t  \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf ;
  assign \go_14_1Lmain_map'_Int_Boolsbos_bufchan_r  = (! \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf [0]);
  assign lizzieLet23_1_argbuf_d = (\go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf [0] ? \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf  :
                                   \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf  <= {67'd0, 1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf [0]))
        \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf  <= {67'd0, 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf [0])))
        \go_14_1Lmain_map'_Int_Boolsbos_bufchan_buf  <= \go_14_1Lmain_map'_Int_Boolsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_14_2,Go) > (go_14_2_argbuf,Go) */
  Go_t go_14_2_bufchan_d;
  logic go_14_2_bufchan_r;
  assign go_14_2_r = ((! go_14_2_bufchan_d[0]) || go_14_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_d <= 1'd0;
    else if (go_14_2_r) go_14_2_bufchan_d <= go_14_2_d;
  Go_t go_14_2_bufchan_buf;
  assign go_14_2_bufchan_r = (! go_14_2_bufchan_buf[0]);
  assign go_14_2_argbuf_d = (go_14_2_bufchan_buf[0] ? go_14_2_bufchan_buf :
                             go_14_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_buf <= 1'd0;
    else
      if ((go_14_2_argbuf_r && go_14_2_bufchan_buf[0]))
        go_14_2_bufchan_buf <= 1'd0;
      else if (((! go_14_2_argbuf_r) && (! go_14_2_bufchan_buf[0])))
        go_14_2_bufchan_buf <= go_14_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool) : [(go_14_2_argbuf,Go),
                                                                                                       (isZa8K_1_1_argbuf,MyDTBool_Bool),
                                                                                                       (ga8L_1_1_argbuf,MyDTInt_Bool),
                                                                                                       (ma8M_1_1_argbuf,Pointer_QTree_Int),
                                                                                                       (lizzieLet4_1_1_argbuf,Pointer_CTmain_map'_Int_Bool)] > (call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1,TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool) */
  assign \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d  = \TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_dc ((& {go_14_2_argbuf_d[0],
                                                                                                                                                                                                                                 isZa8K_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 ga8L_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 ma8M_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 lizzieLet4_1_1_argbuf_d[0]}), go_14_2_argbuf_d, isZa8K_1_1_argbuf_d, ga8L_1_1_argbuf_d, ma8M_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_14_2_argbuf_r,
          isZa8K_1_1_argbuf_r,
          ga8L_1_1_argbuf_r,
          ma8M_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {5 {(\call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_r  && \call_main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int___Pointer_CTmain_map'_Int_Bool_1_d [0])}};
  
  /* fork (Ty C10) : (go_15_goMux_choice,C10) > [(go_15_goMux_choice_1,C10),
                                            (go_15_goMux_choice_2,C10)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[4:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[4:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C10,
     Ty Pointer_QTree_Int) : (go_15_goMux_choice_1,C10) [(lizzieLet5_7QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet8_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet11_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet12_1_1_argbuf,Pointer_QTree_Int),
                                                         (lizzieLet13_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [9:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet5_7QNone_Int_1_argbuf_d};
      4'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd2,
                                                               contRet_0_1_argbuf_d};
      4'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_d};
      4'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet8_1_argbuf_d};
      4'd4:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet9_1_argbuf_d};
      4'd5:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet10_1_argbuf_d};
      4'd6:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_d};
      4'd7:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet11_1_argbuf_d};
      4'd8:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet12_1_1_argbuf_d};
      4'd9:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet13_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet13_1_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet11_1_argbuf_r,
          lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_r,
          lizzieLet10_1_argbuf_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet5_7QNone_Int_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                               10'd0);
  
  /* mux (Ty C10,
     Ty Pointer_CT$wmAdd_Int) : (go_15_goMux_choice_2,C10) [(lizzieLet5_5QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (sc_0_6_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QVal_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_4QNode_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int),
                                                            (lizzieLet5_5QError_Int_1_argbuf,Pointer_CT$wmAdd_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [9:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet5_5QNone_Int_1_argbuf_d};
      4'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd2,
                                                               sc_0_6_1_argbuf_d};
      4'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_d};
      4'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_d};
      4'd4:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_d};
      4'd5:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_d};
      4'd6:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_d};
      4'd7:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_d};
      4'd8:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_d};
      4'd9:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet5_5QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet5_5QError_Int_1_argbuf_r,
          lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_r,
          lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_r,
          lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet5_5QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               10'd0);
  
  /* fork (Ty C4) : (go_16_goMux_choice,C4) > [(go_16_goMux_choice_1,C4),
                                          (go_16_goMux_choice_2,C4)] */
  logic [1:0] go_16_goMux_choice_emitted;
  logic [1:0] go_16_goMux_choice_done;
  assign go_16_goMux_choice_1_d = {go_16_goMux_choice_d[2:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[0]))};
  assign go_16_goMux_choice_2_d = {go_16_goMux_choice_d[2:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[1]))};
  assign go_16_goMux_choice_done = (go_16_goMux_choice_emitted | ({go_16_goMux_choice_2_d[0],
                                                                   go_16_goMux_choice_1_d[0]} & {go_16_goMux_choice_2_r,
                                                                                                 go_16_goMux_choice_1_r}));
  assign go_16_goMux_choice_r = (& go_16_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_goMux_choice_emitted <= 2'd0;
    else
      go_16_goMux_choice_emitted <= (go_16_goMux_choice_r ? 2'd0 :
                                     go_16_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_16_goMux_choice_1,C4) [(lizzieLet5_1_1_argbuf,Int#),
                                           (contRet_0_1_1_argbuf,Int#),
                                           (lizzieLet6_1_1_argbuf,Int#),
                                           (lizzieLet5_2_1_argbuf,Int#)] > (srtarg_0_1_goMux_mux,Int#) */
  logic [32:0] srtarg_0_1_goMux_mux_mux;
  logic [3:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet5_1_1_argbuf_d};
      2'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   contRet_0_1_1_argbuf_d};
      2'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet6_1_1_argbuf_d};
      2'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet5_2_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {32'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[32:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_1_d[0])};
  assign go_16_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet5_2_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = (go_16_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz) : (go_16_goMux_choice_2,C4) [(lizzieLet15_4QNone_Bool_1_argbuf,Pointer_CT$wnnz),
                                                      (sc_0_10_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet15_4QVal_Bool_1_argbuf,Pointer_CT$wnnz),
                                                      (lizzieLet15_4QError_Bool_1_argbuf,Pointer_CT$wnnz)] > (scfarg_0_1_goMux_mux,Pointer_CT$wnnz) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [3:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet15_4QNone_Bool_1_argbuf_d};
      2'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd2,
                                                                   sc_0_10_1_argbuf_d};
      2'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet15_4QVal_Bool_1_argbuf_d};
      2'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet15_4QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_2_d[0])};
  assign go_16_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet15_4QError_Bool_1_argbuf_r,
          lizzieLet15_4QVal_Bool_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet15_4QNone_Bool_1_argbuf_r} = (go_16_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                                 4'd0);
  
  /* fork (Ty C5) : (go_17_goMux_choice,C5) > [(go_17_goMux_choice_1,C5),
                                          (go_17_goMux_choice_2,C5)] */
  logic [1:0] go_17_goMux_choice_emitted;
  logic [1:0] go_17_goMux_choice_done;
  assign go_17_goMux_choice_1_d = {go_17_goMux_choice_d[3:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[0]))};
  assign go_17_goMux_choice_2_d = {go_17_goMux_choice_d[3:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[1]))};
  assign go_17_goMux_choice_done = (go_17_goMux_choice_emitted | ({go_17_goMux_choice_2_d[0],
                                                                   go_17_goMux_choice_1_d[0]} & {go_17_goMux_choice_2_r,
                                                                                                 go_17_goMux_choice_1_r}));
  assign go_17_goMux_choice_r = (& go_17_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_goMux_choice_emitted <= 2'd0;
    else
      go_17_goMux_choice_emitted <= (go_17_goMux_choice_r ? 2'd0 :
                                     go_17_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_17_goMux_choice_1,C5) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [4:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_1_d[0])};
  assign go_17_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_17_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Int_Bool) : (go_17_goMux_choice_2,C5) [(lizzieLet17_6QNone_Int_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (sc_0_14_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (es_0_4_2MyFalse_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (es_0_4_2MyTrue_1_argbuf,Pointer_CTmain_map'_Int_Bool),
                                                                   (lizzieLet17_6QError_Int_1_argbuf,Pointer_CTmain_map'_Int_Bool)] > (scfarg_0_2_goMux_mux,Pointer_CTmain_map'_Int_Bool) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [4:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet17_6QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   sc_0_14_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   es_0_4_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   es_0_4_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet17_6QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_2_d[0])};
  assign go_17_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet17_6QError_Int_1_argbuf_r,
          es_0_4_2MyTrue_1_argbuf_r,
          es_0_4_2MyFalse_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet17_6QNone_Int_1_argbuf_r} = (go_17_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                5'd0);
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_1_argbuf,Go),
                                                             (wsm3_1_0,Pointer_QTree_Int),
                                                             (w1sm4_1_1,Pointer_QTree_Int)] > ($wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_1_argbuf_d[0],
                                                                                                                          wsm3_1_0_d[0],
                                                                                                                          w1sm4_1_1_d[0]}), go_1_argbuf_d, wsm3_1_0_d, w1sm4_1_1_d);
  assign {go_1_argbuf_r,
          wsm3_1_0_r,
          w1sm4_1_1_r} = {3 {(\$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_r  && \$wmainTupGo___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon L$wmAdd_Intsbos) : [(go_6_1,Go)] > (go_6_1L$wmAdd_Intsbos,CT$wmAdd_Int) */
  assign go_6_1L$wmAdd_Intsbos_d = L$wmAdd_Intsbos_dc((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(go_6_1L$wmAdd_Intsbos_r && go_6_1L$wmAdd_Intsbos_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (go_6_1L$wmAdd_Intsbos,CT$wmAdd_Int) > (lizzieLet0_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t go_6_1L$wmAdd_Intsbos_bufchan_d;
  logic go_6_1L$wmAdd_Intsbos_bufchan_r;
  assign go_6_1L$wmAdd_Intsbos_r = ((! go_6_1L$wmAdd_Intsbos_bufchan_d[0]) || go_6_1L$wmAdd_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wmAdd_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_6_1L$wmAdd_Intsbos_r)
        go_6_1L$wmAdd_Intsbos_bufchan_d <= go_6_1L$wmAdd_Intsbos_d;
  CT$wmAdd_Int_t go_6_1L$wmAdd_Intsbos_bufchan_buf;
  assign go_6_1L$wmAdd_Intsbos_bufchan_r = (! go_6_1L$wmAdd_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_6_1L$wmAdd_Intsbos_bufchan_buf[0] ? go_6_1L$wmAdd_Intsbos_bufchan_buf :
                                  go_6_1L$wmAdd_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1L$wmAdd_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_6_1L$wmAdd_Intsbos_bufchan_buf[0]))
        go_6_1L$wmAdd_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_6_1L$wmAdd_Intsbos_bufchan_buf[0])))
        go_6_1L$wmAdd_Intsbos_bufchan_buf <= go_6_1L$wmAdd_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int,
      Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) : [(go_6_2_argbuf,Go),
                                                                                                      (wslR_1_argbuf,MyDTInt_Int_Int),
                                                                                                      (w1slS_1_argbuf,Pointer_QTree_Int),
                                                                                                      (w2slT_1_argbuf,Pointer_QTree_Int),
                                                                                                      (lizzieLet14_1_argbuf,Pointer_CT$wmAdd_Int)] > (call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int) */
  assign call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d = TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_dc((& {go_6_2_argbuf_d[0],
                                                                                                                                                                                                                   wslR_1_argbuf_d[0],
                                                                                                                                                                                                                   w1slS_1_argbuf_d[0],
                                                                                                                                                                                                                   w2slT_1_argbuf_d[0],
                                                                                                                                                                                                                   lizzieLet14_1_argbuf_d[0]}), go_6_2_argbuf_d, wslR_1_argbuf_d, w1slS_1_argbuf_d, w2slT_1_argbuf_d, lizzieLet14_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          wslR_1_argbuf_r,
          w1slS_1_argbuf_r,
          w2slT_1_argbuf_r,
          lizzieLet14_1_argbuf_r} = {5 {(call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_r && call_$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int___Pointer_CT$wmAdd_Int_1_d[0])}};
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_main1) : [(go_7_1,Go)] > (go_7_1Dcon_main1,MyDTInt_Bool) */
  assign go_7_1Dcon_main1_d = Dcon_main1_dc((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(go_7_1Dcon_main1_r && go_7_1Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_7_1Dcon_main1,MyDTInt_Bool) > (es_2_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_7_1Dcon_main1_bufchan_d;
  logic go_7_1Dcon_main1_bufchan_r;
  assign go_7_1Dcon_main1_r = ((! go_7_1Dcon_main1_bufchan_d[0]) || go_7_1Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_1Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_7_1Dcon_main1_r)
        go_7_1Dcon_main1_bufchan_d <= go_7_1Dcon_main1_d;
  MyDTInt_Bool_t go_7_1Dcon_main1_bufchan_buf;
  assign go_7_1Dcon_main1_bufchan_r = (! go_7_1Dcon_main1_bufchan_buf[0]);
  assign es_2_1_argbuf_d = (go_7_1Dcon_main1_bufchan_buf[0] ? go_7_1Dcon_main1_bufchan_buf :
                            go_7_1Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_1Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1_argbuf_r && go_7_1Dcon_main1_bufchan_buf[0]))
        go_7_1Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_2_1_argbuf_r) && (! go_7_1Dcon_main1_bufchan_buf[0])))
        go_7_1Dcon_main1_bufchan_buf <= go_7_1Dcon_main1_bufchan_d;
  
  /* dcon (Ty MyDTBool_Bool,
      Dcon Dcon_main2) : [(go_7_2,Go)] > (go_7_2Dcon_main2,MyDTBool_Bool) */
  assign go_7_2Dcon_main2_d = Dcon_main2_dc((& {go_7_2_d[0]}), go_7_2_d);
  assign {go_7_2_r} = {1 {(go_7_2Dcon_main2_r && go_7_2Dcon_main2_d[0])}};
  
  /* buf (Ty MyDTBool_Bool) : (go_7_2Dcon_main2,MyDTBool_Bool) > (es_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t go_7_2Dcon_main2_bufchan_d;
  logic go_7_2Dcon_main2_bufchan_r;
  assign go_7_2Dcon_main2_r = ((! go_7_2Dcon_main2_bufchan_d[0]) || go_7_2Dcon_main2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2Dcon_main2_bufchan_d <= 1'd0;
    else
      if (go_7_2Dcon_main2_r)
        go_7_2Dcon_main2_bufchan_d <= go_7_2Dcon_main2_d;
  MyDTBool_Bool_t go_7_2Dcon_main2_bufchan_buf;
  assign go_7_2Dcon_main2_bufchan_r = (! go_7_2Dcon_main2_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (go_7_2Dcon_main2_bufchan_buf[0] ? go_7_2Dcon_main2_bufchan_buf :
                            go_7_2Dcon_main2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2Dcon_main2_bufchan_buf <= 1'd0;
    else
      if ((es_1_1_argbuf_r && go_7_2Dcon_main2_bufchan_buf[0]))
        go_7_2Dcon_main2_bufchan_buf <= 1'd0;
      else if (((! es_1_1_argbuf_r) && (! go_7_2Dcon_main2_bufchan_buf[0])))
        go_7_2Dcon_main2_bufchan_buf <= go_7_2Dcon_main2_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c+) : [(go_7_3,Go)] > (go_7_3Dcon_$fNumInt_$c+,MyDTInt_Int_Int) */
  assign \go_7_3Dcon_$fNumInt_$c+_d  = \Dcon_$fNumInt_$c+_dc ((& {go_7_3_d[0]}), go_7_3_d);
  assign {go_7_3_r} = {1 {(\go_7_3Dcon_$fNumInt_$c+_r  && \go_7_3Dcon_$fNumInt_$c+_d [0])}};
  
  /* buf (Ty MyDTInt_Int_Int) : (go_7_3Dcon_$fNumInt_$c+,MyDTInt_Int_Int) > (es_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$c+_bufchan_d ;
  logic \go_7_3Dcon_$fNumInt_$c+_bufchan_r ;
  assign \go_7_3Dcon_$fNumInt_$c+_r  = ((! \go_7_3Dcon_$fNumInt_$c+_bufchan_d [0]) || \go_7_3Dcon_$fNumInt_$c+_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_7_3Dcon_$fNumInt_$c+_bufchan_d  <= 1'd0;
    else
      if (\go_7_3Dcon_$fNumInt_$c+_r )
        \go_7_3Dcon_$fNumInt_$c+_bufchan_d  <= \go_7_3Dcon_$fNumInt_$c+_d ;
  MyDTInt_Int_Int_t \go_7_3Dcon_$fNumInt_$c+_bufchan_buf ;
  assign \go_7_3Dcon_$fNumInt_$c+_bufchan_r  = (! \go_7_3Dcon_$fNumInt_$c+_bufchan_buf [0]);
  assign es_4_1_argbuf_d = (\go_7_3Dcon_$fNumInt_$c+_bufchan_buf [0] ? \go_7_3Dcon_$fNumInt_$c+_bufchan_buf  :
                            \go_7_3Dcon_$fNumInt_$c+_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_7_3Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
    else
      if ((es_4_1_argbuf_r && \go_7_3Dcon_$fNumInt_$c+_bufchan_buf [0]))
        \go_7_3Dcon_$fNumInt_$c+_bufchan_buf  <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! \go_7_3Dcon_$fNumInt_$c+_bufchan_buf [0])))
        \go_7_3Dcon_$fNumInt_$c+_bufchan_buf  <= \go_7_3Dcon_$fNumInt_$c+_bufchan_d ;
  
  /* buf (Ty Go) : (go_7_4,Go) > (go_7_4_argbuf,Go) */
  Go_t go_7_4_bufchan_d;
  logic go_7_4_bufchan_r;
  assign go_7_4_r = ((! go_7_4_bufchan_d[0]) || go_7_4_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_4_bufchan_d <= 1'd0;
    else if (go_7_4_r) go_7_4_bufchan_d <= go_7_4_d;
  Go_t go_7_4_bufchan_buf;
  assign go_7_4_bufchan_r = (! go_7_4_bufchan_buf[0]);
  assign go_7_4_argbuf_d = (go_7_4_bufchan_buf[0] ? go_7_4_bufchan_buf :
                            go_7_4_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_4_bufchan_buf <= 1'd0;
    else
      if ((go_7_4_argbuf_r && go_7_4_bufchan_buf[0]))
        go_7_4_bufchan_buf <= 1'd0;
      else if (((! go_7_4_argbuf_r) && (! go_7_4_bufchan_buf[0])))
        go_7_4_bufchan_buf <= go_7_4_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int,
      Dcon TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) : [(go_7_4_argbuf,Go),
                                                                               (es_4_1_argbuf,MyDTInt_Int_Int),
                                                                               (wsm3_1_argbuf,Pointer_QTree_Int),
                                                                               (w1sm4_1_argbuf,Pointer_QTree_Int)] > ($wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1,TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int) */
  assign \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d  = TupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_dc((& {go_7_4_argbuf_d[0],
                                                                                                                                                                  es_4_1_argbuf_d[0],
                                                                                                                                                                  wsm3_1_argbuf_d[0],
                                                                                                                                                                  w1sm4_1_argbuf_d[0]}), go_7_4_argbuf_d, es_4_1_argbuf_d, wsm3_1_argbuf_d, w1sm4_1_argbuf_d);
  assign {go_7_4_argbuf_r,
          es_4_1_argbuf_r,
          wsm3_1_argbuf_r,
          w1sm4_1_argbuf_r} = {4 {(\$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_r  && \$wmAdd_IntTupGo___MyDTInt_Int_Int___Pointer_QTree_Int___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (go_7_5,Go) > (go_7_5_argbuf,Go) */
  Go_t go_7_5_bufchan_d;
  logic go_7_5_bufchan_r;
  assign go_7_5_r = ((! go_7_5_bufchan_d[0]) || go_7_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_5_bufchan_d <= 1'd0;
    else if (go_7_5_r) go_7_5_bufchan_d <= go_7_5_d;
  Go_t go_7_5_bufchan_buf;
  assign go_7_5_bufchan_r = (! go_7_5_bufchan_buf[0]);
  assign go_7_5_argbuf_d = (go_7_5_bufchan_buf[0] ? go_7_5_bufchan_buf :
                            go_7_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_5_bufchan_buf <= 1'd0;
    else
      if ((go_7_5_argbuf_r && go_7_5_bufchan_buf[0]))
        go_7_5_bufchan_buf <= 1'd0;
      else if (((! go_7_5_argbuf_r) && (! go_7_5_bufchan_buf[0])))
        go_7_5_bufchan_buf <= go_7_5_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int,
      Dcon TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int) : [(go_7_5_argbuf,Go),
                                                                        (es_1_1_argbuf,MyDTBool_Bool),
                                                                        (es_2_1_argbuf,MyDTInt_Bool),
                                                                        (es_3_1_argbuf,Pointer_QTree_Int)] > (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1,TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int) */
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d  = TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_dc((& {go_7_5_argbuf_d[0],
                                                                                                                                                            es_1_1_argbuf_d[0],
                                                                                                                                                            es_2_1_argbuf_d[0],
                                                                                                                                                            es_3_1_argbuf_d[0]}), go_7_5_argbuf_d, es_1_1_argbuf_d, es_2_1_argbuf_d, es_3_1_argbuf_d);
  assign {go_7_5_argbuf_r,
          es_1_1_argbuf_r,
          es_2_1_argbuf_r,
          es_3_1_argbuf_r} = {4 {(\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_r  && \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [0])}};
  
  /* buf (Ty Go) : (go_7_6,Go) > (go_7_6_argbuf,Go) */
  Go_t go_7_6_bufchan_d;
  logic go_7_6_bufchan_r;
  assign go_7_6_r = ((! go_7_6_bufchan_d[0]) || go_7_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_6_bufchan_d <= 1'd0;
    else if (go_7_6_r) go_7_6_bufchan_d <= go_7_6_d;
  Go_t go_7_6_bufchan_buf;
  assign go_7_6_bufchan_r = (! go_7_6_bufchan_buf[0]);
  assign go_7_6_argbuf_d = (go_7_6_bufchan_buf[0] ? go_7_6_bufchan_buf :
                            go_7_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_6_bufchan_buf <= 1'd0;
    else
      if ((go_7_6_argbuf_r && go_7_6_bufchan_buf[0]))
        go_7_6_bufchan_buf <= 1'd0;
      else if (((! go_7_6_argbuf_r) && (! go_7_6_bufchan_buf[0])))
        go_7_6_bufchan_buf <= go_7_6_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool,
      Dcon TupGo___Pointer_QTree_Bool) : [(go_7_6_argbuf,Go),
                                          (es_0_1_1_argbuf,Pointer_QTree_Bool)] > ($wnnzTupGo___Pointer_QTree_Bool_1,TupGo___Pointer_QTree_Bool) */
  assign \$wnnzTupGo___Pointer_QTree_Bool_1_d  = TupGo___Pointer_QTree_Bool_dc((& {go_7_6_argbuf_d[0],
                                                                                   es_0_1_1_argbuf_d[0]}), go_7_6_argbuf_d, es_0_1_1_argbuf_d);
  assign {go_7_6_argbuf_r,
          es_0_1_1_argbuf_r} = {2 {(\$wnnzTupGo___Pointer_QTree_Bool_1_r  && \$wnnzTupGo___Pointer_QTree_Bool_1_d [0])}};
  
  /* dcon (Ty CT$wnnz,
      Dcon L$wnnzsbos) : [(go_8_1,Go)] > (go_8_1L$wnnzsbos,CT$wnnz) */
  assign go_8_1L$wnnzsbos_d = L$wnnzsbos_dc((& {go_8_1_d[0]}), go_8_1_d);
  assign {go_8_1_r} = {1 {(go_8_1L$wnnzsbos_r && go_8_1L$wnnzsbos_d[0])}};
  
  /* buf (Ty CT$wnnz) : (go_8_1L$wnnzsbos,CT$wnnz) > (lizzieLet1_1_argbuf,CT$wnnz) */
  CT$wnnz_t go_8_1L$wnnzsbos_bufchan_d;
  logic go_8_1L$wnnzsbos_bufchan_r;
  assign go_8_1L$wnnzsbos_r = ((! go_8_1L$wnnzsbos_bufchan_d[0]) || go_8_1L$wnnzsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_1L$wnnzsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_8_1L$wnnzsbos_r)
        go_8_1L$wnnzsbos_bufchan_d <= go_8_1L$wnnzsbos_d;
  CT$wnnz_t go_8_1L$wnnzsbos_bufchan_buf;
  assign go_8_1L$wnnzsbos_bufchan_r = (! go_8_1L$wnnzsbos_bufchan_buf[0]);
  assign lizzieLet1_1_argbuf_d = (go_8_1L$wnnzsbos_bufchan_buf[0] ? go_8_1L$wnnzsbos_bufchan_buf :
                                  go_8_1L$wnnzsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_8_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet1_1_argbuf_r && go_8_1L$wnnzsbos_bufchan_buf[0]))
        go_8_1L$wnnzsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet1_1_argbuf_r) && (! go_8_1L$wnnzsbos_bufchan_buf[0])))
        go_8_1L$wnnzsbos_bufchan_buf <= go_8_1L$wnnzsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_8_2,Go) > (go_8_2_argbuf,Go) */
  Go_t go_8_2_bufchan_d;
  logic go_8_2_bufchan_r;
  assign go_8_2_r = ((! go_8_2_bufchan_d[0]) || go_8_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_d <= 1'd0;
    else if (go_8_2_r) go_8_2_bufchan_d <= go_8_2_d;
  Go_t go_8_2_bufchan_buf;
  assign go_8_2_bufchan_r = (! go_8_2_bufchan_buf[0]);
  assign go_8_2_argbuf_d = (go_8_2_bufchan_buf[0] ? go_8_2_bufchan_buf :
                            go_8_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_2_bufchan_buf <= 1'd0;
    else
      if ((go_8_2_argbuf_r && go_8_2_bufchan_buf[0]))
        go_8_2_bufchan_buf <= 1'd0;
      else if (((! go_8_2_argbuf_r) && (! go_8_2_bufchan_buf[0])))
        go_8_2_bufchan_buf <= go_8_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) : [(go_8_2_argbuf,Go),
                                                            (wslW_1_argbuf,Pointer_QTree_Bool),
                                                            (lizzieLet7_1_argbuf,Pointer_CT$wnnz)] > (call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1,TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz) */
  assign call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d = TupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_dc((& {go_8_2_argbuf_d[0],
                                                                                                                          wslW_1_argbuf_d[0],
                                                                                                                          lizzieLet7_1_argbuf_d[0]}), go_8_2_argbuf_d, wslW_1_argbuf_d, lizzieLet7_1_argbuf_d);
  assign {go_8_2_argbuf_r,
          wslW_1_argbuf_r,
          lizzieLet7_1_argbuf_r} = {3 {(call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_r && call_$wnnzTupGo___Pointer_QTree_Bool___Pointer_CT$wnnz_1_d[0])}};
  
  /* buf (Ty MyDTBool_Bool) : (isZa8K_2_2,MyDTBool_Bool) > (isZa8K_2_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZa8K_2_2_bufchan_d;
  logic isZa8K_2_2_bufchan_r;
  assign isZa8K_2_2_r = ((! isZa8K_2_2_bufchan_d[0]) || isZa8K_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_2_2_bufchan_d <= 1'd0;
    else if (isZa8K_2_2_r) isZa8K_2_2_bufchan_d <= isZa8K_2_2_d;
  MyDTBool_Bool_t isZa8K_2_2_bufchan_buf;
  assign isZa8K_2_2_bufchan_r = (! isZa8K_2_2_bufchan_buf[0]);
  assign isZa8K_2_2_argbuf_d = (isZa8K_2_2_bufchan_buf[0] ? isZa8K_2_2_bufchan_buf :
                                isZa8K_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZa8K_2_2_argbuf_r && isZa8K_2_2_bufchan_buf[0]))
        isZa8K_2_2_bufchan_buf <= 1'd0;
      else if (((! isZa8K_2_2_argbuf_r) && (! isZa8K_2_2_bufchan_buf[0])))
        isZa8K_2_2_bufchan_buf <= isZa8K_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZa8K_2_destruct,MyDTBool_Bool) > [(isZa8K_2_1,MyDTBool_Bool),
                                                               (isZa8K_2_2,MyDTBool_Bool)] */
  logic [1:0] isZa8K_2_destruct_emitted;
  logic [1:0] isZa8K_2_destruct_done;
  assign isZa8K_2_1_d = (isZa8K_2_destruct_d[0] && (! isZa8K_2_destruct_emitted[0]));
  assign isZa8K_2_2_d = (isZa8K_2_destruct_d[0] && (! isZa8K_2_destruct_emitted[1]));
  assign isZa8K_2_destruct_done = (isZa8K_2_destruct_emitted | ({isZa8K_2_2_d[0],
                                                                 isZa8K_2_1_d[0]} & {isZa8K_2_2_r,
                                                                                     isZa8K_2_1_r}));
  assign isZa8K_2_destruct_r = (& isZa8K_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_2_destruct_emitted <= 2'd0;
    else
      isZa8K_2_destruct_emitted <= (isZa8K_2_destruct_r ? 2'd0 :
                                    isZa8K_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZa8K_3_2,MyDTBool_Bool) > (isZa8K_3_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZa8K_3_2_bufchan_d;
  logic isZa8K_3_2_bufchan_r;
  assign isZa8K_3_2_r = ((! isZa8K_3_2_bufchan_d[0]) || isZa8K_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_3_2_bufchan_d <= 1'd0;
    else if (isZa8K_3_2_r) isZa8K_3_2_bufchan_d <= isZa8K_3_2_d;
  MyDTBool_Bool_t isZa8K_3_2_bufchan_buf;
  assign isZa8K_3_2_bufchan_r = (! isZa8K_3_2_bufchan_buf[0]);
  assign isZa8K_3_2_argbuf_d = (isZa8K_3_2_bufchan_buf[0] ? isZa8K_3_2_bufchan_buf :
                                isZa8K_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZa8K_3_2_argbuf_r && isZa8K_3_2_bufchan_buf[0]))
        isZa8K_3_2_bufchan_buf <= 1'd0;
      else if (((! isZa8K_3_2_argbuf_r) && (! isZa8K_3_2_bufchan_buf[0])))
        isZa8K_3_2_bufchan_buf <= isZa8K_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZa8K_3_destruct,MyDTBool_Bool) > [(isZa8K_3_1,MyDTBool_Bool),
                                                               (isZa8K_3_2,MyDTBool_Bool)] */
  logic [1:0] isZa8K_3_destruct_emitted;
  logic [1:0] isZa8K_3_destruct_done;
  assign isZa8K_3_1_d = (isZa8K_3_destruct_d[0] && (! isZa8K_3_destruct_emitted[0]));
  assign isZa8K_3_2_d = (isZa8K_3_destruct_d[0] && (! isZa8K_3_destruct_emitted[1]));
  assign isZa8K_3_destruct_done = (isZa8K_3_destruct_emitted | ({isZa8K_3_2_d[0],
                                                                 isZa8K_3_1_d[0]} & {isZa8K_3_2_r,
                                                                                     isZa8K_3_1_r}));
  assign isZa8K_3_destruct_r = (& isZa8K_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_3_destruct_emitted <= 2'd0;
    else
      isZa8K_3_destruct_emitted <= (isZa8K_3_destruct_r ? 2'd0 :
                                    isZa8K_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZa8K_4_destruct,MyDTBool_Bool) > (isZa8K_4_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZa8K_4_destruct_bufchan_d;
  logic isZa8K_4_destruct_bufchan_r;
  assign isZa8K_4_destruct_r = ((! isZa8K_4_destruct_bufchan_d[0]) || isZa8K_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZa8K_4_destruct_r)
        isZa8K_4_destruct_bufchan_d <= isZa8K_4_destruct_d;
  MyDTBool_Bool_t isZa8K_4_destruct_bufchan_buf;
  assign isZa8K_4_destruct_bufchan_r = (! isZa8K_4_destruct_bufchan_buf[0]);
  assign isZa8K_4_1_argbuf_d = (isZa8K_4_destruct_bufchan_buf[0] ? isZa8K_4_destruct_bufchan_buf :
                                isZa8K_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZa8K_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZa8K_4_1_argbuf_r && isZa8K_4_destruct_bufchan_buf[0]))
        isZa8K_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZa8K_4_1_argbuf_r) && (! isZa8K_4_destruct_bufchan_buf[0])))
        isZa8K_4_destruct_bufchan_buf <= isZa8K_4_destruct_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet15_1QNode_Bool,QTree_Bool) > [(q1a92_destruct,Pointer_QTree_Bool),
                                                                     (q2a93_destruct,Pointer_QTree_Bool),
                                                                     (q3a94_destruct,Pointer_QTree_Bool),
                                                                     (q4a95_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet15_1QNode_Bool_emitted;
  logic [3:0] lizzieLet15_1QNode_Bool_done;
  assign q1a92_destruct_d = {lizzieLet15_1QNode_Bool_d[18:3],
                             (lizzieLet15_1QNode_Bool_d[0] && (! lizzieLet15_1QNode_Bool_emitted[0]))};
  assign q2a93_destruct_d = {lizzieLet15_1QNode_Bool_d[34:19],
                             (lizzieLet15_1QNode_Bool_d[0] && (! lizzieLet15_1QNode_Bool_emitted[1]))};
  assign q3a94_destruct_d = {lizzieLet15_1QNode_Bool_d[50:35],
                             (lizzieLet15_1QNode_Bool_d[0] && (! lizzieLet15_1QNode_Bool_emitted[2]))};
  assign q4a95_destruct_d = {lizzieLet15_1QNode_Bool_d[66:51],
                             (lizzieLet15_1QNode_Bool_d[0] && (! lizzieLet15_1QNode_Bool_emitted[3]))};
  assign lizzieLet15_1QNode_Bool_done = (lizzieLet15_1QNode_Bool_emitted | ({q4a95_destruct_d[0],
                                                                             q3a94_destruct_d[0],
                                                                             q2a93_destruct_d[0],
                                                                             q1a92_destruct_d[0]} & {q4a95_destruct_r,
                                                                                                     q3a94_destruct_r,
                                                                                                     q2a93_destruct_r,
                                                                                                     q1a92_destruct_r}));
  assign lizzieLet15_1QNode_Bool_r = (& lizzieLet15_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet15_1QNode_Bool_emitted <= (lizzieLet15_1QNode_Bool_r ? 4'd0 :
                                          lizzieLet15_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet15_2,QTree_Bool) (lizzieLet15_1,QTree_Bool) > [(_58,QTree_Bool),
                                                                                 (_57,QTree_Bool),
                                                                                 (lizzieLet15_1QNode_Bool,QTree_Bool),
                                                                                 (_56,QTree_Bool)] */
  logic [3:0] lizzieLet15_1_onehotd;
  always_comb
    if ((lizzieLet15_2_d[0] && lizzieLet15_1_d[0]))
      unique case (lizzieLet15_2_d[2:1])
        2'd0: lizzieLet15_1_onehotd = 4'd1;
        2'd1: lizzieLet15_1_onehotd = 4'd2;
        2'd2: lizzieLet15_1_onehotd = 4'd4;
        2'd3: lizzieLet15_1_onehotd = 4'd8;
        default: lizzieLet15_1_onehotd = 4'd0;
      endcase
    else lizzieLet15_1_onehotd = 4'd0;
  assign _58_d = {lizzieLet15_1_d[66:1], lizzieLet15_1_onehotd[0]};
  assign _57_d = {lizzieLet15_1_d[66:1], lizzieLet15_1_onehotd[1]};
  assign lizzieLet15_1QNode_Bool_d = {lizzieLet15_1_d[66:1],
                                      lizzieLet15_1_onehotd[2]};
  assign _56_d = {lizzieLet15_1_d[66:1], lizzieLet15_1_onehotd[3]};
  assign lizzieLet15_1_r = (| (lizzieLet15_1_onehotd & {_56_r,
                                                        lizzieLet15_1QNode_Bool_r,
                                                        _57_r,
                                                        _58_r}));
  assign lizzieLet15_2_r = lizzieLet15_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet15_3,QTree_Bool) (go_12_goMux_data,Go) > [(lizzieLet15_3QNone_Bool,Go),
                                                                    (lizzieLet15_3QVal_Bool,Go),
                                                                    (lizzieLet15_3QNode_Bool,Go),
                                                                    (lizzieLet15_3QError_Bool,Go)] */
  logic [3:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet15_3_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet15_3_d[2:1])
        2'd0: go_12_goMux_data_onehotd = 4'd1;
        2'd1: go_12_goMux_data_onehotd = 4'd2;
        2'd2: go_12_goMux_data_onehotd = 4'd4;
        2'd3: go_12_goMux_data_onehotd = 4'd8;
        default: go_12_goMux_data_onehotd = 4'd0;
      endcase
    else go_12_goMux_data_onehotd = 4'd0;
  assign lizzieLet15_3QNone_Bool_d = go_12_goMux_data_onehotd[0];
  assign lizzieLet15_3QVal_Bool_d = go_12_goMux_data_onehotd[1];
  assign lizzieLet15_3QNode_Bool_d = go_12_goMux_data_onehotd[2];
  assign lizzieLet15_3QError_Bool_d = go_12_goMux_data_onehotd[3];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {lizzieLet15_3QError_Bool_r,
                                                              lizzieLet15_3QNode_Bool_r,
                                                              lizzieLet15_3QVal_Bool_r,
                                                              lizzieLet15_3QNone_Bool_r}));
  assign lizzieLet15_3_r = go_12_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet15_3QError_Bool,Go) > [(lizzieLet15_3QError_Bool_1,Go),
                                                (lizzieLet15_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet15_3QError_Bool_emitted;
  logic [1:0] lizzieLet15_3QError_Bool_done;
  assign lizzieLet15_3QError_Bool_1_d = (lizzieLet15_3QError_Bool_d[0] && (! lizzieLet15_3QError_Bool_emitted[0]));
  assign lizzieLet15_3QError_Bool_2_d = (lizzieLet15_3QError_Bool_d[0] && (! lizzieLet15_3QError_Bool_emitted[1]));
  assign lizzieLet15_3QError_Bool_done = (lizzieLet15_3QError_Bool_emitted | ({lizzieLet15_3QError_Bool_2_d[0],
                                                                               lizzieLet15_3QError_Bool_1_d[0]} & {lizzieLet15_3QError_Bool_2_r,
                                                                                                                   lizzieLet15_3QError_Bool_1_r}));
  assign lizzieLet15_3QError_Bool_r = (& lizzieLet15_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet15_3QError_Bool_emitted <= (lizzieLet15_3QError_Bool_r ? 2'd0 :
                                           lizzieLet15_3QError_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet15_3QError_Bool_1,Go) > (lizzieLet15_3QError_Bool_1_argbuf,Go) */
  Go_t lizzieLet15_3QError_Bool_1_bufchan_d;
  logic lizzieLet15_3QError_Bool_1_bufchan_r;
  assign lizzieLet15_3QError_Bool_1_r = ((! lizzieLet15_3QError_Bool_1_bufchan_d[0]) || lizzieLet15_3QError_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QError_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QError_Bool_1_r)
        lizzieLet15_3QError_Bool_1_bufchan_d <= lizzieLet15_3QError_Bool_1_d;
  Go_t lizzieLet15_3QError_Bool_1_bufchan_buf;
  assign lizzieLet15_3QError_Bool_1_bufchan_r = (! lizzieLet15_3QError_Bool_1_bufchan_buf[0]);
  assign lizzieLet15_3QError_Bool_1_argbuf_d = (lizzieLet15_3QError_Bool_1_bufchan_buf[0] ? lizzieLet15_3QError_Bool_1_bufchan_buf :
                                                lizzieLet15_3QError_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QError_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QError_Bool_1_argbuf_r && lizzieLet15_3QError_Bool_1_bufchan_buf[0]))
        lizzieLet15_3QError_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QError_Bool_1_argbuf_r) && (! lizzieLet15_3QError_Bool_1_bufchan_buf[0])))
        lizzieLet15_3QError_Bool_1_bufchan_buf <= lizzieLet15_3QError_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet15_3QError_Bool_1_argbuf,Go) > (lizzieLet15_3QError_Bool_1_argbuf_0,Int#) */
  assign lizzieLet15_3QError_Bool_1_argbuf_0_d = {32'd0,
                                                  lizzieLet15_3QError_Bool_1_argbuf_d[0]};
  assign lizzieLet15_3QError_Bool_1_argbuf_r = lizzieLet15_3QError_Bool_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet15_3QError_Bool_1_argbuf_0,Int#) > (lizzieLet5_2_1_argbuf,Int#) */
  \Int#_t  lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d;
  logic lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_r;
  assign lizzieLet15_3QError_Bool_1_argbuf_0_r = ((! lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d[0]) || lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet15_3QError_Bool_1_argbuf_0_r)
        lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d <= lizzieLet15_3QError_Bool_1_argbuf_0_d;
  \Int#_t  lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf;
  assign lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_r = (! lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet5_2_1_argbuf_d = (lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf[0] ? lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf :
                                    lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet5_2_1_argbuf_r && lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf[0]))
        lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet5_2_1_argbuf_r) && (! lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf[0])))
        lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_buf <= lizzieLet15_3QError_Bool_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet15_3QError_Bool_2,Go) > (lizzieLet15_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet15_3QError_Bool_2_bufchan_d;
  logic lizzieLet15_3QError_Bool_2_bufchan_r;
  assign lizzieLet15_3QError_Bool_2_r = ((! lizzieLet15_3QError_Bool_2_bufchan_d[0]) || lizzieLet15_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QError_Bool_2_r)
        lizzieLet15_3QError_Bool_2_bufchan_d <= lizzieLet15_3QError_Bool_2_d;
  Go_t lizzieLet15_3QError_Bool_2_bufchan_buf;
  assign lizzieLet15_3QError_Bool_2_bufchan_r = (! lizzieLet15_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet15_3QError_Bool_2_argbuf_d = (lizzieLet15_3QError_Bool_2_bufchan_buf[0] ? lizzieLet15_3QError_Bool_2_bufchan_buf :
                                                lizzieLet15_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QError_Bool_2_argbuf_r && lizzieLet15_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet15_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QError_Bool_2_argbuf_r) && (! lizzieLet15_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet15_3QError_Bool_2_bufchan_buf <= lizzieLet15_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet15_3QNode_Bool,Go) > (lizzieLet15_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet15_3QNode_Bool_bufchan_d;
  logic lizzieLet15_3QNode_Bool_bufchan_r;
  assign lizzieLet15_3QNode_Bool_r = ((! lizzieLet15_3QNode_Bool_bufchan_d[0]) || lizzieLet15_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QNode_Bool_r)
        lizzieLet15_3QNode_Bool_bufchan_d <= lizzieLet15_3QNode_Bool_d;
  Go_t lizzieLet15_3QNode_Bool_bufchan_buf;
  assign lizzieLet15_3QNode_Bool_bufchan_r = (! lizzieLet15_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet15_3QNode_Bool_1_argbuf_d = (lizzieLet15_3QNode_Bool_bufchan_buf[0] ? lizzieLet15_3QNode_Bool_bufchan_buf :
                                               lizzieLet15_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QNode_Bool_1_argbuf_r && lizzieLet15_3QNode_Bool_bufchan_buf[0]))
        lizzieLet15_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QNode_Bool_1_argbuf_r) && (! lizzieLet15_3QNode_Bool_bufchan_buf[0])))
        lizzieLet15_3QNode_Bool_bufchan_buf <= lizzieLet15_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet15_3QNone_Bool,Go) > [(lizzieLet15_3QNone_Bool_1,Go),
                                               (lizzieLet15_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet15_3QNone_Bool_emitted;
  logic [1:0] lizzieLet15_3QNone_Bool_done;
  assign lizzieLet15_3QNone_Bool_1_d = (lizzieLet15_3QNone_Bool_d[0] && (! lizzieLet15_3QNone_Bool_emitted[0]));
  assign lizzieLet15_3QNone_Bool_2_d = (lizzieLet15_3QNone_Bool_d[0] && (! lizzieLet15_3QNone_Bool_emitted[1]));
  assign lizzieLet15_3QNone_Bool_done = (lizzieLet15_3QNone_Bool_emitted | ({lizzieLet15_3QNone_Bool_2_d[0],
                                                                             lizzieLet15_3QNone_Bool_1_d[0]} & {lizzieLet15_3QNone_Bool_2_r,
                                                                                                                lizzieLet15_3QNone_Bool_1_r}));
  assign lizzieLet15_3QNone_Bool_r = (& lizzieLet15_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet15_3QNone_Bool_emitted <= (lizzieLet15_3QNone_Bool_r ? 2'd0 :
                                          lizzieLet15_3QNone_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet15_3QNone_Bool_1,Go) > (lizzieLet15_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet15_3QNone_Bool_1_bufchan_d;
  logic lizzieLet15_3QNone_Bool_1_bufchan_r;
  assign lizzieLet15_3QNone_Bool_1_r = ((! lizzieLet15_3QNone_Bool_1_bufchan_d[0]) || lizzieLet15_3QNone_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNone_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QNone_Bool_1_r)
        lizzieLet15_3QNone_Bool_1_bufchan_d <= lizzieLet15_3QNone_Bool_1_d;
  Go_t lizzieLet15_3QNone_Bool_1_bufchan_buf;
  assign lizzieLet15_3QNone_Bool_1_bufchan_r = (! lizzieLet15_3QNone_Bool_1_bufchan_buf[0]);
  assign lizzieLet15_3QNone_Bool_1_argbuf_d = (lizzieLet15_3QNone_Bool_1_bufchan_buf[0] ? lizzieLet15_3QNone_Bool_1_bufchan_buf :
                                               lizzieLet15_3QNone_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNone_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QNone_Bool_1_argbuf_r && lizzieLet15_3QNone_Bool_1_bufchan_buf[0]))
        lizzieLet15_3QNone_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QNone_Bool_1_argbuf_r) && (! lizzieLet15_3QNone_Bool_1_bufchan_buf[0])))
        lizzieLet15_3QNone_Bool_1_bufchan_buf <= lizzieLet15_3QNone_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet15_3QNone_Bool_1_argbuf,Go) > (lizzieLet15_3QNone_Bool_1_argbuf_0,Int#) */
  assign lizzieLet15_3QNone_Bool_1_argbuf_0_d = {32'd0,
                                                 lizzieLet15_3QNone_Bool_1_argbuf_d[0]};
  assign lizzieLet15_3QNone_Bool_1_argbuf_r = lizzieLet15_3QNone_Bool_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet15_3QNone_Bool_1_argbuf_0,Int#) > (lizzieLet5_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d;
  logic lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_r;
  assign lizzieLet15_3QNone_Bool_1_argbuf_0_r = ((! lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d[0]) || lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet15_3QNone_Bool_1_argbuf_0_r)
        lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d <= lizzieLet15_3QNone_Bool_1_argbuf_0_d;
  \Int#_t  lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf;
  assign lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_r = (! lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf[0] ? lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf :
                                    lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf[0]))
        lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf[0])))
        lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_buf <= lizzieLet15_3QNone_Bool_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet15_3QNone_Bool_2,Go) > (lizzieLet15_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet15_3QNone_Bool_2_bufchan_d;
  logic lizzieLet15_3QNone_Bool_2_bufchan_r;
  assign lizzieLet15_3QNone_Bool_2_r = ((! lizzieLet15_3QNone_Bool_2_bufchan_d[0]) || lizzieLet15_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QNone_Bool_2_r)
        lizzieLet15_3QNone_Bool_2_bufchan_d <= lizzieLet15_3QNone_Bool_2_d;
  Go_t lizzieLet15_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet15_3QNone_Bool_2_bufchan_r = (! lizzieLet15_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet15_3QNone_Bool_2_argbuf_d = (lizzieLet15_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet15_3QNone_Bool_2_bufchan_buf :
                                               lizzieLet15_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QNone_Bool_2_argbuf_r && lizzieLet15_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet15_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QNone_Bool_2_argbuf_r) && (! lizzieLet15_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet15_3QNone_Bool_2_bufchan_buf <= lizzieLet15_3QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet15_3QNone_Bool_2_argbuf,Go),
                           (lizzieLet29_3Lcall_$wnnz0_1_argbuf,Go),
                           (lizzieLet15_3QVal_Bool_2_argbuf,Go),
                           (lizzieLet15_3QError_Bool_2_argbuf,Go)] > (go_16_goMux_choice,C4) (go_16_goMux_data,Go) */
  logic [3:0] lizzieLet15_3QNone_Bool_2_argbuf_select_d;
  assign lizzieLet15_3QNone_Bool_2_argbuf_select_d = ((| lizzieLet15_3QNone_Bool_2_argbuf_select_q) ? lizzieLet15_3QNone_Bool_2_argbuf_select_q :
                                                      (lizzieLet15_3QNone_Bool_2_argbuf_d[0] ? 4'd1 :
                                                       (lizzieLet29_3Lcall_$wnnz0_1_argbuf_d[0] ? 4'd2 :
                                                        (lizzieLet15_3QVal_Bool_2_argbuf_d[0] ? 4'd4 :
                                                         (lizzieLet15_3QError_Bool_2_argbuf_d[0] ? 4'd8 :
                                                          4'd0)))));
  logic [3:0] lizzieLet15_3QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QNone_Bool_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet15_3QNone_Bool_2_argbuf_select_q <= (lizzieLet15_3QNone_Bool_2_argbuf_done ? 4'd0 :
                                                    lizzieLet15_3QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet15_3QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet15_3QNone_Bool_2_argbuf_emit_q <= (lizzieLet15_3QNone_Bool_2_argbuf_done ? 2'd0 :
                                                  lizzieLet15_3QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet15_3QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet15_3QNone_Bool_2_argbuf_emit_d = (lizzieLet15_3QNone_Bool_2_argbuf_emit_q | ({go_16_goMux_choice_d[0],
                                                                                                go_16_goMux_data_d[0]} & {go_16_goMux_choice_r,
                                                                                                                          go_16_goMux_data_r}));
  logic lizzieLet15_3QNone_Bool_2_argbuf_done;
  assign lizzieLet15_3QNone_Bool_2_argbuf_done = (& lizzieLet15_3QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet15_3QError_Bool_2_argbuf_r,
          lizzieLet15_3QVal_Bool_2_argbuf_r,
          lizzieLet29_3Lcall_$wnnz0_1_argbuf_r,
          lizzieLet15_3QNone_Bool_2_argbuf_r} = (lizzieLet15_3QNone_Bool_2_argbuf_done ? lizzieLet15_3QNone_Bool_2_argbuf_select_d :
                                                 4'd0);
  assign go_16_goMux_data_d = ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet15_3QNone_Bool_2_argbuf_d :
                               ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet29_3Lcall_$wnnz0_1_argbuf_d :
                                ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet15_3QVal_Bool_2_argbuf_d :
                                 ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet15_3QError_Bool_2_argbuf_d :
                                  1'd0))));
  assign go_16_goMux_choice_d = ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet15_3QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet15_3QNone_Bool_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet15_3QVal_Bool,Go) > [(lizzieLet15_3QVal_Bool_1,Go),
                                              (lizzieLet15_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet15_3QVal_Bool_emitted;
  logic [1:0] lizzieLet15_3QVal_Bool_done;
  assign lizzieLet15_3QVal_Bool_1_d = (lizzieLet15_3QVal_Bool_d[0] && (! lizzieLet15_3QVal_Bool_emitted[0]));
  assign lizzieLet15_3QVal_Bool_2_d = (lizzieLet15_3QVal_Bool_d[0] && (! lizzieLet15_3QVal_Bool_emitted[1]));
  assign lizzieLet15_3QVal_Bool_done = (lizzieLet15_3QVal_Bool_emitted | ({lizzieLet15_3QVal_Bool_2_d[0],
                                                                           lizzieLet15_3QVal_Bool_1_d[0]} & {lizzieLet15_3QVal_Bool_2_r,
                                                                                                             lizzieLet15_3QVal_Bool_1_r}));
  assign lizzieLet15_3QVal_Bool_r = (& lizzieLet15_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet15_3QVal_Bool_emitted <= (lizzieLet15_3QVal_Bool_r ? 2'd0 :
                                         lizzieLet15_3QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet15_3QVal_Bool_1,Go) > (lizzieLet15_3QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet15_3QVal_Bool_1_bufchan_d;
  logic lizzieLet15_3QVal_Bool_1_bufchan_r;
  assign lizzieLet15_3QVal_Bool_1_r = ((! lizzieLet15_3QVal_Bool_1_bufchan_d[0]) || lizzieLet15_3QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QVal_Bool_1_r)
        lizzieLet15_3QVal_Bool_1_bufchan_d <= lizzieLet15_3QVal_Bool_1_d;
  Go_t lizzieLet15_3QVal_Bool_1_bufchan_buf;
  assign lizzieLet15_3QVal_Bool_1_bufchan_r = (! lizzieLet15_3QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet15_3QVal_Bool_1_argbuf_d = (lizzieLet15_3QVal_Bool_1_bufchan_buf[0] ? lizzieLet15_3QVal_Bool_1_bufchan_buf :
                                              lizzieLet15_3QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QVal_Bool_1_argbuf_r && lizzieLet15_3QVal_Bool_1_bufchan_buf[0]))
        lizzieLet15_3QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QVal_Bool_1_argbuf_r) && (! lizzieLet15_3QVal_Bool_1_bufchan_buf[0])))
        lizzieLet15_3QVal_Bool_1_bufchan_buf <= lizzieLet15_3QVal_Bool_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet15_3QVal_Bool_1_argbuf,Go) > (lizzieLet15_3QVal_Bool_1_argbuf_1,Int#) */
  assign lizzieLet15_3QVal_Bool_1_argbuf_1_d = {32'd1,
                                                lizzieLet15_3QVal_Bool_1_argbuf_d[0]};
  assign lizzieLet15_3QVal_Bool_1_argbuf_r = lizzieLet15_3QVal_Bool_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet15_3QVal_Bool_1_argbuf_1,Int#) > (lizzieLet6_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d;
  logic lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_r;
  assign lizzieLet15_3QVal_Bool_1_argbuf_1_r = ((! lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d[0]) || lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet15_3QVal_Bool_1_argbuf_1_r)
        lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d <= lizzieLet15_3QVal_Bool_1_argbuf_1_d;
  \Int#_t  lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf;
  assign lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_r = (! lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf[0] ? lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf :
                                    lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf[0]))
        lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf[0])))
        lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_buf <= lizzieLet15_3QVal_Bool_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet15_3QVal_Bool_2,Go) > (lizzieLet15_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet15_3QVal_Bool_2_bufchan_d;
  logic lizzieLet15_3QVal_Bool_2_bufchan_r;
  assign lizzieLet15_3QVal_Bool_2_r = ((! lizzieLet15_3QVal_Bool_2_bufchan_d[0]) || lizzieLet15_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet15_3QVal_Bool_2_r)
        lizzieLet15_3QVal_Bool_2_bufchan_d <= lizzieLet15_3QVal_Bool_2_d;
  Go_t lizzieLet15_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet15_3QVal_Bool_2_bufchan_r = (! lizzieLet15_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet15_3QVal_Bool_2_argbuf_d = (lizzieLet15_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet15_3QVal_Bool_2_bufchan_buf :
                                              lizzieLet15_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet15_3QVal_Bool_2_argbuf_r && lizzieLet15_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet15_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet15_3QVal_Bool_2_argbuf_r) && (! lizzieLet15_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet15_3QVal_Bool_2_bufchan_buf <= lizzieLet15_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CT$wnnz) : (lizzieLet15_4,QTree_Bool) (sc_0_1_goMux_mux,Pointer_CT$wnnz) > [(lizzieLet15_4QNone_Bool,Pointer_CT$wnnz),
                                                                                              (lizzieLet15_4QVal_Bool,Pointer_CT$wnnz),
                                                                                              (lizzieLet15_4QNode_Bool,Pointer_CT$wnnz),
                                                                                              (lizzieLet15_4QError_Bool,Pointer_CT$wnnz)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet15_4_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet15_4_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet15_4QNone_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet15_4QVal_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet15_4QNode_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet15_4QError_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                       sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet15_4QError_Bool_r,
                                                              lizzieLet15_4QNode_Bool_r,
                                                              lizzieLet15_4QVal_Bool_r,
                                                              lizzieLet15_4QNone_Bool_r}));
  assign lizzieLet15_4_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet15_4QError_Bool,Pointer_CT$wnnz) > (lizzieLet15_4QError_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet15_4QError_Bool_bufchan_d;
  logic lizzieLet15_4QError_Bool_bufchan_r;
  assign lizzieLet15_4QError_Bool_r = ((! lizzieLet15_4QError_Bool_bufchan_d[0]) || lizzieLet15_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet15_4QError_Bool_r)
        lizzieLet15_4QError_Bool_bufchan_d <= lizzieLet15_4QError_Bool_d;
  Pointer_CT$wnnz_t lizzieLet15_4QError_Bool_bufchan_buf;
  assign lizzieLet15_4QError_Bool_bufchan_r = (! lizzieLet15_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet15_4QError_Bool_1_argbuf_d = (lizzieLet15_4QError_Bool_bufchan_buf[0] ? lizzieLet15_4QError_Bool_bufchan_buf :
                                                lizzieLet15_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet15_4QError_Bool_1_argbuf_r && lizzieLet15_4QError_Bool_bufchan_buf[0]))
        lizzieLet15_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet15_4QError_Bool_1_argbuf_r) && (! lizzieLet15_4QError_Bool_bufchan_buf[0])))
        lizzieLet15_4QError_Bool_bufchan_buf <= lizzieLet15_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz3) : [(lizzieLet15_4QNode_Bool,Pointer_CT$wnnz),
                            (q4a95_destruct,Pointer_QTree_Bool),
                            (q3a94_destruct,Pointer_QTree_Bool),
                            (q2a93_destruct,Pointer_QTree_Bool)] > (lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3,CT$wnnz) */
  assign lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_d = Lcall_$wnnz3_dc((& {lizzieLet15_4QNode_Bool_d[0],
                                                                                            q4a95_destruct_d[0],
                                                                                            q3a94_destruct_d[0],
                                                                                            q2a93_destruct_d[0]}), lizzieLet15_4QNode_Bool_d, q4a95_destruct_d, q3a94_destruct_d, q2a93_destruct_d);
  assign {lizzieLet15_4QNode_Bool_r,
          q4a95_destruct_r,
          q3a94_destruct_r,
          q2a93_destruct_r} = {4 {(lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_r && lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3,CT$wnnz) > (lizzieLet16_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d;
  logic lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_r;
  assign lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_r = ((! lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d[0]) || lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d <= {115'd0,
                                                                               1'd0};
    else
      if (lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_r)
        lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d <= lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_d;
  CT$wnnz_t lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_r = (! lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf :
                                   lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf <= {115'd0,
                                                                                   1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_buf <= lizzieLet15_4QNode_Bool_1q4a95_1q3a94_1q2a93_1Lcall_$wnnz3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet15_4QNone_Bool,Pointer_CT$wnnz) > (lizzieLet15_4QNone_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet15_4QNone_Bool_bufchan_d;
  logic lizzieLet15_4QNone_Bool_bufchan_r;
  assign lizzieLet15_4QNone_Bool_r = ((! lizzieLet15_4QNone_Bool_bufchan_d[0]) || lizzieLet15_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet15_4QNone_Bool_r)
        lizzieLet15_4QNone_Bool_bufchan_d <= lizzieLet15_4QNone_Bool_d;
  Pointer_CT$wnnz_t lizzieLet15_4QNone_Bool_bufchan_buf;
  assign lizzieLet15_4QNone_Bool_bufchan_r = (! lizzieLet15_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet15_4QNone_Bool_1_argbuf_d = (lizzieLet15_4QNone_Bool_bufchan_buf[0] ? lizzieLet15_4QNone_Bool_bufchan_buf :
                                               lizzieLet15_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet15_4QNone_Bool_1_argbuf_r && lizzieLet15_4QNone_Bool_bufchan_buf[0]))
        lizzieLet15_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet15_4QNone_Bool_1_argbuf_r) && (! lizzieLet15_4QNone_Bool_bufchan_buf[0])))
        lizzieLet15_4QNone_Bool_bufchan_buf <= lizzieLet15_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (lizzieLet15_4QVal_Bool,Pointer_CT$wnnz) > (lizzieLet15_4QVal_Bool_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t lizzieLet15_4QVal_Bool_bufchan_d;
  logic lizzieLet15_4QVal_Bool_bufchan_r;
  assign lizzieLet15_4QVal_Bool_r = ((! lizzieLet15_4QVal_Bool_bufchan_d[0]) || lizzieLet15_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet15_4QVal_Bool_r)
        lizzieLet15_4QVal_Bool_bufchan_d <= lizzieLet15_4QVal_Bool_d;
  Pointer_CT$wnnz_t lizzieLet15_4QVal_Bool_bufchan_buf;
  assign lizzieLet15_4QVal_Bool_bufchan_r = (! lizzieLet15_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet15_4QVal_Bool_1_argbuf_d = (lizzieLet15_4QVal_Bool_bufchan_buf[0] ? lizzieLet15_4QVal_Bool_bufchan_buf :
                                              lizzieLet15_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet15_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet15_4QVal_Bool_1_argbuf_r && lizzieLet15_4QVal_Bool_bufchan_buf[0]))
        lizzieLet15_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet15_4QVal_Bool_1_argbuf_r) && (! lizzieLet15_4QVal_Bool_bufchan_buf[0])))
        lizzieLet15_4QVal_Bool_bufchan_buf <= lizzieLet15_4QVal_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet17_1QNode_Int,QTree_Int) > [(q1a8O_destruct,Pointer_QTree_Int),
                                                                  (q2a8P_destruct,Pointer_QTree_Int),
                                                                  (q3a8Q_destruct,Pointer_QTree_Int),
                                                                  (q4a8R_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet17_1QNode_Int_emitted;
  logic [3:0] lizzieLet17_1QNode_Int_done;
  assign q1a8O_destruct_d = {lizzieLet17_1QNode_Int_d[18:3],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[0]))};
  assign q2a8P_destruct_d = {lizzieLet17_1QNode_Int_d[34:19],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[1]))};
  assign q3a8Q_destruct_d = {lizzieLet17_1QNode_Int_d[50:35],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[2]))};
  assign q4a8R_destruct_d = {lizzieLet17_1QNode_Int_d[66:51],
                             (lizzieLet17_1QNode_Int_d[0] && (! lizzieLet17_1QNode_Int_emitted[3]))};
  assign lizzieLet17_1QNode_Int_done = (lizzieLet17_1QNode_Int_emitted | ({q4a8R_destruct_d[0],
                                                                           q3a8Q_destruct_d[0],
                                                                           q2a8P_destruct_d[0],
                                                                           q1a8O_destruct_d[0]} & {q4a8R_destruct_r,
                                                                                                   q3a8Q_destruct_r,
                                                                                                   q2a8P_destruct_r,
                                                                                                   q1a8O_destruct_r}));
  assign lizzieLet17_1QNode_Int_r = (& lizzieLet17_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet17_1QNode_Int_emitted <= (lizzieLet17_1QNode_Int_r ? 4'd0 :
                                         lizzieLet17_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet17_1QVal_Int,QTree_Int) > [(va8N_destruct,Int)] */
  assign va8N_destruct_d = {lizzieLet17_1QVal_Int_d[34:3],
                            lizzieLet17_1QVal_Int_d[0]};
  assign lizzieLet17_1QVal_Int_r = va8N_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet17_2,QTree_Int) (lizzieLet17_1,QTree_Int) > [(_55,QTree_Int),
                                                                              (lizzieLet17_1QVal_Int,QTree_Int),
                                                                              (lizzieLet17_1QNode_Int,QTree_Int),
                                                                              (_54,QTree_Int)] */
  logic [3:0] lizzieLet17_1_onehotd;
  always_comb
    if ((lizzieLet17_2_d[0] && lizzieLet17_1_d[0]))
      unique case (lizzieLet17_2_d[2:1])
        2'd0: lizzieLet17_1_onehotd = 4'd1;
        2'd1: lizzieLet17_1_onehotd = 4'd2;
        2'd2: lizzieLet17_1_onehotd = 4'd4;
        2'd3: lizzieLet17_1_onehotd = 4'd8;
        default: lizzieLet17_1_onehotd = 4'd0;
      endcase
    else lizzieLet17_1_onehotd = 4'd0;
  assign _55_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[0]};
  assign lizzieLet17_1QVal_Int_d = {lizzieLet17_1_d[66:1],
                                    lizzieLet17_1_onehotd[1]};
  assign lizzieLet17_1QNode_Int_d = {lizzieLet17_1_d[66:1],
                                     lizzieLet17_1_onehotd[2]};
  assign _54_d = {lizzieLet17_1_d[66:1], lizzieLet17_1_onehotd[3]};
  assign lizzieLet17_1_r = (| (lizzieLet17_1_onehotd & {_54_r,
                                                        lizzieLet17_1QNode_Int_r,
                                                        lizzieLet17_1QVal_Int_r,
                                                        _55_r}));
  assign lizzieLet17_2_r = lizzieLet17_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet17_3,QTree_Int) (ga8L_goMux_mux,MyDTInt_Bool) > [(_53,MyDTInt_Bool),
                                                                                     (lizzieLet17_3QVal_Int,MyDTInt_Bool),
                                                                                     (lizzieLet17_3QNode_Int,MyDTInt_Bool),
                                                                                     (_52,MyDTInt_Bool)] */
  logic [3:0] ga8L_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_3_d[0] && ga8L_goMux_mux_d[0]))
      unique case (lizzieLet17_3_d[2:1])
        2'd0: ga8L_goMux_mux_onehotd = 4'd1;
        2'd1: ga8L_goMux_mux_onehotd = 4'd2;
        2'd2: ga8L_goMux_mux_onehotd = 4'd4;
        2'd3: ga8L_goMux_mux_onehotd = 4'd8;
        default: ga8L_goMux_mux_onehotd = 4'd0;
      endcase
    else ga8L_goMux_mux_onehotd = 4'd0;
  assign _53_d = ga8L_goMux_mux_onehotd[0];
  assign lizzieLet17_3QVal_Int_d = ga8L_goMux_mux_onehotd[1];
  assign lizzieLet17_3QNode_Int_d = ga8L_goMux_mux_onehotd[2];
  assign _52_d = ga8L_goMux_mux_onehotd[3];
  assign ga8L_goMux_mux_r = (| (ga8L_goMux_mux_onehotd & {_52_r,
                                                          lizzieLet17_3QNode_Int_r,
                                                          lizzieLet17_3QVal_Int_r,
                                                          _53_r}));
  assign lizzieLet17_3_r = ga8L_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet17_3QNode_Int,MyDTInt_Bool) > [(lizzieLet17_3QNode_Int_1,MyDTInt_Bool),
                                                                  (lizzieLet17_3QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet17_3QNode_Int_emitted;
  logic [1:0] lizzieLet17_3QNode_Int_done;
  assign lizzieLet17_3QNode_Int_1_d = (lizzieLet17_3QNode_Int_d[0] && (! lizzieLet17_3QNode_Int_emitted[0]));
  assign lizzieLet17_3QNode_Int_2_d = (lizzieLet17_3QNode_Int_d[0] && (! lizzieLet17_3QNode_Int_emitted[1]));
  assign lizzieLet17_3QNode_Int_done = (lizzieLet17_3QNode_Int_emitted | ({lizzieLet17_3QNode_Int_2_d[0],
                                                                           lizzieLet17_3QNode_Int_1_d[0]} & {lizzieLet17_3QNode_Int_2_r,
                                                                                                             lizzieLet17_3QNode_Int_1_r}));
  assign lizzieLet17_3QNode_Int_r = (& lizzieLet17_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_3QNode_Int_emitted <= (lizzieLet17_3QNode_Int_r ? 2'd0 :
                                         lizzieLet17_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_3QNode_Int_2,MyDTInt_Bool) > (lizzieLet17_3QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_2_bufchan_d;
  logic lizzieLet17_3QNode_Int_2_bufchan_r;
  assign lizzieLet17_3QNode_Int_2_r = ((! lizzieLet17_3QNode_Int_2_bufchan_d[0]) || lizzieLet17_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_3QNode_Int_2_r)
        lizzieLet17_3QNode_Int_2_bufchan_d <= lizzieLet17_3QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet17_3QNode_Int_2_bufchan_buf;
  assign lizzieLet17_3QNode_Int_2_bufchan_r = (! lizzieLet17_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_3QNode_Int_2_argbuf_d = (lizzieLet17_3QNode_Int_2_bufchan_buf[0] ? lizzieLet17_3QNode_Int_2_bufchan_buf :
                                              lizzieLet17_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_3QNode_Int_2_argbuf_r && lizzieLet17_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_3QNode_Int_2_argbuf_r) && (! lizzieLet17_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_3QNode_Int_2_bufchan_buf <= lizzieLet17_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet17_3QVal_Int,MyDTInt_Bool) > (lizzieLet17_3QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet17_3QVal_Int_bufchan_d;
  logic lizzieLet17_3QVal_Int_bufchan_r;
  assign lizzieLet17_3QVal_Int_r = ((! lizzieLet17_3QVal_Int_bufchan_d[0]) || lizzieLet17_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_3QVal_Int_r)
        lizzieLet17_3QVal_Int_bufchan_d <= lizzieLet17_3QVal_Int_d;
  MyDTInt_Bool_t lizzieLet17_3QVal_Int_bufchan_buf;
  assign lizzieLet17_3QVal_Int_bufchan_r = (! lizzieLet17_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_3QVal_Int_1_argbuf_d = (lizzieLet17_3QVal_Int_bufchan_buf[0] ? lizzieLet17_3QVal_Int_bufchan_buf :
                                             lizzieLet17_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_3QVal_Int_1_argbuf_r && lizzieLet17_3QVal_Int_bufchan_buf[0]))
        lizzieLet17_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_3QVal_Int_1_argbuf_r) && (! lizzieLet17_3QVal_Int_bufchan_buf[0])))
        lizzieLet17_3QVal_Int_bufchan_buf <= lizzieLet17_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet17_4,QTree_Int) (go_13_goMux_data,Go) > [(lizzieLet17_4QNone_Int,Go),
                                                                   (lizzieLet17_4QVal_Int,Go),
                                                                   (lizzieLet17_4QNode_Int,Go),
                                                                   (lizzieLet17_4QError_Int,Go)] */
  logic [3:0] go_13_goMux_data_onehotd;
  always_comb
    if ((lizzieLet17_4_d[0] && go_13_goMux_data_d[0]))
      unique case (lizzieLet17_4_d[2:1])
        2'd0: go_13_goMux_data_onehotd = 4'd1;
        2'd1: go_13_goMux_data_onehotd = 4'd2;
        2'd2: go_13_goMux_data_onehotd = 4'd4;
        2'd3: go_13_goMux_data_onehotd = 4'd8;
        default: go_13_goMux_data_onehotd = 4'd0;
      endcase
    else go_13_goMux_data_onehotd = 4'd0;
  assign lizzieLet17_4QNone_Int_d = go_13_goMux_data_onehotd[0];
  assign lizzieLet17_4QVal_Int_d = go_13_goMux_data_onehotd[1];
  assign lizzieLet17_4QNode_Int_d = go_13_goMux_data_onehotd[2];
  assign lizzieLet17_4QError_Int_d = go_13_goMux_data_onehotd[3];
  assign go_13_goMux_data_r = (| (go_13_goMux_data_onehotd & {lizzieLet17_4QError_Int_r,
                                                              lizzieLet17_4QNode_Int_r,
                                                              lizzieLet17_4QVal_Int_r,
                                                              lizzieLet17_4QNone_Int_r}));
  assign lizzieLet17_4_r = go_13_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet17_4QError_Int,Go) > [(lizzieLet17_4QError_Int_1,Go),
                                               (lizzieLet17_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet17_4QError_Int_emitted;
  logic [1:0] lizzieLet17_4QError_Int_done;
  assign lizzieLet17_4QError_Int_1_d = (lizzieLet17_4QError_Int_d[0] && (! lizzieLet17_4QError_Int_emitted[0]));
  assign lizzieLet17_4QError_Int_2_d = (lizzieLet17_4QError_Int_d[0] && (! lizzieLet17_4QError_Int_emitted[1]));
  assign lizzieLet17_4QError_Int_done = (lizzieLet17_4QError_Int_emitted | ({lizzieLet17_4QError_Int_2_d[0],
                                                                             lizzieLet17_4QError_Int_1_d[0]} & {lizzieLet17_4QError_Int_2_r,
                                                                                                                lizzieLet17_4QError_Int_1_r}));
  assign lizzieLet17_4QError_Int_r = (& lizzieLet17_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet17_4QError_Int_emitted <= (lizzieLet17_4QError_Int_r ? 2'd0 :
                                          lizzieLet17_4QError_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet17_4QError_Int_1,Go)] > (lizzieLet17_4QError_Int_1QError_Bool,QTree_Bool) */
  assign lizzieLet17_4QError_Int_1QError_Bool_d = QError_Bool_dc((& {lizzieLet17_4QError_Int_1_d[0]}), lizzieLet17_4QError_Int_1_d);
  assign {lizzieLet17_4QError_Int_1_r} = {1 {(lizzieLet17_4QError_Int_1QError_Bool_r && lizzieLet17_4QError_Int_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet17_4QError_Int_1QError_Bool,QTree_Bool) > (lizzieLet22_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet17_4QError_Int_1QError_Bool_bufchan_d;
  logic lizzieLet17_4QError_Int_1QError_Bool_bufchan_r;
  assign lizzieLet17_4QError_Int_1QError_Bool_r = ((! lizzieLet17_4QError_Int_1QError_Bool_bufchan_d[0]) || lizzieLet17_4QError_Int_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QError_Int_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_4QError_Int_1QError_Bool_r)
        lizzieLet17_4QError_Int_1QError_Bool_bufchan_d <= lizzieLet17_4QError_Int_1QError_Bool_d;
  QTree_Bool_t lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf;
  assign lizzieLet17_4QError_Int_1QError_Bool_bufchan_r = (! lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf[0] ? lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf :
                                   lizzieLet17_4QError_Int_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf[0]))
        lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf[0])))
        lizzieLet17_4QError_Int_1QError_Bool_bufchan_buf <= lizzieLet17_4QError_Int_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QError_Int_2,Go) > (lizzieLet17_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet17_4QError_Int_2_bufchan_d;
  logic lizzieLet17_4QError_Int_2_bufchan_r;
  assign lizzieLet17_4QError_Int_2_r = ((! lizzieLet17_4QError_Int_2_bufchan_d[0]) || lizzieLet17_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QError_Int_2_r)
        lizzieLet17_4QError_Int_2_bufchan_d <= lizzieLet17_4QError_Int_2_d;
  Go_t lizzieLet17_4QError_Int_2_bufchan_buf;
  assign lizzieLet17_4QError_Int_2_bufchan_r = (! lizzieLet17_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet17_4QError_Int_2_argbuf_d = (lizzieLet17_4QError_Int_2_bufchan_buf[0] ? lizzieLet17_4QError_Int_2_bufchan_buf :
                                               lizzieLet17_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QError_Int_2_argbuf_r && lizzieLet17_4QError_Int_2_bufchan_buf[0]))
        lizzieLet17_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QError_Int_2_argbuf_r) && (! lizzieLet17_4QError_Int_2_bufchan_buf[0])))
        lizzieLet17_4QError_Int_2_bufchan_buf <= lizzieLet17_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QNode_Int,Go) > (lizzieLet17_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet17_4QNode_Int_bufchan_d;
  logic lizzieLet17_4QNode_Int_bufchan_r;
  assign lizzieLet17_4QNode_Int_r = ((! lizzieLet17_4QNode_Int_bufchan_d[0]) || lizzieLet17_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QNode_Int_r)
        lizzieLet17_4QNode_Int_bufchan_d <= lizzieLet17_4QNode_Int_d;
  Go_t lizzieLet17_4QNode_Int_bufchan_buf;
  assign lizzieLet17_4QNode_Int_bufchan_r = (! lizzieLet17_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet17_4QNode_Int_1_argbuf_d = (lizzieLet17_4QNode_Int_bufchan_buf[0] ? lizzieLet17_4QNode_Int_bufchan_buf :
                                              lizzieLet17_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QNode_Int_1_argbuf_r && lizzieLet17_4QNode_Int_bufchan_buf[0]))
        lizzieLet17_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QNode_Int_1_argbuf_r) && (! lizzieLet17_4QNode_Int_bufchan_buf[0])))
        lizzieLet17_4QNode_Int_bufchan_buf <= lizzieLet17_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet17_4QNone_Int,Go) > [(lizzieLet17_4QNone_Int_1,Go),
                                              (lizzieLet17_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet17_4QNone_Int_emitted;
  logic [1:0] lizzieLet17_4QNone_Int_done;
  assign lizzieLet17_4QNone_Int_1_d = (lizzieLet17_4QNone_Int_d[0] && (! lizzieLet17_4QNone_Int_emitted[0]));
  assign lizzieLet17_4QNone_Int_2_d = (lizzieLet17_4QNone_Int_d[0] && (! lizzieLet17_4QNone_Int_emitted[1]));
  assign lizzieLet17_4QNone_Int_done = (lizzieLet17_4QNone_Int_emitted | ({lizzieLet17_4QNone_Int_2_d[0],
                                                                           lizzieLet17_4QNone_Int_1_d[0]} & {lizzieLet17_4QNone_Int_2_r,
                                                                                                             lizzieLet17_4QNone_Int_1_r}));
  assign lizzieLet17_4QNone_Int_r = (& lizzieLet17_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet17_4QNone_Int_emitted <= (lizzieLet17_4QNone_Int_r ? 2'd0 :
                                         lizzieLet17_4QNone_Int_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet17_4QNone_Int_1,Go)] > (lizzieLet17_4QNone_Int_1QNone_Bool,QTree_Bool) */
  assign lizzieLet17_4QNone_Int_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet17_4QNone_Int_1_d[0]}), lizzieLet17_4QNone_Int_1_d);
  assign {lizzieLet17_4QNone_Int_1_r} = {1 {(lizzieLet17_4QNone_Int_1QNone_Bool_r && lizzieLet17_4QNone_Int_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet17_4QNone_Int_1QNone_Bool,QTree_Bool) > (lizzieLet18_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d;
  logic lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_r;
  assign lizzieLet17_4QNone_Int_1QNone_Bool_r = ((! lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d[0]) || lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet17_4QNone_Int_1QNone_Bool_r)
        lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d <= lizzieLet17_4QNone_Int_1QNone_Bool_d;
  QTree_Bool_t lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf;
  assign lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_r = (! lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf[0] ? lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf :
                                   lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf[0]))
        lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf[0])))
        lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_buf <= lizzieLet17_4QNone_Int_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet17_4QNone_Int_2,Go) > (lizzieLet17_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet17_4QNone_Int_2_bufchan_d;
  logic lizzieLet17_4QNone_Int_2_bufchan_r;
  assign lizzieLet17_4QNone_Int_2_r = ((! lizzieLet17_4QNone_Int_2_bufchan_d[0]) || lizzieLet17_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QNone_Int_2_r)
        lizzieLet17_4QNone_Int_2_bufchan_d <= lizzieLet17_4QNone_Int_2_d;
  Go_t lizzieLet17_4QNone_Int_2_bufchan_buf;
  assign lizzieLet17_4QNone_Int_2_bufchan_r = (! lizzieLet17_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet17_4QNone_Int_2_argbuf_d = (lizzieLet17_4QNone_Int_2_bufchan_buf[0] ? lizzieLet17_4QNone_Int_2_bufchan_buf :
                                              lizzieLet17_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QNone_Int_2_argbuf_r && lizzieLet17_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet17_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QNone_Int_2_argbuf_r) && (! lizzieLet17_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet17_4QNone_Int_2_bufchan_buf <= lizzieLet17_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet17_4QNone_Int_2_argbuf,Go),
                           (lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf,Go),
                           (es_0_4_1MyFalse_1_argbuf,Go),
                           (es_0_4_1MyTrue_2_argbuf,Go),
                           (lizzieLet17_4QError_Int_2_argbuf,Go)] > (go_17_goMux_choice,C5) (go_17_goMux_data,Go) */
  logic [4:0] lizzieLet17_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet17_4QNone_Int_2_argbuf_select_d = ((| lizzieLet17_4QNone_Int_2_argbuf_select_q) ? lizzieLet17_4QNone_Int_2_argbuf_select_q :
                                                     (lizzieLet17_4QNone_Int_2_argbuf_d[0] ? 5'd1 :
                                                      (\lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_d [0] ? 5'd2 :
                                                       (es_0_4_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                        (es_0_4_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                         (lizzieLet17_4QError_Int_2_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] lizzieLet17_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet17_4QNone_Int_2_argbuf_select_q <= (lizzieLet17_4QNone_Int_2_argbuf_done ? 5'd0 :
                                                   lizzieLet17_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet17_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet17_4QNone_Int_2_argbuf_emit_q <= (lizzieLet17_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                 lizzieLet17_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet17_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet17_4QNone_Int_2_argbuf_emit_d = (lizzieLet17_4QNone_Int_2_argbuf_emit_q | ({go_17_goMux_choice_d[0],
                                                                                              go_17_goMux_data_d[0]} & {go_17_goMux_choice_r,
                                                                                                                        go_17_goMux_data_r}));
  logic lizzieLet17_4QNone_Int_2_argbuf_done;
  assign lizzieLet17_4QNone_Int_2_argbuf_done = (& lizzieLet17_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet17_4QError_Int_2_argbuf_r,
          es_0_4_1MyTrue_2_argbuf_r,
          es_0_4_1MyFalse_1_argbuf_r,
          \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_r ,
          lizzieLet17_4QNone_Int_2_argbuf_r} = (lizzieLet17_4QNone_Int_2_argbuf_done ? lizzieLet17_4QNone_Int_2_argbuf_select_d :
                                                5'd0);
  assign go_17_goMux_data_d = ((lizzieLet17_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_4QNone_Int_2_argbuf_d :
                               ((lizzieLet17_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_d  :
                                ((lizzieLet17_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_4_1MyFalse_1_argbuf_d :
                                 ((lizzieLet17_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? es_0_4_1MyTrue_2_argbuf_d :
                                  ((lizzieLet17_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet17_4QError_Int_2_argbuf_d :
                                   1'd0)))));
  assign go_17_goMux_choice_d = ((lizzieLet17_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet17_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet17_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet17_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet17_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet17_4QNone_Int_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet17_4QVal_Int,Go) > [(lizzieLet17_4QVal_Int_1,Go),
                                             (lizzieLet17_4QVal_Int_2,Go),
                                             (lizzieLet17_4QVal_Int_3,Go)] */
  logic [2:0] lizzieLet17_4QVal_Int_emitted;
  logic [2:0] lizzieLet17_4QVal_Int_done;
  assign lizzieLet17_4QVal_Int_1_d = (lizzieLet17_4QVal_Int_d[0] && (! lizzieLet17_4QVal_Int_emitted[0]));
  assign lizzieLet17_4QVal_Int_2_d = (lizzieLet17_4QVal_Int_d[0] && (! lizzieLet17_4QVal_Int_emitted[1]));
  assign lizzieLet17_4QVal_Int_3_d = (lizzieLet17_4QVal_Int_d[0] && (! lizzieLet17_4QVal_Int_emitted[2]));
  assign lizzieLet17_4QVal_Int_done = (lizzieLet17_4QVal_Int_emitted | ({lizzieLet17_4QVal_Int_3_d[0],
                                                                         lizzieLet17_4QVal_Int_2_d[0],
                                                                         lizzieLet17_4QVal_Int_1_d[0]} & {lizzieLet17_4QVal_Int_3_r,
                                                                                                          lizzieLet17_4QVal_Int_2_r,
                                                                                                          lizzieLet17_4QVal_Int_1_r}));
  assign lizzieLet17_4QVal_Int_r = (& lizzieLet17_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_emitted <= 3'd0;
    else
      lizzieLet17_4QVal_Int_emitted <= (lizzieLet17_4QVal_Int_r ? 3'd0 :
                                        lizzieLet17_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet17_4QVal_Int_1,Go) > (lizzieLet17_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet17_4QVal_Int_1_bufchan_d;
  logic lizzieLet17_4QVal_Int_1_bufchan_r;
  assign lizzieLet17_4QVal_Int_1_r = ((! lizzieLet17_4QVal_Int_1_bufchan_d[0]) || lizzieLet17_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QVal_Int_1_r)
        lizzieLet17_4QVal_Int_1_bufchan_d <= lizzieLet17_4QVal_Int_1_d;
  Go_t lizzieLet17_4QVal_Int_1_bufchan_buf;
  assign lizzieLet17_4QVal_Int_1_bufchan_r = (! lizzieLet17_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet17_4QVal_Int_1_argbuf_d = (lizzieLet17_4QVal_Int_1_bufchan_buf[0] ? lizzieLet17_4QVal_Int_1_bufchan_buf :
                                             lizzieLet17_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QVal_Int_1_argbuf_r && lizzieLet17_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet17_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QVal_Int_1_argbuf_r) && (! lizzieLet17_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet17_4QVal_Int_1_bufchan_buf <= lizzieLet17_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet17_4QVal_Int_1_argbuf,Go),
                                          (lizzieLet17_3QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (va8N_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet17_4QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet17_3QVal_Int_1_argbuf_d[0],
                                                                                             va8N_1_argbuf_d[0]}), lizzieLet17_4QVal_Int_1_argbuf_d, lizzieLet17_3QVal_Int_1_argbuf_d, va8N_1_argbuf_d);
  assign {lizzieLet17_4QVal_Int_1_argbuf_r,
          lizzieLet17_3QVal_Int_1_argbuf_r,
          va8N_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet17_4QVal_Int_2,Go) > (lizzieLet17_4QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet17_4QVal_Int_2_bufchan_d;
  logic lizzieLet17_4QVal_Int_2_bufchan_r;
  assign lizzieLet17_4QVal_Int_2_r = ((! lizzieLet17_4QVal_Int_2_bufchan_d[0]) || lizzieLet17_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_4QVal_Int_2_r)
        lizzieLet17_4QVal_Int_2_bufchan_d <= lizzieLet17_4QVal_Int_2_d;
  Go_t lizzieLet17_4QVal_Int_2_bufchan_buf;
  assign lizzieLet17_4QVal_Int_2_bufchan_r = (! lizzieLet17_4QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet17_4QVal_Int_2_argbuf_d = (lizzieLet17_4QVal_Int_2_bufchan_buf[0] ? lizzieLet17_4QVal_Int_2_bufchan_buf :
                                             lizzieLet17_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_4QVal_Int_2_argbuf_r && lizzieLet17_4QVal_Int_2_bufchan_buf[0]))
        lizzieLet17_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_4QVal_Int_2_argbuf_r) && (! lizzieLet17_4QVal_Int_2_bufchan_buf[0])))
        lizzieLet17_4QVal_Int_2_bufchan_buf <= lizzieLet17_4QVal_Int_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyBool,
      Dcon TupGo___MyDTBool_Bool___MyBool) : [(lizzieLet17_4QVal_Int_2_argbuf,Go),
                                              (lizzieLet17_5QVal_Int_1_argbuf,MyDTBool_Bool),
                                              (xa88_1_argbuf,MyBool)] > (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) */
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d = TupGo___MyDTBool_Bool___MyBool_dc((& {lizzieLet17_4QVal_Int_2_argbuf_d[0],
                                                                                                      lizzieLet17_5QVal_Int_1_argbuf_d[0],
                                                                                                      xa88_1_argbuf_d[0]}), lizzieLet17_4QVal_Int_2_argbuf_d, lizzieLet17_5QVal_Int_1_argbuf_d, xa88_1_argbuf_d);
  assign {lizzieLet17_4QVal_Int_2_argbuf_r,
          lizzieLet17_5QVal_Int_1_argbuf_r,
          xa88_1_argbuf_r} = {3 {(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTBool_Bool) : (lizzieLet17_5,QTree_Int) (isZa8K_goMux_mux,MyDTBool_Bool) > [(_51,MyDTBool_Bool),
                                                                                         (lizzieLet17_5QVal_Int,MyDTBool_Bool),
                                                                                         (lizzieLet17_5QNode_Int,MyDTBool_Bool),
                                                                                         (_50,MyDTBool_Bool)] */
  logic [3:0] isZa8K_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_5_d[0] && isZa8K_goMux_mux_d[0]))
      unique case (lizzieLet17_5_d[2:1])
        2'd0: isZa8K_goMux_mux_onehotd = 4'd1;
        2'd1: isZa8K_goMux_mux_onehotd = 4'd2;
        2'd2: isZa8K_goMux_mux_onehotd = 4'd4;
        2'd3: isZa8K_goMux_mux_onehotd = 4'd8;
        default: isZa8K_goMux_mux_onehotd = 4'd0;
      endcase
    else isZa8K_goMux_mux_onehotd = 4'd0;
  assign _51_d = isZa8K_goMux_mux_onehotd[0];
  assign lizzieLet17_5QVal_Int_d = isZa8K_goMux_mux_onehotd[1];
  assign lizzieLet17_5QNode_Int_d = isZa8K_goMux_mux_onehotd[2];
  assign _50_d = isZa8K_goMux_mux_onehotd[3];
  assign isZa8K_goMux_mux_r = (| (isZa8K_goMux_mux_onehotd & {_50_r,
                                                              lizzieLet17_5QNode_Int_r,
                                                              lizzieLet17_5QVal_Int_r,
                                                              _51_r}));
  assign lizzieLet17_5_r = isZa8K_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool) : (lizzieLet17_5QNode_Int,MyDTBool_Bool) > [(lizzieLet17_5QNode_Int_1,MyDTBool_Bool),
                                                                    (lizzieLet17_5QNode_Int_2,MyDTBool_Bool)] */
  logic [1:0] lizzieLet17_5QNode_Int_emitted;
  logic [1:0] lizzieLet17_5QNode_Int_done;
  assign lizzieLet17_5QNode_Int_1_d = (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[0]));
  assign lizzieLet17_5QNode_Int_2_d = (lizzieLet17_5QNode_Int_d[0] && (! lizzieLet17_5QNode_Int_emitted[1]));
  assign lizzieLet17_5QNode_Int_done = (lizzieLet17_5QNode_Int_emitted | ({lizzieLet17_5QNode_Int_2_d[0],
                                                                           lizzieLet17_5QNode_Int_1_d[0]} & {lizzieLet17_5QNode_Int_2_r,
                                                                                                             lizzieLet17_5QNode_Int_1_r}));
  assign lizzieLet17_5QNode_Int_r = (& lizzieLet17_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet17_5QNode_Int_emitted <= (lizzieLet17_5QNode_Int_r ? 2'd0 :
                                         lizzieLet17_5QNode_Int_done);
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet17_5QNode_Int_2,MyDTBool_Bool) > (lizzieLet17_5QNode_Int_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_2_bufchan_d;
  logic lizzieLet17_5QNode_Int_2_bufchan_r;
  assign lizzieLet17_5QNode_Int_2_r = ((! lizzieLet17_5QNode_Int_2_bufchan_d[0]) || lizzieLet17_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QNode_Int_2_r)
        lizzieLet17_5QNode_Int_2_bufchan_d <= lizzieLet17_5QNode_Int_2_d;
  MyDTBool_Bool_t lizzieLet17_5QNode_Int_2_bufchan_buf;
  assign lizzieLet17_5QNode_Int_2_bufchan_r = (! lizzieLet17_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet17_5QNode_Int_2_argbuf_d = (lizzieLet17_5QNode_Int_2_bufchan_buf[0] ? lizzieLet17_5QNode_Int_2_bufchan_buf :
                                              lizzieLet17_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QNode_Int_2_argbuf_r && lizzieLet17_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet17_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QNode_Int_2_argbuf_r) && (! lizzieLet17_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet17_5QNode_Int_2_bufchan_buf <= lizzieLet17_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet17_5QVal_Int,MyDTBool_Bool) > (lizzieLet17_5QVal_Int_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet17_5QVal_Int_bufchan_d;
  logic lizzieLet17_5QVal_Int_bufchan_r;
  assign lizzieLet17_5QVal_Int_r = ((! lizzieLet17_5QVal_Int_bufchan_d[0]) || lizzieLet17_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet17_5QVal_Int_r)
        lizzieLet17_5QVal_Int_bufchan_d <= lizzieLet17_5QVal_Int_d;
  MyDTBool_Bool_t lizzieLet17_5QVal_Int_bufchan_buf;
  assign lizzieLet17_5QVal_Int_bufchan_r = (! lizzieLet17_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet17_5QVal_Int_1_argbuf_d = (lizzieLet17_5QVal_Int_bufchan_buf[0] ? lizzieLet17_5QVal_Int_bufchan_buf :
                                             lizzieLet17_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet17_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet17_5QVal_Int_1_argbuf_r && lizzieLet17_5QVal_Int_bufchan_buf[0]))
        lizzieLet17_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet17_5QVal_Int_1_argbuf_r) && (! lizzieLet17_5QVal_Int_bufchan_buf[0])))
        lizzieLet17_5QVal_Int_bufchan_buf <= lizzieLet17_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTmain_map'_Int_Bool) : (lizzieLet17_6,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTmain_map'_Int_Bool) > [(lizzieLet17_6QNone_Int,Pointer_CTmain_map'_Int_Bool),
                                                                                                                       (lizzieLet17_6QVal_Int,Pointer_CTmain_map'_Int_Bool),
                                                                                                                       (lizzieLet17_6QNode_Int,Pointer_CTmain_map'_Int_Bool),
                                                                                                                       (lizzieLet17_6QError_Int,Pointer_CTmain_map'_Int_Bool)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet17_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet17_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet17_6QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet17_6QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                    sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet17_6QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                     sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet17_6QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet17_6QError_Int_r,
                                                              lizzieLet17_6QNode_Int_r,
                                                              lizzieLet17_6QVal_Int_r,
                                                              lizzieLet17_6QNone_Int_r}));
  assign lizzieLet17_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (lizzieLet17_6QError_Int,Pointer_CTmain_map'_Int_Bool) > (lizzieLet17_6QError_Int_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QError_Int_bufchan_d;
  logic lizzieLet17_6QError_Int_bufchan_r;
  assign lizzieLet17_6QError_Int_r = ((! lizzieLet17_6QError_Int_bufchan_d[0]) || lizzieLet17_6QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_6QError_Int_r)
        lizzieLet17_6QError_Int_bufchan_d <= lizzieLet17_6QError_Int_d;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QError_Int_bufchan_buf;
  assign lizzieLet17_6QError_Int_bufchan_r = (! lizzieLet17_6QError_Int_bufchan_buf[0]);
  assign lizzieLet17_6QError_Int_1_argbuf_d = (lizzieLet17_6QError_Int_bufchan_buf[0] ? lizzieLet17_6QError_Int_bufchan_buf :
                                               lizzieLet17_6QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_6QError_Int_1_argbuf_r && lizzieLet17_6QError_Int_bufchan_buf[0]))
        lizzieLet17_6QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_6QError_Int_1_argbuf_r) && (! lizzieLet17_6QError_Int_bufchan_buf[0])))
        lizzieLet17_6QError_Int_bufchan_buf <= lizzieLet17_6QError_Int_bufchan_d;
  
  /* dcon (Ty CTmain_map'_Int_Bool,
      Dcon Lcall_main_map'_Int_Bool3) : [(lizzieLet17_6QNode_Int,Pointer_CTmain_map'_Int_Bool),
                                         (lizzieLet17_5QNode_Int_1,MyDTBool_Bool),
                                         (lizzieLet17_3QNode_Int_1,MyDTInt_Bool),
                                         (q1a8O_destruct,Pointer_QTree_Int),
                                         (q2a8P_destruct,Pointer_QTree_Int),
                                         (q3a8Q_destruct,Pointer_QTree_Int)] > (lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3,CTmain_map'_Int_Bool) */
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_d  = \Lcall_main_map'_Int_Bool3_dc ((& {lizzieLet17_6QNode_Int_d[0],
                                                                                                                                                                         lizzieLet17_5QNode_Int_1_d[0],
                                                                                                                                                                         lizzieLet17_3QNode_Int_1_d[0],
                                                                                                                                                                         q1a8O_destruct_d[0],
                                                                                                                                                                         q2a8P_destruct_d[0],
                                                                                                                                                                         q3a8Q_destruct_d[0]}), lizzieLet17_6QNode_Int_d, lizzieLet17_5QNode_Int_1_d, lizzieLet17_3QNode_Int_1_d, q1a8O_destruct_d, q2a8P_destruct_d, q3a8Q_destruct_d);
  assign {lizzieLet17_6QNode_Int_r,
          lizzieLet17_5QNode_Int_1_r,
          lizzieLet17_3QNode_Int_1_r,
          q1a8O_destruct_r,
          q2a8P_destruct_r,
          q3a8Q_destruct_r} = {6 {(\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_r  && \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Bool) : (lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3,CTmain_map'_Int_Bool) > (lizzieLet21_1_argbuf,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d ;
  logic \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_r ;
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_r  = ((! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d [0]) || \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d  <= {67'd0,
                                                                                                                                             1'd0};
    else
      if (\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_r )
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d  <= \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_d ;
  \CTmain_map'_Int_Bool_t  \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf ;
  assign \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_r  = (! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf [0]);
  assign lizzieLet21_1_argbuf_d = (\lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf [0] ? \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf  :
                                   \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf  <= {67'd0,
                                                                                                                                               1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf [0]))
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf  <= {67'd0,
                                                                                                                                                 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf [0])))
        \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_buf  <= \lizzieLet17_6QNode_Int_1lizzieLet17_5QNode_Int_1lizzieLet17_3QNode_Int_1q1a8O_1q2a8P_1q3a8Q_1Lcall_main_map'_Int_Bool3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (lizzieLet17_6QNone_Int,Pointer_CTmain_map'_Int_Bool) > (lizzieLet17_6QNone_Int_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QNone_Int_bufchan_d;
  logic lizzieLet17_6QNone_Int_bufchan_r;
  assign lizzieLet17_6QNone_Int_r = ((! lizzieLet17_6QNone_Int_bufchan_d[0]) || lizzieLet17_6QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet17_6QNone_Int_r)
        lizzieLet17_6QNone_Int_bufchan_d <= lizzieLet17_6QNone_Int_d;
  \Pointer_CTmain_map'_Int_Bool_t  lizzieLet17_6QNone_Int_bufchan_buf;
  assign lizzieLet17_6QNone_Int_bufchan_r = (! lizzieLet17_6QNone_Int_bufchan_buf[0]);
  assign lizzieLet17_6QNone_Int_1_argbuf_d = (lizzieLet17_6QNone_Int_bufchan_buf[0] ? lizzieLet17_6QNone_Int_bufchan_buf :
                                              lizzieLet17_6QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet17_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet17_6QNone_Int_1_argbuf_r && lizzieLet17_6QNone_Int_bufchan_buf[0]))
        lizzieLet17_6QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet17_6QNone_Int_1_argbuf_r) && (! lizzieLet17_6QNone_Int_bufchan_buf[0])))
        lizzieLet17_6QNone_Int_bufchan_buf <= lizzieLet17_6QNone_Int_bufchan_d;
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int0) : (lizzieLet24_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) > [(es_2_1_destruct,Pointer_QTree_Int),
                                                                                     (es_3_2_destruct,Pointer_QTree_Int),
                                                                                     (es_4_3_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_6_destruct,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet24_1Lcall_$wmAdd_Int0_emitted;
  logic [3:0] lizzieLet24_1Lcall_$wmAdd_Int0_done;
  assign es_2_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int0_d[19:4],
                              (lizzieLet24_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int0_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int0_d[35:20],
                              (lizzieLet24_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int0_emitted[1]))};
  assign es_4_3_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int0_d[51:36],
                              (lizzieLet24_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int0_d[67:52],
                              (lizzieLet24_1Lcall_$wmAdd_Int0_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int0_emitted[3]))};
  assign lizzieLet24_1Lcall_$wmAdd_Int0_done = (lizzieLet24_1Lcall_$wmAdd_Int0_emitted | ({sc_0_6_destruct_d[0],
                                                                                           es_4_3_destruct_d[0],
                                                                                           es_3_2_destruct_d[0],
                                                                                           es_2_1_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                                    es_4_3_destruct_r,
                                                                                                                    es_3_2_destruct_r,
                                                                                                                    es_2_1_destruct_r}));
  assign lizzieLet24_1Lcall_$wmAdd_Int0_r = (& lizzieLet24_1Lcall_$wmAdd_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_$wmAdd_Int0_emitted <= 4'd0;
    else
      lizzieLet24_1Lcall_$wmAdd_Int0_emitted <= (lizzieLet24_1Lcall_$wmAdd_Int0_r ? 4'd0 :
                                                 lizzieLet24_1Lcall_$wmAdd_Int0_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int1) : (lizzieLet24_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) > [(es_3_1_destruct,Pointer_QTree_Int),
                                                                                     (es_4_2_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_5_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wslR_4_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8j_3_destruct,Pointer_QTree_Int),
                                                                                     (t1a8o_3_destruct,Pointer_QTree_Int)] */
  logic [5:0] lizzieLet24_1Lcall_$wmAdd_Int1_emitted;
  logic [5:0] lizzieLet24_1Lcall_$wmAdd_Int1_done;
  assign es_3_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int1_d[19:4],
                              (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[0]))};
  assign es_4_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int1_d[35:20],
                              (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int1_d[51:36],
                              (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[2]))};
  assign wslR_4_destruct_d = (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[3]));
  assign q1a8j_3_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int1_d[67:52],
                               (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[4]))};
  assign t1a8o_3_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int1_d[83:68],
                               (lizzieLet24_1Lcall_$wmAdd_Int1_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int1_emitted[5]))};
  assign lizzieLet24_1Lcall_$wmAdd_Int1_done = (lizzieLet24_1Lcall_$wmAdd_Int1_emitted | ({t1a8o_3_destruct_d[0],
                                                                                           q1a8j_3_destruct_d[0],
                                                                                           wslR_4_destruct_d[0],
                                                                                           sc_0_5_destruct_d[0],
                                                                                           es_4_2_destruct_d[0],
                                                                                           es_3_1_destruct_d[0]} & {t1a8o_3_destruct_r,
                                                                                                                    q1a8j_3_destruct_r,
                                                                                                                    wslR_4_destruct_r,
                                                                                                                    sc_0_5_destruct_r,
                                                                                                                    es_4_2_destruct_r,
                                                                                                                    es_3_1_destruct_r}));
  assign lizzieLet24_1Lcall_$wmAdd_Int1_r = (& lizzieLet24_1Lcall_$wmAdd_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_$wmAdd_Int1_emitted <= 6'd0;
    else
      lizzieLet24_1Lcall_$wmAdd_Int1_emitted <= (lizzieLet24_1Lcall_$wmAdd_Int1_r ? 6'd0 :
                                                 lizzieLet24_1Lcall_$wmAdd_Int1_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int2) : (lizzieLet24_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) > [(es_4_1_destruct,Pointer_QTree_Int),
                                                                                     (sc_0_4_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wslR_3_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8j_2_destruct,Pointer_QTree_Int),
                                                                                     (t1a8o_2_destruct,Pointer_QTree_Int),
                                                                                     (q2a8k_2_destruct,Pointer_QTree_Int),
                                                                                     (t2a8p_2_destruct,Pointer_QTree_Int)] */
  logic [6:0] lizzieLet24_1Lcall_$wmAdd_Int2_emitted;
  logic [6:0] lizzieLet24_1Lcall_$wmAdd_Int2_done;
  assign es_4_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[19:4],
                              (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[35:20],
                              (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[1]))};
  assign wslR_3_destruct_d = (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[2]));
  assign q1a8j_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[51:36],
                               (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[3]))};
  assign t1a8o_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[67:52],
                               (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[4]))};
  assign q2a8k_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[83:68],
                               (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[5]))};
  assign t2a8p_2_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int2_d[99:84],
                               (lizzieLet24_1Lcall_$wmAdd_Int2_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int2_emitted[6]))};
  assign lizzieLet24_1Lcall_$wmAdd_Int2_done = (lizzieLet24_1Lcall_$wmAdd_Int2_emitted | ({t2a8p_2_destruct_d[0],
                                                                                           q2a8k_2_destruct_d[0],
                                                                                           t1a8o_2_destruct_d[0],
                                                                                           q1a8j_2_destruct_d[0],
                                                                                           wslR_3_destruct_d[0],
                                                                                           sc_0_4_destruct_d[0],
                                                                                           es_4_1_destruct_d[0]} & {t2a8p_2_destruct_r,
                                                                                                                    q2a8k_2_destruct_r,
                                                                                                                    t1a8o_2_destruct_r,
                                                                                                                    q1a8j_2_destruct_r,
                                                                                                                    wslR_3_destruct_r,
                                                                                                                    sc_0_4_destruct_r,
                                                                                                                    es_4_1_destruct_r}));
  assign lizzieLet24_1Lcall_$wmAdd_Int2_r = (& lizzieLet24_1Lcall_$wmAdd_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_$wmAdd_Int2_emitted <= 7'd0;
    else
      lizzieLet24_1Lcall_$wmAdd_Int2_emitted <= (lizzieLet24_1Lcall_$wmAdd_Int2_r ? 7'd0 :
                                                 lizzieLet24_1Lcall_$wmAdd_Int2_done);
  
  /* destruct (Ty CT$wmAdd_Int,
          Dcon Lcall_$wmAdd_Int3) : (lizzieLet24_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) > [(sc_0_3_destruct,Pointer_CT$wmAdd_Int),
                                                                                     (wslR_2_destruct,MyDTInt_Int_Int),
                                                                                     (q1a8j_1_destruct,Pointer_QTree_Int),
                                                                                     (t1a8o_1_destruct,Pointer_QTree_Int),
                                                                                     (q2a8k_1_destruct,Pointer_QTree_Int),
                                                                                     (t2a8p_1_destruct,Pointer_QTree_Int),
                                                                                     (q3a8l_1_destruct,Pointer_QTree_Int),
                                                                                     (t3a8q_1_destruct,Pointer_QTree_Int)] */
  logic [7:0] lizzieLet24_1Lcall_$wmAdd_Int3_emitted;
  logic [7:0] lizzieLet24_1Lcall_$wmAdd_Int3_done;
  assign sc_0_3_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[19:4],
                              (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[0]))};
  assign wslR_2_destruct_d = (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[1]));
  assign q1a8j_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[35:20],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[2]))};
  assign t1a8o_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[51:36],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[3]))};
  assign q2a8k_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[67:52],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[4]))};
  assign t2a8p_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[83:68],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[5]))};
  assign q3a8l_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[99:84],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[6]))};
  assign t3a8q_1_destruct_d = {lizzieLet24_1Lcall_$wmAdd_Int3_d[115:100],
                               (lizzieLet24_1Lcall_$wmAdd_Int3_d[0] && (! lizzieLet24_1Lcall_$wmAdd_Int3_emitted[7]))};
  assign lizzieLet24_1Lcall_$wmAdd_Int3_done = (lizzieLet24_1Lcall_$wmAdd_Int3_emitted | ({t3a8q_1_destruct_d[0],
                                                                                           q3a8l_1_destruct_d[0],
                                                                                           t2a8p_1_destruct_d[0],
                                                                                           q2a8k_1_destruct_d[0],
                                                                                           t1a8o_1_destruct_d[0],
                                                                                           q1a8j_1_destruct_d[0],
                                                                                           wslR_2_destruct_d[0],
                                                                                           sc_0_3_destruct_d[0]} & {t3a8q_1_destruct_r,
                                                                                                                    q3a8l_1_destruct_r,
                                                                                                                    t2a8p_1_destruct_r,
                                                                                                                    q2a8k_1_destruct_r,
                                                                                                                    t1a8o_1_destruct_r,
                                                                                                                    q1a8j_1_destruct_r,
                                                                                                                    wslR_2_destruct_r,
                                                                                                                    sc_0_3_destruct_r}));
  assign lizzieLet24_1Lcall_$wmAdd_Int3_r = (& lizzieLet24_1Lcall_$wmAdd_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_$wmAdd_Int3_emitted <= 8'd0;
    else
      lizzieLet24_1Lcall_$wmAdd_Int3_emitted <= (lizzieLet24_1Lcall_$wmAdd_Int3_r ? 8'd0 :
                                                 lizzieLet24_1Lcall_$wmAdd_Int3_done);
  
  /* demux (Ty CT$wmAdd_Int,
       Ty CT$wmAdd_Int) : (lizzieLet24_2,CT$wmAdd_Int) (lizzieLet24_1,CT$wmAdd_Int) > [(_49,CT$wmAdd_Int),
                                                                                       (lizzieLet24_1Lcall_$wmAdd_Int3,CT$wmAdd_Int),
                                                                                       (lizzieLet24_1Lcall_$wmAdd_Int2,CT$wmAdd_Int),
                                                                                       (lizzieLet24_1Lcall_$wmAdd_Int1,CT$wmAdd_Int),
                                                                                       (lizzieLet24_1Lcall_$wmAdd_Int0,CT$wmAdd_Int)] */
  logic [4:0] lizzieLet24_1_onehotd;
  always_comb
    if ((lizzieLet24_2_d[0] && lizzieLet24_1_d[0]))
      unique case (lizzieLet24_2_d[3:1])
        3'd0: lizzieLet24_1_onehotd = 5'd1;
        3'd1: lizzieLet24_1_onehotd = 5'd2;
        3'd2: lizzieLet24_1_onehotd = 5'd4;
        3'd3: lizzieLet24_1_onehotd = 5'd8;
        3'd4: lizzieLet24_1_onehotd = 5'd16;
        default: lizzieLet24_1_onehotd = 5'd0;
      endcase
    else lizzieLet24_1_onehotd = 5'd0;
  assign _49_d = {lizzieLet24_1_d[115:1], lizzieLet24_1_onehotd[0]};
  assign lizzieLet24_1Lcall_$wmAdd_Int3_d = {lizzieLet24_1_d[115:1],
                                             lizzieLet24_1_onehotd[1]};
  assign lizzieLet24_1Lcall_$wmAdd_Int2_d = {lizzieLet24_1_d[115:1],
                                             lizzieLet24_1_onehotd[2]};
  assign lizzieLet24_1Lcall_$wmAdd_Int1_d = {lizzieLet24_1_d[115:1],
                                             lizzieLet24_1_onehotd[3]};
  assign lizzieLet24_1Lcall_$wmAdd_Int0_d = {lizzieLet24_1_d[115:1],
                                             lizzieLet24_1_onehotd[4]};
  assign lizzieLet24_1_r = (| (lizzieLet24_1_onehotd & {lizzieLet24_1Lcall_$wmAdd_Int0_r,
                                                        lizzieLet24_1Lcall_$wmAdd_Int1_r,
                                                        lizzieLet24_1Lcall_$wmAdd_Int2_r,
                                                        lizzieLet24_1Lcall_$wmAdd_Int3_r,
                                                        _49_r}));
  assign lizzieLet24_2_r = lizzieLet24_1_r;
  
  /* demux (Ty CT$wmAdd_Int,
       Ty Go) : (lizzieLet24_3,CT$wmAdd_Int) (go_15_goMux_data,Go) > [(_48,Go),
                                                                      (lizzieLet24_3Lcall_$wmAdd_Int3,Go),
                                                                      (lizzieLet24_3Lcall_$wmAdd_Int2,Go),
                                                                      (lizzieLet24_3Lcall_$wmAdd_Int1,Go),
                                                                      (lizzieLet24_3Lcall_$wmAdd_Int0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet24_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet24_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _48_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet24_3Lcall_$wmAdd_Int3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet24_3Lcall_$wmAdd_Int2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet24_3Lcall_$wmAdd_Int1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet24_3Lcall_$wmAdd_Int0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet24_3Lcall_$wmAdd_Int0_r,
                                                              lizzieLet24_3Lcall_$wmAdd_Int1_r,
                                                              lizzieLet24_3Lcall_$wmAdd_Int2_r,
                                                              lizzieLet24_3Lcall_$wmAdd_Int3_r,
                                                              _48_r}));
  assign lizzieLet24_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_$wmAdd_Int0,Go) > (lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_r;
  assign lizzieLet24_3Lcall_$wmAdd_Int0_r = ((! lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d[0]) || lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_$wmAdd_Int0_r)
        lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d <= lizzieLet24_3Lcall_$wmAdd_Int0_d;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf;
  assign lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_r = (! lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_d = (lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf[0] ? lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf :
                                                      lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_r && lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf[0]))
        lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_r) && (! lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf[0])))
        lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_buf <= lizzieLet24_3Lcall_$wmAdd_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_$wmAdd_Int1,Go) > (lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_r;
  assign lizzieLet24_3Lcall_$wmAdd_Int1_r = ((! lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d[0]) || lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_$wmAdd_Int1_r)
        lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d <= lizzieLet24_3Lcall_$wmAdd_Int1_d;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf;
  assign lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_r = (! lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_d = (lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf[0] ? lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf :
                                                      lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_r && lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf[0]))
        lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_$wmAdd_Int1_1_argbuf_r) && (! lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf[0])))
        lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_buf <= lizzieLet24_3Lcall_$wmAdd_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_$wmAdd_Int2,Go) > (lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_r;
  assign lizzieLet24_3Lcall_$wmAdd_Int2_r = ((! lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d[0]) || lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_$wmAdd_Int2_r)
        lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d <= lizzieLet24_3Lcall_$wmAdd_Int2_d;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf;
  assign lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_r = (! lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_d = (lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf[0] ? lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf :
                                                      lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_r && lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf[0]))
        lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_$wmAdd_Int2_1_argbuf_r) && (! lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf[0])))
        lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_buf <= lizzieLet24_3Lcall_$wmAdd_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_$wmAdd_Int3,Go) > (lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d;
  logic lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_r;
  assign lizzieLet24_3Lcall_$wmAdd_Int3_r = ((! lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d[0]) || lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_$wmAdd_Int3_r)
        lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d <= lizzieLet24_3Lcall_$wmAdd_Int3_d;
  Go_t lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf;
  assign lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_r = (! lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_d = (lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf[0] ? lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf :
                                                      lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_r && lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf[0]))
        lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_$wmAdd_Int3_1_argbuf_r) && (! lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf[0])))
        lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_buf <= lizzieLet24_3Lcall_$wmAdd_Int3_bufchan_d;
  
  /* demux (Ty CT$wmAdd_Int,
       Ty Pointer_QTree_Int) : (lizzieLet24_4,CT$wmAdd_Int) (srtarg_0_goMux_mux,Pointer_QTree_Int) > [(lizzieLet24_4L$wmAdd_Intsbos,Pointer_QTree_Int),
                                                                                                      (lizzieLet24_4Lcall_$wmAdd_Int3,Pointer_QTree_Int),
                                                                                                      (lizzieLet24_4Lcall_$wmAdd_Int2,Pointer_QTree_Int),
                                                                                                      (lizzieLet24_4Lcall_$wmAdd_Int1,Pointer_QTree_Int),
                                                                                                      (lizzieLet24_4Lcall_$wmAdd_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet24_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet24_4L$wmAdd_Intsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                           srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet24_4Lcall_$wmAdd_Int3_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet24_4Lcall_$wmAdd_Int2_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet24_4Lcall_$wmAdd_Int1_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet24_4Lcall_$wmAdd_Int0_d = {srtarg_0_goMux_mux_d[16:1],
                                             srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet24_4Lcall_$wmAdd_Int0_r,
                                                                  lizzieLet24_4Lcall_$wmAdd_Int1_r,
                                                                  lizzieLet24_4Lcall_$wmAdd_Int2_r,
                                                                  lizzieLet24_4Lcall_$wmAdd_Int3_r,
                                                                  lizzieLet24_4L$wmAdd_Intsbos_r}));
  assign lizzieLet24_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet24_4L$wmAdd_Intsbos,Pointer_QTree_Int) > [(lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                  (lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet24_4L$wmAdd_Intsbos_emitted;
  logic [1:0] lizzieLet24_4L$wmAdd_Intsbos_done;
  assign lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d = {lizzieLet24_4L$wmAdd_Intsbos_d[16:1],
                                                                (lizzieLet24_4L$wmAdd_Intsbos_d[0] && (! lizzieLet24_4L$wmAdd_Intsbos_emitted[0]))};
  assign lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d = {lizzieLet24_4L$wmAdd_Intsbos_d[16:1],
                                                                (lizzieLet24_4L$wmAdd_Intsbos_d[0] && (! lizzieLet24_4L$wmAdd_Intsbos_emitted[1]))};
  assign lizzieLet24_4L$wmAdd_Intsbos_done = (lizzieLet24_4L$wmAdd_Intsbos_emitted | ({lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                       lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                  lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet24_4L$wmAdd_Intsbos_r = (& lizzieLet24_4L$wmAdd_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet24_4L$wmAdd_Intsbos_emitted <= 2'd0;
    else
      lizzieLet24_4L$wmAdd_Intsbos_emitted <= (lizzieLet24_4L$wmAdd_Intsbos_r ? 2'd0 :
                                               lizzieLet24_4L$wmAdd_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_$wmAdd_Int_goConst,Go) */
  assign call_$wmAdd_Int_goConst_d = lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_1_r = call_$wmAdd_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > ($wmAdd_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                      1'd0};
    else
      if (lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wmAdd_Int_resbuf_d  = (lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                  lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                        1'd0};
    else
      if ((\$wmAdd_Int_resbuf_r  && lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                          1'd0};
      else if (((! \$wmAdd_Int_resbuf_r ) && (! lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet24_4L$wmAdd_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet24_4Lcall_$wmAdd_Int0,Pointer_QTree_Int),
                         (es_2_1_destruct,Pointer_QTree_Int),
                         (es_3_2_destruct,Pointer_QTree_Int),
                         (es_4_3_destruct,Pointer_QTree_Int)] > (lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int,QTree_Int) */
  assign lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_d = QNode_Int_dc((& {lizzieLet24_4Lcall_$wmAdd_Int0_d[0],
                                                                                                es_2_1_destruct_d[0],
                                                                                                es_3_2_destruct_d[0],
                                                                                                es_4_3_destruct_d[0]}), lizzieLet24_4Lcall_$wmAdd_Int0_d, es_2_1_destruct_d, es_3_2_destruct_d, es_4_3_destruct_d);
  assign {lizzieLet24_4Lcall_$wmAdd_Int0_r,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          es_4_3_destruct_r} = {4 {(lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_r && lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int,QTree_Int) > (lizzieLet28_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_r;
  assign lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_r = ((! lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d[0]) || lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d <= {66'd0,
                                                                                      1'd0};
    else
      if (lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_r)
        lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d <= lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_d;
  QTree_Int_t lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf;
  assign lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_r = (! lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf[0] ? lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf :
                                   lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf[0]))
        lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                          1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf[0])))
        lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_buf <= lizzieLet24_4Lcall_$wmAdd_Int0_1es_2_1_1es_3_2_1es_4_3_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int0) : [(lizzieLet24_4Lcall_$wmAdd_Int1,Pointer_QTree_Int),
                                 (es_3_1_destruct,Pointer_QTree_Int),
                                 (es_4_2_destruct,Pointer_QTree_Int),
                                 (sc_0_5_destruct,Pointer_CT$wmAdd_Int)] > (lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) */
  assign lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_d = Lcall_$wmAdd_Int0_dc((& {lizzieLet24_4Lcall_$wmAdd_Int1_d[0],
                                                                                                                es_3_1_destruct_d[0],
                                                                                                                es_4_2_destruct_d[0],
                                                                                                                sc_0_5_destruct_d[0]}), lizzieLet24_4Lcall_$wmAdd_Int1_d, es_3_1_destruct_d, es_4_2_destruct_d, sc_0_5_destruct_d);
  assign {lizzieLet24_4Lcall_$wmAdd_Int1_r,
          es_3_1_destruct_r,
          es_4_2_destruct_r,
          sc_0_5_destruct_r} = {4 {(lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_r && lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0,CT$wmAdd_Int) > (lizzieLet27_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r;
  assign lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_r = ((! lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d[0]) || lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_r)
        lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d <= lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_d;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf;
  assign lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_r = (! lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0] ? lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf :
                                   lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0]))
        lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf[0])))
        lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_buf <= lizzieLet24_4Lcall_$wmAdd_Int1_1es_3_1_1es_4_2_1sc_0_5_1Lcall_$wmAdd_Int0_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int1) : [(lizzieLet24_4Lcall_$wmAdd_Int2,Pointer_QTree_Int),
                                 (es_4_1_destruct,Pointer_QTree_Int),
                                 (sc_0_4_destruct,Pointer_CT$wmAdd_Int),
                                 (wslR_3_1,MyDTInt_Int_Int),
                                 (q1a8j_2_destruct,Pointer_QTree_Int),
                                 (t1a8o_2_destruct,Pointer_QTree_Int)] > (lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) */
  assign lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_d = Lcall_$wmAdd_Int1_dc((& {lizzieLet24_4Lcall_$wmAdd_Int2_d[0],
                                                                                                                                  es_4_1_destruct_d[0],
                                                                                                                                  sc_0_4_destruct_d[0],
                                                                                                                                  wslR_3_1_d[0],
                                                                                                                                  q1a8j_2_destruct_d[0],
                                                                                                                                  t1a8o_2_destruct_d[0]}), lizzieLet24_4Lcall_$wmAdd_Int2_d, es_4_1_destruct_d, sc_0_4_destruct_d, wslR_3_1_d, q1a8j_2_destruct_d, t1a8o_2_destruct_d);
  assign {lizzieLet24_4Lcall_$wmAdd_Int2_r,
          es_4_1_destruct_r,
          sc_0_4_destruct_r,
          wslR_3_1_r,
          q1a8j_2_destruct_r,
          t1a8o_2_destruct_r} = {6 {(lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_r && lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1,CT$wmAdd_Int) > (lizzieLet26_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_r;
  assign lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_r = ((! lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d[0]) || lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d <= {115'd0,
                                                                                                                1'd0};
    else
      if (lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_r)
        lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d <= lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_d;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf;
  assign lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_r = (! lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf[0] ? lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf :
                                   lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf <= {115'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf[0]))
        lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf <= {115'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf[0])))
        lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_buf <= lizzieLet24_4Lcall_$wmAdd_Int2_1es_4_1_1sc_0_4_1wslR_3_1q1a8j_2_1t1a8o_2_1Lcall_$wmAdd_Int1_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int2) : [(lizzieLet24_4Lcall_$wmAdd_Int3,Pointer_QTree_Int),
                                 (sc_0_3_destruct,Pointer_CT$wmAdd_Int),
                                 (wslR_2_1,MyDTInt_Int_Int),
                                 (q1a8j_1_destruct,Pointer_QTree_Int),
                                 (t1a8o_1_destruct,Pointer_QTree_Int),
                                 (q2a8k_1_destruct,Pointer_QTree_Int),
                                 (t2a8p_1_destruct,Pointer_QTree_Int)] > (lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) */
  assign lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_d = Lcall_$wmAdd_Int2_dc((& {lizzieLet24_4Lcall_$wmAdd_Int3_d[0],
                                                                                                                                            sc_0_3_destruct_d[0],
                                                                                                                                            wslR_2_1_d[0],
                                                                                                                                            q1a8j_1_destruct_d[0],
                                                                                                                                            t1a8o_1_destruct_d[0],
                                                                                                                                            q2a8k_1_destruct_d[0],
                                                                                                                                            t2a8p_1_destruct_d[0]}), lizzieLet24_4Lcall_$wmAdd_Int3_d, sc_0_3_destruct_d, wslR_2_1_d, q1a8j_1_destruct_d, t1a8o_1_destruct_d, q2a8k_1_destruct_d, t2a8p_1_destruct_d);
  assign {lizzieLet24_4Lcall_$wmAdd_Int3_r,
          sc_0_3_destruct_r,
          wslR_2_1_r,
          q1a8j_1_destruct_r,
          t1a8o_1_destruct_r,
          q2a8k_1_destruct_r,
          t2a8p_1_destruct_r} = {7 {(lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_r && lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2,CT$wmAdd_Int) > (lizzieLet25_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d;
  logic lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_r;
  assign lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_r = ((! lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d[0]) || lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d <= {115'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_r)
        lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d <= lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_d;
  CT$wmAdd_Int_t lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf;
  assign lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_r = (! lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf[0] ? lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf :
                                   lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf <= {115'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf[0]))
        lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf <= {115'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf[0])))
        lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_buf <= lizzieLet24_4Lcall_$wmAdd_Int3_1sc_0_3_1wslR_2_1q1a8j_1_1t1a8o_1_1q2a8k_1_1t2a8p_1_1Lcall_$wmAdd_Int2_bufchan_d;
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz0) : (lizzieLet29_1Lcall_$wnnz0,CT$wnnz) > [(wwslZ_3_destruct,Int#),
                                                                      (ww1XmJ_2_destruct,Int#),
                                                                      (ww2XmM_1_destruct,Int#),
                                                                      (sc_0_10_destruct,Pointer_CT$wnnz)] */
  logic [3:0] lizzieLet29_1Lcall_$wnnz0_emitted;
  logic [3:0] lizzieLet29_1Lcall_$wnnz0_done;
  assign wwslZ_3_destruct_d = {lizzieLet29_1Lcall_$wnnz0_d[35:4],
                               (lizzieLet29_1Lcall_$wnnz0_d[0] && (! lizzieLet29_1Lcall_$wnnz0_emitted[0]))};
  assign ww1XmJ_2_destruct_d = {lizzieLet29_1Lcall_$wnnz0_d[67:36],
                                (lizzieLet29_1Lcall_$wnnz0_d[0] && (! lizzieLet29_1Lcall_$wnnz0_emitted[1]))};
  assign ww2XmM_1_destruct_d = {lizzieLet29_1Lcall_$wnnz0_d[99:68],
                                (lizzieLet29_1Lcall_$wnnz0_d[0] && (! lizzieLet29_1Lcall_$wnnz0_emitted[2]))};
  assign sc_0_10_destruct_d = {lizzieLet29_1Lcall_$wnnz0_d[115:100],
                               (lizzieLet29_1Lcall_$wnnz0_d[0] && (! lizzieLet29_1Lcall_$wnnz0_emitted[3]))};
  assign lizzieLet29_1Lcall_$wnnz0_done = (lizzieLet29_1Lcall_$wnnz0_emitted | ({sc_0_10_destruct_d[0],
                                                                                 ww2XmM_1_destruct_d[0],
                                                                                 ww1XmJ_2_destruct_d[0],
                                                                                 wwslZ_3_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                           ww2XmM_1_destruct_r,
                                                                                                           ww1XmJ_2_destruct_r,
                                                                                                           wwslZ_3_destruct_r}));
  assign lizzieLet29_1Lcall_$wnnz0_r = (& lizzieLet29_1Lcall_$wnnz0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1Lcall_$wnnz0_emitted <= 4'd0;
    else
      lizzieLet29_1Lcall_$wnnz0_emitted <= (lizzieLet29_1Lcall_$wnnz0_r ? 4'd0 :
                                            lizzieLet29_1Lcall_$wnnz0_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz1) : (lizzieLet29_1Lcall_$wnnz1,CT$wnnz) > [(wwslZ_2_destruct,Int#),
                                                                      (ww1XmJ_1_destruct,Int#),
                                                                      (sc_0_9_destruct,Pointer_CT$wnnz),
                                                                      (q4a95_3_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet29_1Lcall_$wnnz1_emitted;
  logic [3:0] lizzieLet29_1Lcall_$wnnz1_done;
  assign wwslZ_2_destruct_d = {lizzieLet29_1Lcall_$wnnz1_d[35:4],
                               (lizzieLet29_1Lcall_$wnnz1_d[0] && (! lizzieLet29_1Lcall_$wnnz1_emitted[0]))};
  assign ww1XmJ_1_destruct_d = {lizzieLet29_1Lcall_$wnnz1_d[67:36],
                                (lizzieLet29_1Lcall_$wnnz1_d[0] && (! lizzieLet29_1Lcall_$wnnz1_emitted[1]))};
  assign sc_0_9_destruct_d = {lizzieLet29_1Lcall_$wnnz1_d[83:68],
                              (lizzieLet29_1Lcall_$wnnz1_d[0] && (! lizzieLet29_1Lcall_$wnnz1_emitted[2]))};
  assign q4a95_3_destruct_d = {lizzieLet29_1Lcall_$wnnz1_d[99:84],
                               (lizzieLet29_1Lcall_$wnnz1_d[0] && (! lizzieLet29_1Lcall_$wnnz1_emitted[3]))};
  assign lizzieLet29_1Lcall_$wnnz1_done = (lizzieLet29_1Lcall_$wnnz1_emitted | ({q4a95_3_destruct_d[0],
                                                                                 sc_0_9_destruct_d[0],
                                                                                 ww1XmJ_1_destruct_d[0],
                                                                                 wwslZ_2_destruct_d[0]} & {q4a95_3_destruct_r,
                                                                                                           sc_0_9_destruct_r,
                                                                                                           ww1XmJ_1_destruct_r,
                                                                                                           wwslZ_2_destruct_r}));
  assign lizzieLet29_1Lcall_$wnnz1_r = (& lizzieLet29_1Lcall_$wnnz1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1Lcall_$wnnz1_emitted <= 4'd0;
    else
      lizzieLet29_1Lcall_$wnnz1_emitted <= (lizzieLet29_1Lcall_$wnnz1_r ? 4'd0 :
                                            lizzieLet29_1Lcall_$wnnz1_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz2) : (lizzieLet29_1Lcall_$wnnz2,CT$wnnz) > [(wwslZ_1_destruct,Int#),
                                                                      (sc_0_8_destruct,Pointer_CT$wnnz),
                                                                      (q4a95_2_destruct,Pointer_QTree_Bool),
                                                                      (q3a94_2_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet29_1Lcall_$wnnz2_emitted;
  logic [3:0] lizzieLet29_1Lcall_$wnnz2_done;
  assign wwslZ_1_destruct_d = {lizzieLet29_1Lcall_$wnnz2_d[35:4],
                               (lizzieLet29_1Lcall_$wnnz2_d[0] && (! lizzieLet29_1Lcall_$wnnz2_emitted[0]))};
  assign sc_0_8_destruct_d = {lizzieLet29_1Lcall_$wnnz2_d[51:36],
                              (lizzieLet29_1Lcall_$wnnz2_d[0] && (! lizzieLet29_1Lcall_$wnnz2_emitted[1]))};
  assign q4a95_2_destruct_d = {lizzieLet29_1Lcall_$wnnz2_d[67:52],
                               (lizzieLet29_1Lcall_$wnnz2_d[0] && (! lizzieLet29_1Lcall_$wnnz2_emitted[2]))};
  assign q3a94_2_destruct_d = {lizzieLet29_1Lcall_$wnnz2_d[83:68],
                               (lizzieLet29_1Lcall_$wnnz2_d[0] && (! lizzieLet29_1Lcall_$wnnz2_emitted[3]))};
  assign lizzieLet29_1Lcall_$wnnz2_done = (lizzieLet29_1Lcall_$wnnz2_emitted | ({q3a94_2_destruct_d[0],
                                                                                 q4a95_2_destruct_d[0],
                                                                                 sc_0_8_destruct_d[0],
                                                                                 wwslZ_1_destruct_d[0]} & {q3a94_2_destruct_r,
                                                                                                           q4a95_2_destruct_r,
                                                                                                           sc_0_8_destruct_r,
                                                                                                           wwslZ_1_destruct_r}));
  assign lizzieLet29_1Lcall_$wnnz2_r = (& lizzieLet29_1Lcall_$wnnz2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1Lcall_$wnnz2_emitted <= 4'd0;
    else
      lizzieLet29_1Lcall_$wnnz2_emitted <= (lizzieLet29_1Lcall_$wnnz2_r ? 4'd0 :
                                            lizzieLet29_1Lcall_$wnnz2_done);
  
  /* destruct (Ty CT$wnnz,
          Dcon Lcall_$wnnz3) : (lizzieLet29_1Lcall_$wnnz3,CT$wnnz) > [(sc_0_7_destruct,Pointer_CT$wnnz),
                                                                      (q4a95_1_destruct,Pointer_QTree_Bool),
                                                                      (q3a94_1_destruct,Pointer_QTree_Bool),
                                                                      (q2a93_1_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet29_1Lcall_$wnnz3_emitted;
  logic [3:0] lizzieLet29_1Lcall_$wnnz3_done;
  assign sc_0_7_destruct_d = {lizzieLet29_1Lcall_$wnnz3_d[19:4],
                              (lizzieLet29_1Lcall_$wnnz3_d[0] && (! lizzieLet29_1Lcall_$wnnz3_emitted[0]))};
  assign q4a95_1_destruct_d = {lizzieLet29_1Lcall_$wnnz3_d[35:20],
                               (lizzieLet29_1Lcall_$wnnz3_d[0] && (! lizzieLet29_1Lcall_$wnnz3_emitted[1]))};
  assign q3a94_1_destruct_d = {lizzieLet29_1Lcall_$wnnz3_d[51:36],
                               (lizzieLet29_1Lcall_$wnnz3_d[0] && (! lizzieLet29_1Lcall_$wnnz3_emitted[2]))};
  assign q2a93_1_destruct_d = {lizzieLet29_1Lcall_$wnnz3_d[67:52],
                               (lizzieLet29_1Lcall_$wnnz3_d[0] && (! lizzieLet29_1Lcall_$wnnz3_emitted[3]))};
  assign lizzieLet29_1Lcall_$wnnz3_done = (lizzieLet29_1Lcall_$wnnz3_emitted | ({q2a93_1_destruct_d[0],
                                                                                 q3a94_1_destruct_d[0],
                                                                                 q4a95_1_destruct_d[0],
                                                                                 sc_0_7_destruct_d[0]} & {q2a93_1_destruct_r,
                                                                                                          q3a94_1_destruct_r,
                                                                                                          q4a95_1_destruct_r,
                                                                                                          sc_0_7_destruct_r}));
  assign lizzieLet29_1Lcall_$wnnz3_r = (& lizzieLet29_1Lcall_$wnnz3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_1Lcall_$wnnz3_emitted <= 4'd0;
    else
      lizzieLet29_1Lcall_$wnnz3_emitted <= (lizzieLet29_1Lcall_$wnnz3_r ? 4'd0 :
                                            lizzieLet29_1Lcall_$wnnz3_done);
  
  /* demux (Ty CT$wnnz,
       Ty CT$wnnz) : (lizzieLet29_2,CT$wnnz) (lizzieLet29_1,CT$wnnz) > [(_47,CT$wnnz),
                                                                        (lizzieLet29_1Lcall_$wnnz3,CT$wnnz),
                                                                        (lizzieLet29_1Lcall_$wnnz2,CT$wnnz),
                                                                        (lizzieLet29_1Lcall_$wnnz1,CT$wnnz),
                                                                        (lizzieLet29_1Lcall_$wnnz0,CT$wnnz)] */
  logic [4:0] lizzieLet29_1_onehotd;
  always_comb
    if ((lizzieLet29_2_d[0] && lizzieLet29_1_d[0]))
      unique case (lizzieLet29_2_d[3:1])
        3'd0: lizzieLet29_1_onehotd = 5'd1;
        3'd1: lizzieLet29_1_onehotd = 5'd2;
        3'd2: lizzieLet29_1_onehotd = 5'd4;
        3'd3: lizzieLet29_1_onehotd = 5'd8;
        3'd4: lizzieLet29_1_onehotd = 5'd16;
        default: lizzieLet29_1_onehotd = 5'd0;
      endcase
    else lizzieLet29_1_onehotd = 5'd0;
  assign _47_d = {lizzieLet29_1_d[115:1], lizzieLet29_1_onehotd[0]};
  assign lizzieLet29_1Lcall_$wnnz3_d = {lizzieLet29_1_d[115:1],
                                        lizzieLet29_1_onehotd[1]};
  assign lizzieLet29_1Lcall_$wnnz2_d = {lizzieLet29_1_d[115:1],
                                        lizzieLet29_1_onehotd[2]};
  assign lizzieLet29_1Lcall_$wnnz1_d = {lizzieLet29_1_d[115:1],
                                        lizzieLet29_1_onehotd[3]};
  assign lizzieLet29_1Lcall_$wnnz0_d = {lizzieLet29_1_d[115:1],
                                        lizzieLet29_1_onehotd[4]};
  assign lizzieLet29_1_r = (| (lizzieLet29_1_onehotd & {lizzieLet29_1Lcall_$wnnz0_r,
                                                        lizzieLet29_1Lcall_$wnnz1_r,
                                                        lizzieLet29_1Lcall_$wnnz2_r,
                                                        lizzieLet29_1Lcall_$wnnz3_r,
                                                        _47_r}));
  assign lizzieLet29_2_r = lizzieLet29_1_r;
  
  /* demux (Ty CT$wnnz,
       Ty Go) : (lizzieLet29_3,CT$wnnz) (go_16_goMux_data,Go) > [(_46,Go),
                                                                 (lizzieLet29_3Lcall_$wnnz3,Go),
                                                                 (lizzieLet29_3Lcall_$wnnz2,Go),
                                                                 (lizzieLet29_3Lcall_$wnnz1,Go),
                                                                 (lizzieLet29_3Lcall_$wnnz0,Go)] */
  logic [4:0] go_16_goMux_data_onehotd;
  always_comb
    if ((lizzieLet29_3_d[0] && go_16_goMux_data_d[0]))
      unique case (lizzieLet29_3_d[3:1])
        3'd0: go_16_goMux_data_onehotd = 5'd1;
        3'd1: go_16_goMux_data_onehotd = 5'd2;
        3'd2: go_16_goMux_data_onehotd = 5'd4;
        3'd3: go_16_goMux_data_onehotd = 5'd8;
        3'd4: go_16_goMux_data_onehotd = 5'd16;
        default: go_16_goMux_data_onehotd = 5'd0;
      endcase
    else go_16_goMux_data_onehotd = 5'd0;
  assign _46_d = go_16_goMux_data_onehotd[0];
  assign lizzieLet29_3Lcall_$wnnz3_d = go_16_goMux_data_onehotd[1];
  assign lizzieLet29_3Lcall_$wnnz2_d = go_16_goMux_data_onehotd[2];
  assign lizzieLet29_3Lcall_$wnnz1_d = go_16_goMux_data_onehotd[3];
  assign lizzieLet29_3Lcall_$wnnz0_d = go_16_goMux_data_onehotd[4];
  assign go_16_goMux_data_r = (| (go_16_goMux_data_onehotd & {lizzieLet29_3Lcall_$wnnz0_r,
                                                              lizzieLet29_3Lcall_$wnnz1_r,
                                                              lizzieLet29_3Lcall_$wnnz2_r,
                                                              lizzieLet29_3Lcall_$wnnz3_r,
                                                              _46_r}));
  assign lizzieLet29_3_r = go_16_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_$wnnz0,Go) > (lizzieLet29_3Lcall_$wnnz0_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_$wnnz0_bufchan_d;
  logic lizzieLet29_3Lcall_$wnnz0_bufchan_r;
  assign lizzieLet29_3Lcall_$wnnz0_r = ((! lizzieLet29_3Lcall_$wnnz0_bufchan_d[0]) || lizzieLet29_3Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz0_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_$wnnz0_r)
        lizzieLet29_3Lcall_$wnnz0_bufchan_d <= lizzieLet29_3Lcall_$wnnz0_d;
  Go_t lizzieLet29_3Lcall_$wnnz0_bufchan_buf;
  assign lizzieLet29_3Lcall_$wnnz0_bufchan_r = (! lizzieLet29_3Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_$wnnz0_1_argbuf_d = (lizzieLet29_3Lcall_$wnnz0_bufchan_buf[0] ? lizzieLet29_3Lcall_$wnnz0_bufchan_buf :
                                                 lizzieLet29_3Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_$wnnz0_1_argbuf_r && lizzieLet29_3Lcall_$wnnz0_bufchan_buf[0]))
        lizzieLet29_3Lcall_$wnnz0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_$wnnz0_1_argbuf_r) && (! lizzieLet29_3Lcall_$wnnz0_bufchan_buf[0])))
        lizzieLet29_3Lcall_$wnnz0_bufchan_buf <= lizzieLet29_3Lcall_$wnnz0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_$wnnz1,Go) > (lizzieLet29_3Lcall_$wnnz1_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_$wnnz1_bufchan_d;
  logic lizzieLet29_3Lcall_$wnnz1_bufchan_r;
  assign lizzieLet29_3Lcall_$wnnz1_r = ((! lizzieLet29_3Lcall_$wnnz1_bufchan_d[0]) || lizzieLet29_3Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz1_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_$wnnz1_r)
        lizzieLet29_3Lcall_$wnnz1_bufchan_d <= lizzieLet29_3Lcall_$wnnz1_d;
  Go_t lizzieLet29_3Lcall_$wnnz1_bufchan_buf;
  assign lizzieLet29_3Lcall_$wnnz1_bufchan_r = (! lizzieLet29_3Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_$wnnz1_1_argbuf_d = (lizzieLet29_3Lcall_$wnnz1_bufchan_buf[0] ? lizzieLet29_3Lcall_$wnnz1_bufchan_buf :
                                                 lizzieLet29_3Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_$wnnz1_1_argbuf_r && lizzieLet29_3Lcall_$wnnz1_bufchan_buf[0]))
        lizzieLet29_3Lcall_$wnnz1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_$wnnz1_1_argbuf_r) && (! lizzieLet29_3Lcall_$wnnz1_bufchan_buf[0])))
        lizzieLet29_3Lcall_$wnnz1_bufchan_buf <= lizzieLet29_3Lcall_$wnnz1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_$wnnz2,Go) > (lizzieLet29_3Lcall_$wnnz2_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_$wnnz2_bufchan_d;
  logic lizzieLet29_3Lcall_$wnnz2_bufchan_r;
  assign lizzieLet29_3Lcall_$wnnz2_r = ((! lizzieLet29_3Lcall_$wnnz2_bufchan_d[0]) || lizzieLet29_3Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz2_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_$wnnz2_r)
        lizzieLet29_3Lcall_$wnnz2_bufchan_d <= lizzieLet29_3Lcall_$wnnz2_d;
  Go_t lizzieLet29_3Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet29_3Lcall_$wnnz2_bufchan_r = (! lizzieLet29_3Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_$wnnz2_1_argbuf_d = (lizzieLet29_3Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet29_3Lcall_$wnnz2_bufchan_buf :
                                                 lizzieLet29_3Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_$wnnz2_1_argbuf_r && lizzieLet29_3Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet29_3Lcall_$wnnz2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_$wnnz2_1_argbuf_r) && (! lizzieLet29_3Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet29_3Lcall_$wnnz2_bufchan_buf <= lizzieLet29_3Lcall_$wnnz2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_$wnnz3,Go) > (lizzieLet29_3Lcall_$wnnz3_1_argbuf,Go) */
  Go_t lizzieLet29_3Lcall_$wnnz3_bufchan_d;
  logic lizzieLet29_3Lcall_$wnnz3_bufchan_r;
  assign lizzieLet29_3Lcall_$wnnz3_r = ((! lizzieLet29_3Lcall_$wnnz3_bufchan_d[0]) || lizzieLet29_3Lcall_$wnnz3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz3_bufchan_d <= 1'd0;
    else
      if (lizzieLet29_3Lcall_$wnnz3_r)
        lizzieLet29_3Lcall_$wnnz3_bufchan_d <= lizzieLet29_3Lcall_$wnnz3_d;
  Go_t lizzieLet29_3Lcall_$wnnz3_bufchan_buf;
  assign lizzieLet29_3Lcall_$wnnz3_bufchan_r = (! lizzieLet29_3Lcall_$wnnz3_bufchan_buf[0]);
  assign lizzieLet29_3Lcall_$wnnz3_1_argbuf_d = (lizzieLet29_3Lcall_$wnnz3_bufchan_buf[0] ? lizzieLet29_3Lcall_$wnnz3_bufchan_buf :
                                                 lizzieLet29_3Lcall_$wnnz3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet29_3Lcall_$wnnz3_1_argbuf_r && lizzieLet29_3Lcall_$wnnz3_bufchan_buf[0]))
        lizzieLet29_3Lcall_$wnnz3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet29_3Lcall_$wnnz3_1_argbuf_r) && (! lizzieLet29_3Lcall_$wnnz3_bufchan_buf[0])))
        lizzieLet29_3Lcall_$wnnz3_bufchan_buf <= lizzieLet29_3Lcall_$wnnz3_bufchan_d;
  
  /* demux (Ty CT$wnnz,
       Ty Int#) : (lizzieLet29_4,CT$wnnz) (srtarg_0_1_goMux_mux,Int#) > [(lizzieLet29_4L$wnnzsbos,Int#),
                                                                         (lizzieLet29_4Lcall_$wnnz3,Int#),
                                                                         (lizzieLet29_4Lcall_$wnnz2,Int#),
                                                                         (lizzieLet29_4Lcall_$wnnz1,Int#),
                                                                         (lizzieLet29_4Lcall_$wnnz0,Int#)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet29_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet29_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet29_4L$wnnzsbos_d = {srtarg_0_1_goMux_mux_d[32:1],
                                      srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet29_4Lcall_$wnnz3_d = {srtarg_0_1_goMux_mux_d[32:1],
                                        srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet29_4Lcall_$wnnz2_d = {srtarg_0_1_goMux_mux_d[32:1],
                                        srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet29_4Lcall_$wnnz1_d = {srtarg_0_1_goMux_mux_d[32:1],
                                        srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet29_4Lcall_$wnnz0_d = {srtarg_0_1_goMux_mux_d[32:1],
                                        srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet29_4Lcall_$wnnz0_r,
                                                                      lizzieLet29_4Lcall_$wnnz1_r,
                                                                      lizzieLet29_4Lcall_$wnnz2_r,
                                                                      lizzieLet29_4Lcall_$wnnz3_r,
                                                                      lizzieLet29_4L$wnnzsbos_r}));
  assign lizzieLet29_4_r = srtarg_0_1_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet29_4L$wnnzsbos,Int#) > [(lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1,Int#),
                                                   (lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet29_4L$wnnzsbos_emitted;
  logic [1:0] lizzieLet29_4L$wnnzsbos_done;
  assign lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_d = {lizzieLet29_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet29_4L$wnnzsbos_d[0] && (! lizzieLet29_4L$wnnzsbos_emitted[0]))};
  assign lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_d = {lizzieLet29_4L$wnnzsbos_d[32:1],
                                                           (lizzieLet29_4L$wnnzsbos_d[0] && (! lizzieLet29_4L$wnnzsbos_emitted[1]))};
  assign lizzieLet29_4L$wnnzsbos_done = (lizzieLet29_4L$wnnzsbos_emitted | ({lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_d[0],
                                                                             lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_r,
                                                                                                                                   lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet29_4L$wnnzsbos_r = (& lizzieLet29_4L$wnnzsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet29_4L$wnnzsbos_emitted <= 2'd0;
    else
      lizzieLet29_4L$wnnzsbos_emitted <= (lizzieLet29_4L$wnnzsbos_r ? 2'd0 :
                                          lizzieLet29_4L$wnnzsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_goConst,Go) */
  assign call_$wnnz_goConst_d = lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_1_r = call_$wnnz_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2,Int#) > ($wnnz_resbuf,Int#) */
  \Int#_t  lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_r = ((! lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                 1'd0};
    else
      if (lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_r)
        lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_resbuf_d  = (lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf :
                             lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                   1'd0};
    else
      if ((\$wnnz_resbuf_r  && lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                     1'd0};
      else if (((! \$wnnz_resbuf_r ) && (! lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet29_4L$wnnzsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz,
      Dcon Lcall_$wnnz2) : [(lizzieLet29_4Lcall_$wnnz3,Int#),
                            (sc_0_7_destruct,Pointer_CT$wnnz),
                            (q4a95_1_destruct,Pointer_QTree_Bool),
                            (q3a94_1_destruct,Pointer_QTree_Bool)] > (lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2,CT$wnnz) */
  assign lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_d = Lcall_$wnnz2_dc((& {lizzieLet29_4Lcall_$wnnz3_d[0],
                                                                                                   sc_0_7_destruct_d[0],
                                                                                                   q4a95_1_destruct_d[0],
                                                                                                   q3a94_1_destruct_d[0]}), lizzieLet29_4Lcall_$wnnz3_d, sc_0_7_destruct_d, q4a95_1_destruct_d, q3a94_1_destruct_d);
  assign {lizzieLet29_4Lcall_$wnnz3_r,
          sc_0_7_destruct_r,
          q4a95_1_destruct_r,
          q3a94_1_destruct_r} = {4 {(lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_r && lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_d[0])}};
  
  /* buf (Ty CT$wnnz) : (lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2,CT$wnnz) > (lizzieLet30_1_argbuf,CT$wnnz) */
  CT$wnnz_t lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d;
  logic lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_r;
  assign lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_r = ((! lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d[0]) || lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_r)
        lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d <= lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_d;
  CT$wnnz_t lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf;
  assign lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_r = (! lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf[0] ? lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf :
                                   lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf[0]))
        lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf[0])))
        lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_buf <= lizzieLet29_4Lcall_$wnnz3_1sc_0_7_1q4a95_1_1q3a94_1_1Lcall_$wnnz2_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet2_1wild1XF_1_Eq,Bool) > (lizzieLet3_1_argbuf,Bool) */
  Bool_t lizzieLet2_1wild1XF_1_Eq_bufchan_d;
  logic lizzieLet2_1wild1XF_1_Eq_bufchan_r;
  assign lizzieLet2_1wild1XF_1_Eq_r = ((! lizzieLet2_1wild1XF_1_Eq_bufchan_d[0]) || lizzieLet2_1wild1XF_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_1wild1XF_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet2_1wild1XF_1_Eq_r)
        lizzieLet2_1wild1XF_1_Eq_bufchan_d <= lizzieLet2_1wild1XF_1_Eq_d;
  Bool_t lizzieLet2_1wild1XF_1_Eq_bufchan_buf;
  assign lizzieLet2_1wild1XF_1_Eq_bufchan_r = (! lizzieLet2_1wild1XF_1_Eq_bufchan_buf[0]);
  assign lizzieLet3_1_argbuf_d = (lizzieLet2_1wild1XF_1_Eq_bufchan_buf[0] ? lizzieLet2_1wild1XF_1_Eq_bufchan_buf :
                                  lizzieLet2_1wild1XF_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_1wild1XF_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet3_1_argbuf_r && lizzieLet2_1wild1XF_1_Eq_bufchan_buf[0]))
        lizzieLet2_1wild1XF_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet3_1_argbuf_r) && (! lizzieLet2_1wild1XF_1_Eq_bufchan_buf[0])))
        lizzieLet2_1wild1XF_1_Eq_bufchan_buf <= lizzieLet2_1wild1XF_1_Eq_bufchan_d;
  
  /* destruct (Ty CTmain_map'_Int_Bool,
          Dcon Lcall_main_map'_Int_Bool0) : (lizzieLet33_1Lcall_main_map'_Int_Bool0,CTmain_map'_Int_Bool) > [(es_2_2_destruct,Pointer_QTree_Bool),
                                                                                                             (es_3_4_destruct,Pointer_QTree_Bool),
                                                                                                             (es_4_7_destruct,Pointer_QTree_Bool),
                                                                                                             (sc_0_14_destruct,Pointer_CTmain_map'_Int_Bool)] */
  logic [3:0] \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted ;
  logic [3:0] \lizzieLet33_1Lcall_main_map'_Int_Bool0_done ;
  assign es_2_2_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [19:4],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted [0]))};
  assign es_3_4_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [35:20],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted [1]))};
  assign es_4_7_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [51:36],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted [2]))};
  assign sc_0_14_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [67:52],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool0_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted [3]))};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool0_done  = (\lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted  | ({sc_0_14_destruct_d[0],
                                                                                                               es_4_7_destruct_d[0],
                                                                                                               es_3_4_destruct_d[0],
                                                                                                               es_2_2_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                                        es_4_7_destruct_r,
                                                                                                                                        es_3_4_destruct_r,
                                                                                                                                        es_2_2_destruct_r}));
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool0_r  = (& \lizzieLet33_1Lcall_main_map'_Int_Bool0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted  <= 4'd0;
    else
      \lizzieLet33_1Lcall_main_map'_Int_Bool0_emitted  <= (\lizzieLet33_1Lcall_main_map'_Int_Bool0_r  ? 4'd0 :
                                                           \lizzieLet33_1Lcall_main_map'_Int_Bool0_done );
  
  /* destruct (Ty CTmain_map'_Int_Bool,
          Dcon Lcall_main_map'_Int_Bool1) : (lizzieLet33_1Lcall_main_map'_Int_Bool1,CTmain_map'_Int_Bool) > [(es_3_3_destruct,Pointer_QTree_Bool),
                                                                                                             (es_4_6_destruct,Pointer_QTree_Bool),
                                                                                                             (sc_0_13_destruct,Pointer_CTmain_map'_Int_Bool),
                                                                                                             (isZa8K_4_destruct,MyDTBool_Bool),
                                                                                                             (ga8L_4_destruct,MyDTInt_Bool),
                                                                                                             (q1a8O_3_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted ;
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool1_done ;
  assign es_3_3_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [19:4],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [0]))};
  assign es_4_6_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [35:20],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [1]))};
  assign sc_0_13_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [51:36],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [2]))};
  assign isZa8K_4_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [3]));
  assign ga8L_4_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [4]));
  assign q1a8O_3_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [67:52],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool1_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted [5]))};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool1_done  = (\lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted  | ({q1a8O_3_destruct_d[0],
                                                                                                               ga8L_4_destruct_d[0],
                                                                                                               isZa8K_4_destruct_d[0],
                                                                                                               sc_0_13_destruct_d[0],
                                                                                                               es_4_6_destruct_d[0],
                                                                                                               es_3_3_destruct_d[0]} & {q1a8O_3_destruct_r,
                                                                                                                                        ga8L_4_destruct_r,
                                                                                                                                        isZa8K_4_destruct_r,
                                                                                                                                        sc_0_13_destruct_r,
                                                                                                                                        es_4_6_destruct_r,
                                                                                                                                        es_3_3_destruct_r}));
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool1_r  = (& \lizzieLet33_1Lcall_main_map'_Int_Bool1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted  <= 6'd0;
    else
      \lizzieLet33_1Lcall_main_map'_Int_Bool1_emitted  <= (\lizzieLet33_1Lcall_main_map'_Int_Bool1_r  ? 6'd0 :
                                                           \lizzieLet33_1Lcall_main_map'_Int_Bool1_done );
  
  /* destruct (Ty CTmain_map'_Int_Bool,
          Dcon Lcall_main_map'_Int_Bool2) : (lizzieLet33_1Lcall_main_map'_Int_Bool2,CTmain_map'_Int_Bool) > [(es_4_5_destruct,Pointer_QTree_Bool),
                                                                                                             (sc_0_12_destruct,Pointer_CTmain_map'_Int_Bool),
                                                                                                             (isZa8K_3_destruct,MyDTBool_Bool),
                                                                                                             (ga8L_3_destruct,MyDTInt_Bool),
                                                                                                             (q1a8O_2_destruct,Pointer_QTree_Int),
                                                                                                             (q2a8P_2_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted ;
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool2_done ;
  assign es_4_5_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [19:4],
                              (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [0]))};
  assign sc_0_12_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [35:20],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [1]))};
  assign isZa8K_3_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [2]));
  assign ga8L_3_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [3]));
  assign q1a8O_2_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [51:36],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [4]))};
  assign q2a8P_2_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [67:52],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool2_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted [5]))};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool2_done  = (\lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted  | ({q2a8P_2_destruct_d[0],
                                                                                                               q1a8O_2_destruct_d[0],
                                                                                                               ga8L_3_destruct_d[0],
                                                                                                               isZa8K_3_destruct_d[0],
                                                                                                               sc_0_12_destruct_d[0],
                                                                                                               es_4_5_destruct_d[0]} & {q2a8P_2_destruct_r,
                                                                                                                                        q1a8O_2_destruct_r,
                                                                                                                                        ga8L_3_destruct_r,
                                                                                                                                        isZa8K_3_destruct_r,
                                                                                                                                        sc_0_12_destruct_r,
                                                                                                                                        es_4_5_destruct_r}));
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool2_r  = (& \lizzieLet33_1Lcall_main_map'_Int_Bool2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted  <= 6'd0;
    else
      \lizzieLet33_1Lcall_main_map'_Int_Bool2_emitted  <= (\lizzieLet33_1Lcall_main_map'_Int_Bool2_r  ? 6'd0 :
                                                           \lizzieLet33_1Lcall_main_map'_Int_Bool2_done );
  
  /* destruct (Ty CTmain_map'_Int_Bool,
          Dcon Lcall_main_map'_Int_Bool3) : (lizzieLet33_1Lcall_main_map'_Int_Bool3,CTmain_map'_Int_Bool) > [(sc_0_11_destruct,Pointer_CTmain_map'_Int_Bool),
                                                                                                             (isZa8K_2_destruct,MyDTBool_Bool),
                                                                                                             (ga8L_2_destruct,MyDTInt_Bool),
                                                                                                             (q1a8O_1_destruct,Pointer_QTree_Int),
                                                                                                             (q2a8P_1_destruct,Pointer_QTree_Int),
                                                                                                             (q3a8Q_1_destruct,Pointer_QTree_Int)] */
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted ;
  logic [5:0] \lizzieLet33_1Lcall_main_map'_Int_Bool3_done ;
  assign sc_0_11_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [19:4],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [0]))};
  assign isZa8K_2_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [1]));
  assign ga8L_2_destruct_d = (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [2]));
  assign q1a8O_1_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [35:20],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [3]))};
  assign q2a8P_1_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [51:36],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [4]))};
  assign q3a8Q_1_destruct_d = {\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [67:52],
                               (\lizzieLet33_1Lcall_main_map'_Int_Bool3_d [0] && (! \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted [5]))};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool3_done  = (\lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted  | ({q3a8Q_1_destruct_d[0],
                                                                                                               q2a8P_1_destruct_d[0],
                                                                                                               q1a8O_1_destruct_d[0],
                                                                                                               ga8L_2_destruct_d[0],
                                                                                                               isZa8K_2_destruct_d[0],
                                                                                                               sc_0_11_destruct_d[0]} & {q3a8Q_1_destruct_r,
                                                                                                                                         q2a8P_1_destruct_r,
                                                                                                                                         q1a8O_1_destruct_r,
                                                                                                                                         ga8L_2_destruct_r,
                                                                                                                                         isZa8K_2_destruct_r,
                                                                                                                                         sc_0_11_destruct_r}));
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool3_r  = (& \lizzieLet33_1Lcall_main_map'_Int_Bool3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted  <= 6'd0;
    else
      \lizzieLet33_1Lcall_main_map'_Int_Bool3_emitted  <= (\lizzieLet33_1Lcall_main_map'_Int_Bool3_r  ? 6'd0 :
                                                           \lizzieLet33_1Lcall_main_map'_Int_Bool3_done );
  
  /* demux (Ty CTmain_map'_Int_Bool,
       Ty CTmain_map'_Int_Bool) : (lizzieLet33_2,CTmain_map'_Int_Bool) (lizzieLet33_1,CTmain_map'_Int_Bool) > [(_45,CTmain_map'_Int_Bool),
                                                                                                               (lizzieLet33_1Lcall_main_map'_Int_Bool3,CTmain_map'_Int_Bool),
                                                                                                               (lizzieLet33_1Lcall_main_map'_Int_Bool2,CTmain_map'_Int_Bool),
                                                                                                               (lizzieLet33_1Lcall_main_map'_Int_Bool1,CTmain_map'_Int_Bool),
                                                                                                               (lizzieLet33_1Lcall_main_map'_Int_Bool0,CTmain_map'_Int_Bool)] */
  logic [4:0] lizzieLet33_1_onehotd;
  always_comb
    if ((lizzieLet33_2_d[0] && lizzieLet33_1_d[0]))
      unique case (lizzieLet33_2_d[3:1])
        3'd0: lizzieLet33_1_onehotd = 5'd1;
        3'd1: lizzieLet33_1_onehotd = 5'd2;
        3'd2: lizzieLet33_1_onehotd = 5'd4;
        3'd3: lizzieLet33_1_onehotd = 5'd8;
        3'd4: lizzieLet33_1_onehotd = 5'd16;
        default: lizzieLet33_1_onehotd = 5'd0;
      endcase
    else lizzieLet33_1_onehotd = 5'd0;
  assign _45_d = {lizzieLet33_1_d[67:1], lizzieLet33_1_onehotd[0]};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool3_d  = {lizzieLet33_1_d[67:1],
                                                       lizzieLet33_1_onehotd[1]};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool2_d  = {lizzieLet33_1_d[67:1],
                                                       lizzieLet33_1_onehotd[2]};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool1_d  = {lizzieLet33_1_d[67:1],
                                                       lizzieLet33_1_onehotd[3]};
  assign \lizzieLet33_1Lcall_main_map'_Int_Bool0_d  = {lizzieLet33_1_d[67:1],
                                                       lizzieLet33_1_onehotd[4]};
  assign lizzieLet33_1_r = (| (lizzieLet33_1_onehotd & {\lizzieLet33_1Lcall_main_map'_Int_Bool0_r ,
                                                        \lizzieLet33_1Lcall_main_map'_Int_Bool1_r ,
                                                        \lizzieLet33_1Lcall_main_map'_Int_Bool2_r ,
                                                        \lizzieLet33_1Lcall_main_map'_Int_Bool3_r ,
                                                        _45_r}));
  assign lizzieLet33_2_r = lizzieLet33_1_r;
  
  /* demux (Ty CTmain_map'_Int_Bool,
       Ty Go) : (lizzieLet33_3,CTmain_map'_Int_Bool) (go_17_goMux_data,Go) > [(_44,Go),
                                                                              (lizzieLet33_3Lcall_main_map'_Int_Bool3,Go),
                                                                              (lizzieLet33_3Lcall_main_map'_Int_Bool2,Go),
                                                                              (lizzieLet33_3Lcall_main_map'_Int_Bool1,Go),
                                                                              (lizzieLet33_3Lcall_main_map'_Int_Bool0,Go)] */
  logic [4:0] go_17_goMux_data_onehotd;
  always_comb
    if ((lizzieLet33_3_d[0] && go_17_goMux_data_d[0]))
      unique case (lizzieLet33_3_d[3:1])
        3'd0: go_17_goMux_data_onehotd = 5'd1;
        3'd1: go_17_goMux_data_onehotd = 5'd2;
        3'd2: go_17_goMux_data_onehotd = 5'd4;
        3'd3: go_17_goMux_data_onehotd = 5'd8;
        3'd4: go_17_goMux_data_onehotd = 5'd16;
        default: go_17_goMux_data_onehotd = 5'd0;
      endcase
    else go_17_goMux_data_onehotd = 5'd0;
  assign _44_d = go_17_goMux_data_onehotd[0];
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool3_d  = go_17_goMux_data_onehotd[1];
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool2_d  = go_17_goMux_data_onehotd[2];
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool1_d  = go_17_goMux_data_onehotd[3];
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool0_d  = go_17_goMux_data_onehotd[4];
  assign go_17_goMux_data_r = (| (go_17_goMux_data_onehotd & {\lizzieLet33_3Lcall_main_map'_Int_Bool0_r ,
                                                              \lizzieLet33_3Lcall_main_map'_Int_Bool1_r ,
                                                              \lizzieLet33_3Lcall_main_map'_Int_Bool2_r ,
                                                              \lizzieLet33_3Lcall_main_map'_Int_Bool3_r ,
                                                              _44_r}));
  assign lizzieLet33_3_r = go_17_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet33_3Lcall_main_map'_Int_Bool0,Go) > (lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf,Go) */
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_r ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool0_r  = ((! \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d [0]) || \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet33_3Lcall_main_map'_Int_Bool0_r )
        \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d  <= \lizzieLet33_3Lcall_main_map'_Int_Bool0_d ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_r  = (! \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf [0]);
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_d  = (\lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf [0] ? \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf  :
                                                                \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_r  && \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf [0]))
        \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet33_3Lcall_main_map'_Int_Bool0_1_argbuf_r ) && (! \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf [0])))
        \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_buf  <= \lizzieLet33_3Lcall_main_map'_Int_Bool0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet33_3Lcall_main_map'_Int_Bool1,Go) > (lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf,Go) */
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_r ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool1_r  = ((! \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d [0]) || \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet33_3Lcall_main_map'_Int_Bool1_r )
        \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d  <= \lizzieLet33_3Lcall_main_map'_Int_Bool1_d ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_r  = (! \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf [0]);
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_d  = (\lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf [0] ? \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf  :
                                                                \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_r  && \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf [0]))
        \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet33_3Lcall_main_map'_Int_Bool1_1_argbuf_r ) && (! \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf [0])))
        \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_buf  <= \lizzieLet33_3Lcall_main_map'_Int_Bool1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet33_3Lcall_main_map'_Int_Bool2,Go) > (lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf,Go) */
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_r ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool2_r  = ((! \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d [0]) || \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet33_3Lcall_main_map'_Int_Bool2_r )
        \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d  <= \lizzieLet33_3Lcall_main_map'_Int_Bool2_d ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_r  = (! \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf [0]);
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_d  = (\lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf [0] ? \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf  :
                                                                \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_r  && \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf [0]))
        \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet33_3Lcall_main_map'_Int_Bool2_1_argbuf_r ) && (! \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf [0])))
        \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_buf  <= \lizzieLet33_3Lcall_main_map'_Int_Bool2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet33_3Lcall_main_map'_Int_Bool3,Go) > (lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf,Go) */
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d ;
  logic \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_r ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool3_r  = ((! \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d [0]) || \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet33_3Lcall_main_map'_Int_Bool3_r )
        \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d  <= \lizzieLet33_3Lcall_main_map'_Int_Bool3_d ;
  Go_t \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf ;
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_r  = (! \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf [0]);
  assign \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_d  = (\lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf [0] ? \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf  :
                                                                \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_r  && \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf [0]))
        \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet33_3Lcall_main_map'_Int_Bool3_1_argbuf_r ) && (! \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf [0])))
        \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_buf  <= \lizzieLet33_3Lcall_main_map'_Int_Bool3_bufchan_d ;
  
  /* demux (Ty CTmain_map'_Int_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet33_4,CTmain_map'_Int_Bool) (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet33_4Lmain_map'_Int_Boolsbos,Pointer_QTree_Bool),
                                                                                                                  (lizzieLet33_4Lcall_main_map'_Int_Bool3,Pointer_QTree_Bool),
                                                                                                                  (lizzieLet33_4Lcall_main_map'_Int_Bool2,Pointer_QTree_Bool),
                                                                                                                  (lizzieLet33_4Lcall_main_map'_Int_Bool1,Pointer_QTree_Bool),
                                                                                                                  (lizzieLet33_4Lcall_main_map'_Int_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet33_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet33_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                     srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                       srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                       srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                       srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                       srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet33_4Lcall_main_map'_Int_Bool0_r ,
                                                                      \lizzieLet33_4Lcall_main_map'_Int_Bool1_r ,
                                                                      \lizzieLet33_4Lcall_main_map'_Int_Bool2_r ,
                                                                      \lizzieLet33_4Lcall_main_map'_Int_Bool3_r ,
                                                                      \lizzieLet33_4Lmain_map'_Int_Boolsbos_r }));
  assign lizzieLet33_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet33_4Lcall_main_map'_Int_Bool0,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_4_destruct,Pointer_QTree_Bool),
                          (es_4_7_destruct,Pointer_QTree_Bool)] > (lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet33_4Lcall_main_map'_Int_Bool0_d [0],
                                                                                                            es_2_2_destruct_d[0],
                                                                                                            es_3_4_destruct_d[0],
                                                                                                            es_4_7_destruct_d[0]}), \lizzieLet33_4Lcall_main_map'_Int_Bool0_d , es_2_2_destruct_d, es_3_4_destruct_d, es_4_7_destruct_d);
  assign {\lizzieLet33_4Lcall_main_map'_Int_Bool0_r ,
          es_2_2_destruct_r,
          es_3_4_destruct_r,
          es_4_7_destruct_r} = {4 {(\lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_r  && \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool,QTree_Bool) > (lizzieLet37_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_r ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_r  = ((! \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d [0]) || \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                                 1'd0};
    else
      if (\lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_r )
        \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d  <= \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_r  = (! \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet37_1_argbuf_d = (\lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf [0] ? \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                   1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                     1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_buf  <= \lizzieLet33_4Lcall_main_map'_Int_Bool0_1es_2_2_1es_3_4_1es_4_7_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Bool,
      Dcon Lcall_main_map'_Int_Bool0) : [(lizzieLet33_4Lcall_main_map'_Int_Bool1,Pointer_QTree_Bool),
                                         (es_3_3_destruct,Pointer_QTree_Bool),
                                         (es_4_6_destruct,Pointer_QTree_Bool),
                                         (sc_0_13_destruct,Pointer_CTmain_map'_Int_Bool)] > (lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0,CTmain_map'_Int_Bool) */
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_d  = \Lcall_main_map'_Int_Bool0_dc ((& {\lizzieLet33_4Lcall_main_map'_Int_Bool1_d [0],
                                                                                                                                             es_3_3_destruct_d[0],
                                                                                                                                             es_4_6_destruct_d[0],
                                                                                                                                             sc_0_13_destruct_d[0]}), \lizzieLet33_4Lcall_main_map'_Int_Bool1_d , es_3_3_destruct_d, es_4_6_destruct_d, sc_0_13_destruct_d);
  assign {\lizzieLet33_4Lcall_main_map'_Int_Bool1_r ,
          es_3_3_destruct_r,
          es_4_6_destruct_r,
          sc_0_13_destruct_r} = {4 {(\lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_r  && \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Bool) : (lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0,CTmain_map'_Int_Bool) > (lizzieLet36_1_argbuf,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_r ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_r  = ((! \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d [0]) || \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d  <= {67'd0,
                                                                                                                 1'd0};
    else
      if (\lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_r )
        \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d  <= \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_d ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_r  = (! \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf [0]);
  assign lizzieLet36_1_argbuf_d = (\lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf [0] ? \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf  :
                                   \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf  <= {67'd0,
                                                                                                                   1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf [0]))
        \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf  <= {67'd0,
                                                                                                                     1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf [0])))
        \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_buf  <= \lizzieLet33_4Lcall_main_map'_Int_Bool1_1es_3_3_1es_4_6_1sc_0_13_1Lcall_main_map'_Int_Bool0_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Bool,
      Dcon Lcall_main_map'_Int_Bool1) : [(lizzieLet33_4Lcall_main_map'_Int_Bool2,Pointer_QTree_Bool),
                                         (es_4_5_destruct,Pointer_QTree_Bool),
                                         (sc_0_12_destruct,Pointer_CTmain_map'_Int_Bool),
                                         (isZa8K_3_1,MyDTBool_Bool),
                                         (ga8L_3_1,MyDTInt_Bool),
                                         (q1a8O_2_destruct,Pointer_QTree_Int)] > (lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1,CTmain_map'_Int_Bool) */
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_d  = \Lcall_main_map'_Int_Bool1_dc ((& {\lizzieLet33_4Lcall_main_map'_Int_Bool2_d [0],
                                                                                                                                                                es_4_5_destruct_d[0],
                                                                                                                                                                sc_0_12_destruct_d[0],
                                                                                                                                                                isZa8K_3_1_d[0],
                                                                                                                                                                ga8L_3_1_d[0],
                                                                                                                                                                q1a8O_2_destruct_d[0]}), \lizzieLet33_4Lcall_main_map'_Int_Bool2_d , es_4_5_destruct_d, sc_0_12_destruct_d, isZa8K_3_1_d, ga8L_3_1_d, q1a8O_2_destruct_d);
  assign {\lizzieLet33_4Lcall_main_map'_Int_Bool2_r ,
          es_4_5_destruct_r,
          sc_0_12_destruct_r,
          isZa8K_3_1_r,
          ga8L_3_1_r,
          q1a8O_2_destruct_r} = {6 {(\lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_r  && \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Bool) : (lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1,CTmain_map'_Int_Bool) > (lizzieLet35_1_argbuf,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_r ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_r  = ((! \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d [0]) || \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d  <= {67'd0,
                                                                                                                                    1'd0};
    else
      if (\lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_r )
        \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d  <= \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_d ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_r  = (! \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf [0]);
  assign lizzieLet35_1_argbuf_d = (\lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf [0] ? \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf  :
                                   \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf  <= {67'd0,
                                                                                                                                      1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf [0]))
        \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf  <= {67'd0,
                                                                                                                                        1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf [0])))
        \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_buf  <= \lizzieLet33_4Lcall_main_map'_Int_Bool2_1es_4_5_1sc_0_12_1isZa8K_3_1ga8L_3_1q1a8O_2_1Lcall_main_map'_Int_Bool1_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Int_Bool,
      Dcon Lcall_main_map'_Int_Bool2) : [(lizzieLet33_4Lcall_main_map'_Int_Bool3,Pointer_QTree_Bool),
                                         (sc_0_11_destruct,Pointer_CTmain_map'_Int_Bool),
                                         (isZa8K_2_1,MyDTBool_Bool),
                                         (ga8L_2_1,MyDTInt_Bool),
                                         (q1a8O_1_destruct,Pointer_QTree_Int),
                                         (q2a8P_1_destruct,Pointer_QTree_Int)] > (lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2,CTmain_map'_Int_Bool) */
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_d  = \Lcall_main_map'_Int_Bool2_dc ((& {\lizzieLet33_4Lcall_main_map'_Int_Bool3_d [0],
                                                                                                                                                                 sc_0_11_destruct_d[0],
                                                                                                                                                                 isZa8K_2_1_d[0],
                                                                                                                                                                 ga8L_2_1_d[0],
                                                                                                                                                                 q1a8O_1_destruct_d[0],
                                                                                                                                                                 q2a8P_1_destruct_d[0]}), \lizzieLet33_4Lcall_main_map'_Int_Bool3_d , sc_0_11_destruct_d, isZa8K_2_1_d, ga8L_2_1_d, q1a8O_1_destruct_d, q2a8P_1_destruct_d);
  assign {\lizzieLet33_4Lcall_main_map'_Int_Bool3_r ,
          sc_0_11_destruct_r,
          isZa8K_2_1_r,
          ga8L_2_1_r,
          q1a8O_1_destruct_r,
          q2a8P_1_destruct_r} = {6 {(\lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_r  && \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_d [0])}};
  
  /* buf (Ty CTmain_map'_Int_Bool) : (lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2,CTmain_map'_Int_Bool) > (lizzieLet34_1_argbuf,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d ;
  logic \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_r ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_r  = ((! \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d [0]) || \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d  <= {67'd0,
                                                                                                                                     1'd0};
    else
      if (\lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_r )
        \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d  <= \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_d ;
  \CTmain_map'_Int_Bool_t  \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf ;
  assign \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_r  = (! \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf [0]);
  assign lizzieLet34_1_argbuf_d = (\lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf [0] ? \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf  :
                                   \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf  <= {67'd0,
                                                                                                                                       1'd0};
    else
      if ((lizzieLet34_1_argbuf_r && \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf [0]))
        \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf  <= {67'd0,
                                                                                                                                         1'd0};
      else if (((! lizzieLet34_1_argbuf_r) && (! \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf [0])))
        \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_buf  <= \lizzieLet33_4Lcall_main_map'_Int_Bool3_1sc_0_11_1isZa8K_2_1ga8L_2_1q1a8O_1_1q2a8P_1_1Lcall_main_map'_Int_Bool2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet33_4Lmain_map'_Int_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                            (lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted ;
  logic [1:0] \lizzieLet33_4Lmain_map'_Int_Boolsbos_done ;
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_d  = {\lizzieLet33_4Lmain_map'_Int_Boolsbos_d [16:1],
                                                                          (\lizzieLet33_4Lmain_map'_Int_Boolsbos_d [0] && (! \lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted [0]))};
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_d  = {\lizzieLet33_4Lmain_map'_Int_Boolsbos_d [16:1],
                                                                          (\lizzieLet33_4Lmain_map'_Int_Boolsbos_d [0] && (! \lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted [1]))};
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_done  = (\lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted  | ({\lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_d [0],
                                                                                                           \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_r  = (& \lizzieLet33_4Lmain_map'_Int_Boolsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted  <= 2'd0;
    else
      \lizzieLet33_4Lmain_map'_Int_Boolsbos_emitted  <= (\lizzieLet33_4Lmain_map'_Int_Boolsbos_r  ? 2'd0 :
                                                         \lizzieLet33_4Lmain_map'_Int_Boolsbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_main_map'_Int_Bool_goConst,Go) */
  assign \call_main_map'_Int_Bool_goConst_d  = \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_1_r  = \call_main_map'_Int_Bool_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (main_map'_Int_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_r )
        \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Bool_t \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \main_map'_Int_Bool_resbuf_d  = (\lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf  :
                                          \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((\main_map'_Int_Bool_resbuf_r  && \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! \main_map'_Int_Bool_resbuf_r ) && (! \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet33_4Lmain_map'_Int_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet4_1,MyBool) (arg0_2_1Dcon_main1_3I#_3,Go) > [(lizzieLet4_1MyFalse,Go),
                                                                       (lizzieLet4_1MyTrue,Go)] */
  logic [1:0] \arg0_2_1Dcon_main1_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet4_1_d[0] && \arg0_2_1Dcon_main1_3I#_3_d [0]))
      unique case (lizzieLet4_1_d[1:1])
        1'd0: \arg0_2_1Dcon_main1_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_2_1Dcon_main1_3I#_3_onehotd  = 2'd2;
        default: \arg0_2_1Dcon_main1_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_2_1Dcon_main1_3I#_3_onehotd  = 2'd0;
  assign lizzieLet4_1MyFalse_d = \arg0_2_1Dcon_main1_3I#_3_onehotd [0];
  assign lizzieLet4_1MyTrue_d = \arg0_2_1Dcon_main1_3I#_3_onehotd [1];
  assign \arg0_2_1Dcon_main1_3I#_3_r  = (| (\arg0_2_1Dcon_main1_3I#_3_onehotd  & {lizzieLet4_1MyTrue_r,
                                                                                  lizzieLet4_1MyFalse_r}));
  assign lizzieLet4_1_r = \arg0_2_1Dcon_main1_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet4_1MyFalse,Go)] > (lizzieLet4_1MyFalse_1MyTrue,MyBool) */
  assign lizzieLet4_1MyFalse_1MyTrue_d = MyTrue_dc((& {lizzieLet4_1MyFalse_d[0]}), lizzieLet4_1MyFalse_d);
  assign {lizzieLet4_1MyFalse_r} = {1 {(lizzieLet4_1MyFalse_1MyTrue_r && lizzieLet4_1MyFalse_1MyTrue_d[0])}};
  
  /* buf (Ty MyBool) : (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d;
  logic lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_r;
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_r = ((! lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d[0]) || lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d <= {1'd0,
                                                                                       1'd0};
    else
      if (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_r)
        lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d <= lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_d;
  MyBool_t lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf;
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_r = (! lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf[0] ? lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf :
                                       lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf <= {1'd0,
                                                                                         1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf[0]))
        lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf <= {1'd0,
                                                                                           1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf[0])))
        lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_buf <= lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet4_1MyTrue,Go)] > (lizzieLet4_1MyTrue_1MyFalse,MyBool) */
  assign lizzieLet4_1MyTrue_1MyFalse_d = MyFalse_dc((& {lizzieLet4_1MyTrue_d[0]}), lizzieLet4_1MyTrue_d);
  assign {lizzieLet4_1MyTrue_r} = {1 {(lizzieLet4_1MyTrue_1MyFalse_r && lizzieLet4_1MyTrue_1MyFalse_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet4_2,MyBool) [(lizzieLet4_1MyFalse_1MyTrue,MyBool),
                                         (lizzieLet4_1MyTrue_1MyFalse,MyBool)] > (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux,MyBool) */
  logic [1:0] lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux;
  logic [1:0] lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_onehot;
  always_comb
    unique case (lizzieLet4_2_d[1:1])
      1'd0:
        {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_onehot,
         lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux} = {2'd1,
                                                                            lizzieLet4_1MyFalse_1MyTrue_d};
      1'd1:
        {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_onehot,
         lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux} = {2'd2,
                                                                            lizzieLet4_1MyTrue_1MyFalse_d};
      default:
        {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_onehot,
         lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d = {lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux[1:1],
                                                                         (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_mux[0] && lizzieLet4_2_d[0])};
  assign lizzieLet4_2_r = (lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_d[0] && lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_r);
  assign {lizzieLet4_1MyTrue_1MyFalse_r,
          lizzieLet4_1MyFalse_1MyTrue_r} = (lizzieLet4_2_r ? lizzieLet4_1MyFalse_1MyTruelizzieLet4_1MyTrue_1MyFalse_mux_onehot :
                                            2'd0);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet5_1QNode_Int,QTree_Int) > [(q1a8j_destruct,Pointer_QTree_Int),
                                                                 (q2a8k_destruct,Pointer_QTree_Int),
                                                                 (q3a8l_destruct,Pointer_QTree_Int),
                                                                 (q4a8m_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet5_1QNode_Int_emitted;
  logic [3:0] lizzieLet5_1QNode_Int_done;
  assign q1a8j_destruct_d = {lizzieLet5_1QNode_Int_d[18:3],
                             (lizzieLet5_1QNode_Int_d[0] && (! lizzieLet5_1QNode_Int_emitted[0]))};
  assign q2a8k_destruct_d = {lizzieLet5_1QNode_Int_d[34:19],
                             (lizzieLet5_1QNode_Int_d[0] && (! lizzieLet5_1QNode_Int_emitted[1]))};
  assign q3a8l_destruct_d = {lizzieLet5_1QNode_Int_d[50:35],
                             (lizzieLet5_1QNode_Int_d[0] && (! lizzieLet5_1QNode_Int_emitted[2]))};
  assign q4a8m_destruct_d = {lizzieLet5_1QNode_Int_d[66:51],
                             (lizzieLet5_1QNode_Int_d[0] && (! lizzieLet5_1QNode_Int_emitted[3]))};
  assign lizzieLet5_1QNode_Int_done = (lizzieLet5_1QNode_Int_emitted | ({q4a8m_destruct_d[0],
                                                                         q3a8l_destruct_d[0],
                                                                         q2a8k_destruct_d[0],
                                                                         q1a8j_destruct_d[0]} & {q4a8m_destruct_r,
                                                                                                 q3a8l_destruct_r,
                                                                                                 q2a8k_destruct_r,
                                                                                                 q1a8j_destruct_r}));
  assign lizzieLet5_1QNode_Int_r = (& lizzieLet5_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet5_1QNode_Int_emitted <= (lizzieLet5_1QNode_Int_r ? 4'd0 :
                                        lizzieLet5_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet5_1QVal_Int,QTree_Int) > [(v1a8d_destruct,Int)] */
  assign v1a8d_destruct_d = {lizzieLet5_1QVal_Int_d[34:3],
                             lizzieLet5_1QVal_Int_d[0]};
  assign lizzieLet5_1QVal_Int_r = v1a8d_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet5_2,QTree_Int) (lizzieLet5_1,QTree_Int) > [(_43,QTree_Int),
                                                                            (lizzieLet5_1QVal_Int,QTree_Int),
                                                                            (lizzieLet5_1QNode_Int,QTree_Int),
                                                                            (_42,QTree_Int)] */
  logic [3:0] lizzieLet5_1_onehotd;
  always_comb
    if ((lizzieLet5_2_d[0] && lizzieLet5_1_d[0]))
      unique case (lizzieLet5_2_d[2:1])
        2'd0: lizzieLet5_1_onehotd = 4'd1;
        2'd1: lizzieLet5_1_onehotd = 4'd2;
        2'd2: lizzieLet5_1_onehotd = 4'd4;
        2'd3: lizzieLet5_1_onehotd = 4'd8;
        default: lizzieLet5_1_onehotd = 4'd0;
      endcase
    else lizzieLet5_1_onehotd = 4'd0;
  assign _43_d = {lizzieLet5_1_d[66:1], lizzieLet5_1_onehotd[0]};
  assign lizzieLet5_1QVal_Int_d = {lizzieLet5_1_d[66:1],
                                   lizzieLet5_1_onehotd[1]};
  assign lizzieLet5_1QNode_Int_d = {lizzieLet5_1_d[66:1],
                                    lizzieLet5_1_onehotd[2]};
  assign _42_d = {lizzieLet5_1_d[66:1], lizzieLet5_1_onehotd[3]};
  assign lizzieLet5_1_r = (| (lizzieLet5_1_onehotd & {_42_r,
                                                      lizzieLet5_1QNode_Int_r,
                                                      lizzieLet5_1QVal_Int_r,
                                                      _43_r}));
  assign lizzieLet5_2_r = lizzieLet5_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet5_3,QTree_Int) (go_11_goMux_data,Go) > [(lizzieLet5_3QNone_Int,Go),
                                                                  (lizzieLet5_3QVal_Int,Go),
                                                                  (lizzieLet5_3QNode_Int,Go),
                                                                  (lizzieLet5_3QError_Int,Go)] */
  logic [3:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet5_3_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet5_3_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 4'd1;
        2'd1: go_11_goMux_data_onehotd = 4'd2;
        2'd2: go_11_goMux_data_onehotd = 4'd4;
        2'd3: go_11_goMux_data_onehotd = 4'd8;
        default: go_11_goMux_data_onehotd = 4'd0;
      endcase
    else go_11_goMux_data_onehotd = 4'd0;
  assign lizzieLet5_3QNone_Int_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet5_3QVal_Int_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet5_3QNode_Int_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet5_3QError_Int_d = go_11_goMux_data_onehotd[3];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet5_3QError_Int_r,
                                                              lizzieLet5_3QNode_Int_r,
                                                              lizzieLet5_3QVal_Int_r,
                                                              lizzieLet5_3QNone_Int_r}));
  assign lizzieLet5_3_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet5_3QError_Int,Go) > [(lizzieLet5_3QError_Int_1,Go),
                                              (lizzieLet5_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet5_3QError_Int_emitted;
  logic [1:0] lizzieLet5_3QError_Int_done;
  assign lizzieLet5_3QError_Int_1_d = (lizzieLet5_3QError_Int_d[0] && (! lizzieLet5_3QError_Int_emitted[0]));
  assign lizzieLet5_3QError_Int_2_d = (lizzieLet5_3QError_Int_d[0] && (! lizzieLet5_3QError_Int_emitted[1]));
  assign lizzieLet5_3QError_Int_done = (lizzieLet5_3QError_Int_emitted | ({lizzieLet5_3QError_Int_2_d[0],
                                                                           lizzieLet5_3QError_Int_1_d[0]} & {lizzieLet5_3QError_Int_2_r,
                                                                                                             lizzieLet5_3QError_Int_1_r}));
  assign lizzieLet5_3QError_Int_r = (& lizzieLet5_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet5_3QError_Int_emitted <= (lizzieLet5_3QError_Int_r ? 2'd0 :
                                         lizzieLet5_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet5_3QError_Int_1,Go)] > (lizzieLet5_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet5_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet5_3QError_Int_1_d[0]}), lizzieLet5_3QError_Int_1_d);
  assign {lizzieLet5_3QError_Int_1_r} = {1 {(lizzieLet5_3QError_Int_1QError_Int_r && lizzieLet5_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet5_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet14_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet5_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet5_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet5_3QError_Int_1QError_Int_r = ((! lizzieLet5_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet5_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_3QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet5_3QError_Int_1QError_Int_r)
        lizzieLet5_3QError_Int_1QError_Int_bufchan_d <= lizzieLet5_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet5_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet5_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet5_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (lizzieLet5_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet5_3QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet5_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && lizzieLet5_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet5_3QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! lizzieLet5_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet5_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet5_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_3QError_Int_2,Go) > (lizzieLet5_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet5_3QError_Int_2_bufchan_d;
  logic lizzieLet5_3QError_Int_2_bufchan_r;
  assign lizzieLet5_3QError_Int_2_r = ((! lizzieLet5_3QError_Int_2_bufchan_d[0]) || lizzieLet5_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_3QError_Int_2_r)
        lizzieLet5_3QError_Int_2_bufchan_d <= lizzieLet5_3QError_Int_2_d;
  Go_t lizzieLet5_3QError_Int_2_bufchan_buf;
  assign lizzieLet5_3QError_Int_2_bufchan_r = (! lizzieLet5_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet5_3QError_Int_2_argbuf_d = (lizzieLet5_3QError_Int_2_bufchan_buf[0] ? lizzieLet5_3QError_Int_2_bufchan_buf :
                                              lizzieLet5_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_3QError_Int_2_argbuf_r && lizzieLet5_3QError_Int_2_bufchan_buf[0]))
        lizzieLet5_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_3QError_Int_2_argbuf_r) && (! lizzieLet5_3QError_Int_2_bufchan_buf[0])))
        lizzieLet5_3QError_Int_2_bufchan_buf <= lizzieLet5_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_3QNone_Int,Go) > (lizzieLet5_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet5_3QNone_Int_bufchan_d;
  logic lizzieLet5_3QNone_Int_bufchan_r;
  assign lizzieLet5_3QNone_Int_r = ((! lizzieLet5_3QNone_Int_bufchan_d[0]) || lizzieLet5_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_3QNone_Int_r)
        lizzieLet5_3QNone_Int_bufchan_d <= lizzieLet5_3QNone_Int_d;
  Go_t lizzieLet5_3QNone_Int_bufchan_buf;
  assign lizzieLet5_3QNone_Int_bufchan_r = (! lizzieLet5_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_3QNone_Int_1_argbuf_d = (lizzieLet5_3QNone_Int_bufchan_buf[0] ? lizzieLet5_3QNone_Int_bufchan_buf :
                                             lizzieLet5_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_3QNone_Int_1_argbuf_r && lizzieLet5_3QNone_Int_bufchan_buf[0]))
        lizzieLet5_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_3QNone_Int_1_argbuf_r) && (! lizzieLet5_3QNone_Int_bufchan_buf[0])))
        lizzieLet5_3QNone_Int_bufchan_buf <= lizzieLet5_3QNone_Int_bufchan_d;
  
  /* mergectrl (Ty C10,Ty Go) : [(lizzieLet5_3QNone_Int_1_argbuf,Go),
                            (lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf,Go),
                            (lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf,Go),
                            (lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf,Go),
                            (lizzieLet5_4QVal_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf,Go),
                            (lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf,Go),
                            (lizzieLet5_4QNode_Int_3QError_Int_2_argbuf,Go),
                            (lizzieLet5_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C10) (go_15_goMux_data,Go) */
  logic [9:0] lizzieLet5_3QNone_Int_1_argbuf_select_d;
  assign lizzieLet5_3QNone_Int_1_argbuf_select_d = ((| lizzieLet5_3QNone_Int_1_argbuf_select_q) ? lizzieLet5_3QNone_Int_1_argbuf_select_q :
                                                    (lizzieLet5_3QNone_Int_1_argbuf_d[0] ? 10'd1 :
                                                     (lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_d[0] ? 10'd2 :
                                                      (lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_d[0] ? 10'd4 :
                                                       (lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_d[0] ? 10'd8 :
                                                        (lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_d[0] ? 10'd16 :
                                                         (lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_d[0] ? 10'd32 :
                                                          (lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_d[0] ? 10'd64 :
                                                           (lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_d[0] ? 10'd128 :
                                                            (lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_d[0] ? 10'd256 :
                                                             (lizzieLet5_3QError_Int_2_argbuf_d[0] ? 10'd512 :
                                                              10'd0)))))))))));
  logic [9:0] lizzieLet5_3QNone_Int_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_3QNone_Int_1_argbuf_select_q <= 10'd0;
    else
      lizzieLet5_3QNone_Int_1_argbuf_select_q <= (lizzieLet5_3QNone_Int_1_argbuf_done ? 10'd0 :
                                                  lizzieLet5_3QNone_Int_1_argbuf_select_d);
  logic [1:0] lizzieLet5_3QNone_Int_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_3QNone_Int_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet5_3QNone_Int_1_argbuf_emit_q <= (lizzieLet5_3QNone_Int_1_argbuf_done ? 2'd0 :
                                                lizzieLet5_3QNone_Int_1_argbuf_emit_d);
  logic [1:0] lizzieLet5_3QNone_Int_1_argbuf_emit_d;
  assign lizzieLet5_3QNone_Int_1_argbuf_emit_d = (lizzieLet5_3QNone_Int_1_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                            go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                      go_15_goMux_data_r}));
  logic lizzieLet5_3QNone_Int_1_argbuf_done;
  assign lizzieLet5_3QNone_Int_1_argbuf_done = (& lizzieLet5_3QNone_Int_1_argbuf_emit_d);
  assign {lizzieLet5_3QError_Int_2_argbuf_r,
          lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_r,
          lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_r,
          lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_r,
          lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_r,
          lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_r,
          lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_r,
          lizzieLet5_3QNone_Int_1_argbuf_r} = (lizzieLet5_3QNone_Int_1_argbuf_done ? lizzieLet5_3QNone_Int_1_argbuf_select_d :
                                               10'd0);
  assign go_15_goMux_data_d = ((lizzieLet5_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_3QNone_Int_1_argbuf_d :
                               ((lizzieLet5_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet24_3Lcall_$wmAdd_Int0_1_argbuf_d :
                                ((lizzieLet5_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_d :
                                 ((lizzieLet5_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_d :
                                  ((lizzieLet5_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_d :
                                   ((lizzieLet5_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_d :
                                    ((lizzieLet5_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_d :
                                     ((lizzieLet5_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_d :
                                      ((lizzieLet5_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_d :
                                       ((lizzieLet5_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[0])) ? lizzieLet5_3QError_Int_2_argbuf_d :
                                        1'd0))))))))));
  assign go_15_goMux_choice_d = ((lizzieLet5_3QNone_Int_1_argbuf_select_d[0] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C1_10_dc(1'd1) :
                                 ((lizzieLet5_3QNone_Int_1_argbuf_select_d[1] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C2_10_dc(1'd1) :
                                  ((lizzieLet5_3QNone_Int_1_argbuf_select_d[2] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C3_10_dc(1'd1) :
                                   ((lizzieLet5_3QNone_Int_1_argbuf_select_d[3] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C4_10_dc(1'd1) :
                                    ((lizzieLet5_3QNone_Int_1_argbuf_select_d[4] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C5_10_dc(1'd1) :
                                     ((lizzieLet5_3QNone_Int_1_argbuf_select_d[5] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C6_10_dc(1'd1) :
                                      ((lizzieLet5_3QNone_Int_1_argbuf_select_d[6] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C7_10_dc(1'd1) :
                                       ((lizzieLet5_3QNone_Int_1_argbuf_select_d[7] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C8_10_dc(1'd1) :
                                        ((lizzieLet5_3QNone_Int_1_argbuf_select_d[8] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C9_10_dc(1'd1) :
                                         ((lizzieLet5_3QNone_Int_1_argbuf_select_d[9] && (! lizzieLet5_3QNone_Int_1_argbuf_emit_q[1])) ? C10_10_dc(1'd1) :
                                          {4'd0, 1'd0}))))))))));
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet5_4,QTree_Int) (readPointer_QTree_Intw2slT_1_1_argbuf_rwb,QTree_Int) > [(_41,QTree_Int),
                                                                                                         (lizzieLet5_4QVal_Int,QTree_Int),
                                                                                                         (lizzieLet5_4QNode_Int,QTree_Int),
                                                                                                         (_40,QTree_Int)] */
  logic [3:0] readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet5_4_d[0] && readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d[0]))
      unique case (lizzieLet5_4_d[2:1])
        2'd0: readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd = 4'd0;
  assign _41_d = {readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet5_4QVal_Int_d = {readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d[66:1],
                                   readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet5_4QNode_Int_d = {readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd[2]};
  assign _40_d = {readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Intw2slT_1_1_argbuf_rwb_r = (| (readPointer_QTree_Intw2slT_1_1_argbuf_rwb_onehotd & {_40_r,
                                                                                                                lizzieLet5_4QNode_Int_r,
                                                                                                                lizzieLet5_4QVal_Int_r,
                                                                                                                _41_r}));
  assign lizzieLet5_4_r = readPointer_QTree_Intw2slT_1_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet5_4QNode_Int,QTree_Int) > [(lizzieLet5_4QNode_Int_1,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_2,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_3,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_4,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_5,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_6,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_7,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_8,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_9,QTree_Int),
                                                           (lizzieLet5_4QNode_Int_10,QTree_Int)] */
  logic [9:0] lizzieLet5_4QNode_Int_emitted;
  logic [9:0] lizzieLet5_4QNode_Int_done;
  assign lizzieLet5_4QNode_Int_1_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[0]))};
  assign lizzieLet5_4QNode_Int_2_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[1]))};
  assign lizzieLet5_4QNode_Int_3_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[2]))};
  assign lizzieLet5_4QNode_Int_4_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[3]))};
  assign lizzieLet5_4QNode_Int_5_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[4]))};
  assign lizzieLet5_4QNode_Int_6_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[5]))};
  assign lizzieLet5_4QNode_Int_7_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[6]))};
  assign lizzieLet5_4QNode_Int_8_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[7]))};
  assign lizzieLet5_4QNode_Int_9_d = {lizzieLet5_4QNode_Int_d[66:1],
                                      (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[8]))};
  assign lizzieLet5_4QNode_Int_10_d = {lizzieLet5_4QNode_Int_d[66:1],
                                       (lizzieLet5_4QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_emitted[9]))};
  assign lizzieLet5_4QNode_Int_done = (lizzieLet5_4QNode_Int_emitted | ({lizzieLet5_4QNode_Int_10_d[0],
                                                                         lizzieLet5_4QNode_Int_9_d[0],
                                                                         lizzieLet5_4QNode_Int_8_d[0],
                                                                         lizzieLet5_4QNode_Int_7_d[0],
                                                                         lizzieLet5_4QNode_Int_6_d[0],
                                                                         lizzieLet5_4QNode_Int_5_d[0],
                                                                         lizzieLet5_4QNode_Int_4_d[0],
                                                                         lizzieLet5_4QNode_Int_3_d[0],
                                                                         lizzieLet5_4QNode_Int_2_d[0],
                                                                         lizzieLet5_4QNode_Int_1_d[0]} & {lizzieLet5_4QNode_Int_10_r,
                                                                                                          lizzieLet5_4QNode_Int_9_r,
                                                                                                          lizzieLet5_4QNode_Int_8_r,
                                                                                                          lizzieLet5_4QNode_Int_7_r,
                                                                                                          lizzieLet5_4QNode_Int_6_r,
                                                                                                          lizzieLet5_4QNode_Int_5_r,
                                                                                                          lizzieLet5_4QNode_Int_4_r,
                                                                                                          lizzieLet5_4QNode_Int_3_r,
                                                                                                          lizzieLet5_4QNode_Int_2_r,
                                                                                                          lizzieLet5_4QNode_Int_1_r}));
  assign lizzieLet5_4QNode_Int_r = (& lizzieLet5_4QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_4QNode_Int_emitted <= 10'd0;
    else
      lizzieLet5_4QNode_Int_emitted <= (lizzieLet5_4QNode_Int_r ? 10'd0 :
                                        lizzieLet5_4QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_10,QTree_Int) (q4a8m_destruct,Pointer_QTree_Int) > [(_39,Pointer_QTree_Int),
                                                                                                          (_38,Pointer_QTree_Int),
                                                                                                          (lizzieLet5_4QNode_Int_10QNode_Int,Pointer_QTree_Int),
                                                                                                          (_37,Pointer_QTree_Int)] */
  logic [3:0] q4a8m_destruct_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_10_d[0] && q4a8m_destruct_d[0]))
      unique case (lizzieLet5_4QNode_Int_10_d[2:1])
        2'd0: q4a8m_destruct_onehotd = 4'd1;
        2'd1: q4a8m_destruct_onehotd = 4'd2;
        2'd2: q4a8m_destruct_onehotd = 4'd4;
        2'd3: q4a8m_destruct_onehotd = 4'd8;
        default: q4a8m_destruct_onehotd = 4'd0;
      endcase
    else q4a8m_destruct_onehotd = 4'd0;
  assign _39_d = {q4a8m_destruct_d[16:1], q4a8m_destruct_onehotd[0]};
  assign _38_d = {q4a8m_destruct_d[16:1], q4a8m_destruct_onehotd[1]};
  assign lizzieLet5_4QNode_Int_10QNode_Int_d = {q4a8m_destruct_d[16:1],
                                                q4a8m_destruct_onehotd[2]};
  assign _37_d = {q4a8m_destruct_d[16:1], q4a8m_destruct_onehotd[3]};
  assign q4a8m_destruct_r = (| (q4a8m_destruct_onehotd & {_37_r,
                                                          lizzieLet5_4QNode_Int_10QNode_Int_r,
                                                          _38_r,
                                                          _39_r}));
  assign lizzieLet5_4QNode_Int_10_r = q4a8m_destruct_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_10QNode_Int,Pointer_QTree_Int) > (lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_10QNode_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_10QNode_Int_r = ((! lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_10QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QNode_Int_10QNode_Int_r)
        lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d <= lizzieLet5_4QNode_Int_10QNode_Int_d;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_10QNode_Int_bufchan_r = (! lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf :
                                                         lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_r && lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QNode_Int_10QNode_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_10QNode_Int_bufchan_buf <= lizzieLet5_4QNode_Int_10QNode_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet5_4QNode_Int_1QNode_Int,QTree_Int) > [(t1a8o_destruct,Pointer_QTree_Int),
                                                                            (t2a8p_destruct,Pointer_QTree_Int),
                                                                            (t3a8q_destruct,Pointer_QTree_Int),
                                                                            (t4a8r_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet5_4QNode_Int_1QNode_Int_emitted;
  logic [3:0] lizzieLet5_4QNode_Int_1QNode_Int_done;
  assign t1a8o_destruct_d = {lizzieLet5_4QNode_Int_1QNode_Int_d[18:3],
                             (lizzieLet5_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_1QNode_Int_emitted[0]))};
  assign t2a8p_destruct_d = {lizzieLet5_4QNode_Int_1QNode_Int_d[34:19],
                             (lizzieLet5_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_1QNode_Int_emitted[1]))};
  assign t3a8q_destruct_d = {lizzieLet5_4QNode_Int_1QNode_Int_d[50:35],
                             (lizzieLet5_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_1QNode_Int_emitted[2]))};
  assign t4a8r_destruct_d = {lizzieLet5_4QNode_Int_1QNode_Int_d[66:51],
                             (lizzieLet5_4QNode_Int_1QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_1QNode_Int_emitted[3]))};
  assign lizzieLet5_4QNode_Int_1QNode_Int_done = (lizzieLet5_4QNode_Int_1QNode_Int_emitted | ({t4a8r_destruct_d[0],
                                                                                               t3a8q_destruct_d[0],
                                                                                               t2a8p_destruct_d[0],
                                                                                               t1a8o_destruct_d[0]} & {t4a8r_destruct_r,
                                                                                                                       t3a8q_destruct_r,
                                                                                                                       t2a8p_destruct_r,
                                                                                                                       t1a8o_destruct_r}));
  assign lizzieLet5_4QNode_Int_1QNode_Int_r = (& lizzieLet5_4QNode_Int_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet5_4QNode_Int_1QNode_Int_emitted <= (lizzieLet5_4QNode_Int_1QNode_Int_r ? 4'd0 :
                                                   lizzieLet5_4QNode_Int_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet5_4QNode_Int_2,QTree_Int) (lizzieLet5_4QNode_Int_1,QTree_Int) > [(_36,QTree_Int),
                                                                                                  (_35,QTree_Int),
                                                                                                  (lizzieLet5_4QNode_Int_1QNode_Int,QTree_Int),
                                                                                                  (_34,QTree_Int)] */
  logic [3:0] lizzieLet5_4QNode_Int_1_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_2_d[0] && lizzieLet5_4QNode_Int_1_d[0]))
      unique case (lizzieLet5_4QNode_Int_2_d[2:1])
        2'd0: lizzieLet5_4QNode_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet5_4QNode_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet5_4QNode_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet5_4QNode_Int_1_onehotd = 4'd8;
        default: lizzieLet5_4QNode_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet5_4QNode_Int_1_onehotd = 4'd0;
  assign _36_d = {lizzieLet5_4QNode_Int_1_d[66:1],
                  lizzieLet5_4QNode_Int_1_onehotd[0]};
  assign _35_d = {lizzieLet5_4QNode_Int_1_d[66:1],
                  lizzieLet5_4QNode_Int_1_onehotd[1]};
  assign lizzieLet5_4QNode_Int_1QNode_Int_d = {lizzieLet5_4QNode_Int_1_d[66:1],
                                               lizzieLet5_4QNode_Int_1_onehotd[2]};
  assign _34_d = {lizzieLet5_4QNode_Int_1_d[66:1],
                  lizzieLet5_4QNode_Int_1_onehotd[3]};
  assign lizzieLet5_4QNode_Int_1_r = (| (lizzieLet5_4QNode_Int_1_onehotd & {_34_r,
                                                                            lizzieLet5_4QNode_Int_1QNode_Int_r,
                                                                            _35_r,
                                                                            _36_r}));
  assign lizzieLet5_4QNode_Int_2_r = lizzieLet5_4QNode_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet5_4QNode_Int_3,QTree_Int) (lizzieLet5_3QNode_Int,Go) > [(lizzieLet5_4QNode_Int_3QNone_Int,Go),
                                                                                  (lizzieLet5_4QNode_Int_3QVal_Int,Go),
                                                                                  (lizzieLet5_4QNode_Int_3QNode_Int,Go),
                                                                                  (lizzieLet5_4QNode_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet5_3QNode_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_3_d[0] && lizzieLet5_3QNode_Int_d[0]))
      unique case (lizzieLet5_4QNode_Int_3_d[2:1])
        2'd0: lizzieLet5_3QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_3QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_3QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_3QNode_Int_onehotd = 4'd8;
        default: lizzieLet5_3QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_3QNode_Int_onehotd = 4'd0;
  assign lizzieLet5_4QNode_Int_3QNone_Int_d = lizzieLet5_3QNode_Int_onehotd[0];
  assign lizzieLet5_4QNode_Int_3QVal_Int_d = lizzieLet5_3QNode_Int_onehotd[1];
  assign lizzieLet5_4QNode_Int_3QNode_Int_d = lizzieLet5_3QNode_Int_onehotd[2];
  assign lizzieLet5_4QNode_Int_3QError_Int_d = lizzieLet5_3QNode_Int_onehotd[3];
  assign lizzieLet5_3QNode_Int_r = (| (lizzieLet5_3QNode_Int_onehotd & {lizzieLet5_4QNode_Int_3QError_Int_r,
                                                                        lizzieLet5_4QNode_Int_3QNode_Int_r,
                                                                        lizzieLet5_4QNode_Int_3QVal_Int_r,
                                                                        lizzieLet5_4QNode_Int_3QNone_Int_r}));
  assign lizzieLet5_4QNode_Int_3_r = lizzieLet5_3QNode_Int_r;
  
  /* fork (Ty Go) : (lizzieLet5_4QNode_Int_3QError_Int,Go) > [(lizzieLet5_4QNode_Int_3QError_Int_1,Go),
                                                         (lizzieLet5_4QNode_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet5_4QNode_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet5_4QNode_Int_3QError_Int_done;
  assign lizzieLet5_4QNode_Int_3QError_Int_1_d = (lizzieLet5_4QNode_Int_3QError_Int_d[0] && (! lizzieLet5_4QNode_Int_3QError_Int_emitted[0]));
  assign lizzieLet5_4QNode_Int_3QError_Int_2_d = (lizzieLet5_4QNode_Int_3QError_Int_d[0] && (! lizzieLet5_4QNode_Int_3QError_Int_emitted[1]));
  assign lizzieLet5_4QNode_Int_3QError_Int_done = (lizzieLet5_4QNode_Int_3QError_Int_emitted | ({lizzieLet5_4QNode_Int_3QError_Int_2_d[0],
                                                                                                 lizzieLet5_4QNode_Int_3QError_Int_1_d[0]} & {lizzieLet5_4QNode_Int_3QError_Int_2_r,
                                                                                                                                              lizzieLet5_4QNode_Int_3QError_Int_1_r}));
  assign lizzieLet5_4QNode_Int_3QError_Int_r = (& lizzieLet5_4QNode_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet5_4QNode_Int_3QError_Int_emitted <= (lizzieLet5_4QNode_Int_3QError_Int_r ? 2'd0 :
                                                    lizzieLet5_4QNode_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet5_4QNode_Int_3QError_Int_1,Go)] > (lizzieLet5_4QNode_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet5_4QNode_Int_3QError_Int_1_d[0]}), lizzieLet5_4QNode_Int_3QError_Int_1_d);
  assign {lizzieLet5_4QNode_Int_3QError_Int_1_r} = {1 {(lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_r && lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet5_4QNode_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet13_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_r = ((! lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_r)
        lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet5_4QNode_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QNode_Int_3QError_Int_2,Go) > (lizzieLet5_4QNode_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QError_Int_2_r = ((! lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QNode_Int_3QError_Int_2_r)
        lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d <= lizzieLet5_4QNode_Int_3QError_Int_2_d;
  Go_t lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_r = (! lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_d = (lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf :
                                                         lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_r && lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QNode_Int_3QError_Int_2_argbuf_r) && (! lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_buf <= lizzieLet5_4QNode_Int_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QNode_Int_3QNode_Int,Go) > (lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QNode_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QNode_Int_r = ((! lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QNode_Int_3QNode_Int_r)
        lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d <= lizzieLet5_4QNode_Int_3QNode_Int_d;
  Go_t lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QNode_Int_bufchan_r = (! lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf :
                                                        lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_r && lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QNode_Int_3QNode_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QNode_Int_bufchan_buf <= lizzieLet5_4QNode_Int_3QNode_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QNode_Int_3QNone_Int,Go) > (lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QNone_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QNone_Int_r = ((! lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QNode_Int_3QNone_Int_r)
        lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d <= lizzieLet5_4QNode_Int_3QNone_Int_d;
  Go_t lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QNone_Int_bufchan_r = (! lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf :
                                                        lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_r && lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QNode_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QNone_Int_bufchan_buf <= lizzieLet5_4QNode_Int_3QNone_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet5_4QNode_Int_3QVal_Int,Go) > [(lizzieLet5_4QNode_Int_3QVal_Int_1,Go),
                                                       (lizzieLet5_4QNode_Int_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet5_4QNode_Int_3QVal_Int_emitted;
  logic [1:0] lizzieLet5_4QNode_Int_3QVal_Int_done;
  assign lizzieLet5_4QNode_Int_3QVal_Int_1_d = (lizzieLet5_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet5_4QNode_Int_3QVal_Int_emitted[0]));
  assign lizzieLet5_4QNode_Int_3QVal_Int_2_d = (lizzieLet5_4QNode_Int_3QVal_Int_d[0] && (! lizzieLet5_4QNode_Int_3QVal_Int_emitted[1]));
  assign lizzieLet5_4QNode_Int_3QVal_Int_done = (lizzieLet5_4QNode_Int_3QVal_Int_emitted | ({lizzieLet5_4QNode_Int_3QVal_Int_2_d[0],
                                                                                             lizzieLet5_4QNode_Int_3QVal_Int_1_d[0]} & {lizzieLet5_4QNode_Int_3QVal_Int_2_r,
                                                                                                                                        lizzieLet5_4QNode_Int_3QVal_Int_1_r}));
  assign lizzieLet5_4QNode_Int_3QVal_Int_r = (& lizzieLet5_4QNode_Int_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet5_4QNode_Int_3QVal_Int_emitted <= (lizzieLet5_4QNode_Int_3QVal_Int_r ? 2'd0 :
                                                  lizzieLet5_4QNode_Int_3QVal_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet5_4QNode_Int_3QVal_Int_1,Go)] > (lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int,QTree_Int) */
  assign lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet5_4QNode_Int_3QVal_Int_1_d[0]}), lizzieLet5_4QNode_Int_3QVal_Int_1_d);
  assign {lizzieLet5_4QNode_Int_3QVal_Int_1_r} = {1 {(lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_r && lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int,QTree_Int) > (lizzieLet11_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_r = ((! lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_r)
        lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d <= lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_d;
  QTree_Int_t lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_r = (! lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf :
                                     lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_buf <= lizzieLet5_4QNode_Int_3QVal_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QNode_Int_3QVal_Int_2,Go) > (lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d;
  logic lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_r;
  assign lizzieLet5_4QNode_Int_3QVal_Int_2_r = ((! lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d[0]) || lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QNode_Int_3QVal_Int_2_r)
        lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d <= lizzieLet5_4QNode_Int_3QVal_Int_2_d;
  Go_t lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf;
  assign lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_r = (! lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_d = (lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf[0] ? lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf :
                                                       lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_r && lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QNode_Int_3QVal_Int_2_argbuf_r) && (! lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_buf <= lizzieLet5_4QNode_Int_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QNode_Int_4,QTree_Int) (lizzieLet5_5QNode_Int,Pointer_CT$wmAdd_Int) > [(lizzieLet5_4QNode_Int_4QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet5_4QNode_Int_4QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet5_4QNode_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                                      (lizzieLet5_4QNode_Int_4QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet5_5QNode_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_4_d[0] && lizzieLet5_5QNode_Int_d[0]))
      unique case (lizzieLet5_4QNode_Int_4_d[2:1])
        2'd0: lizzieLet5_5QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_5QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_5QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_5QNode_Int_onehotd = 4'd8;
        default: lizzieLet5_5QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_5QNode_Int_onehotd = 4'd0;
  assign lizzieLet5_4QNode_Int_4QNone_Int_d = {lizzieLet5_5QNode_Int_d[16:1],
                                               lizzieLet5_5QNode_Int_onehotd[0]};
  assign lizzieLet5_4QNode_Int_4QVal_Int_d = {lizzieLet5_5QNode_Int_d[16:1],
                                              lizzieLet5_5QNode_Int_onehotd[1]};
  assign lizzieLet5_4QNode_Int_4QNode_Int_d = {lizzieLet5_5QNode_Int_d[16:1],
                                               lizzieLet5_5QNode_Int_onehotd[2]};
  assign lizzieLet5_4QNode_Int_4QError_Int_d = {lizzieLet5_5QNode_Int_d[16:1],
                                                lizzieLet5_5QNode_Int_onehotd[3]};
  assign lizzieLet5_5QNode_Int_r = (| (lizzieLet5_5QNode_Int_onehotd & {lizzieLet5_4QNode_Int_4QError_Int_r,
                                                                        lizzieLet5_4QNode_Int_4QNode_Int_r,
                                                                        lizzieLet5_4QNode_Int_4QVal_Int_r,
                                                                        lizzieLet5_4QNode_Int_4QNone_Int_r}));
  assign lizzieLet5_4QNode_Int_4_r = lizzieLet5_5QNode_Int_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QNode_Int_4QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QNode_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QError_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_4QError_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_4QError_Int_r = ((! lizzieLet5_4QNode_Int_4QError_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QNode_Int_4QError_Int_r)
        lizzieLet5_4QNode_Int_4QError_Int_bufchan_d <= lizzieLet5_4QNode_Int_4QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_4QError_Int_bufchan_r = (! lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf :
                                                         lizzieLet5_4QNode_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_r && lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QNode_Int_4QError_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_4QError_Int_bufchan_buf <= lizzieLet5_4QNode_Int_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Int,
      Dcon Lcall_$wmAdd_Int3) : [(lizzieLet5_4QNode_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                 (lizzieLet5_4QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                 (lizzieLet5_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                                 (t1a8o_destruct,Pointer_QTree_Int),
                                 (lizzieLet5_4QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                 (t2a8p_destruct,Pointer_QTree_Int),
                                 (lizzieLet5_4QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                 (t3a8q_destruct,Pointer_QTree_Int)] > (lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) */
  assign lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_d = Lcall_$wmAdd_Int3_dc((& {lizzieLet5_4QNode_Int_4QNode_Int_d[0],
                                                                                                                                                                                                                                                       lizzieLet5_4QNode_Int_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                       lizzieLet5_4QNode_Int_7QNode_Int_d[0],
                                                                                                                                                                                                                                                       t1a8o_destruct_d[0],
                                                                                                                                                                                                                                                       lizzieLet5_4QNode_Int_8QNode_Int_d[0],
                                                                                                                                                                                                                                                       t2a8p_destruct_d[0],
                                                                                                                                                                                                                                                       lizzieLet5_4QNode_Int_9QNode_Int_d[0],
                                                                                                                                                                                                                                                       t3a8q_destruct_d[0]}), lizzieLet5_4QNode_Int_4QNode_Int_d, lizzieLet5_4QNode_Int_6QNode_Int_1_d, lizzieLet5_4QNode_Int_7QNode_Int_d, t1a8o_destruct_d, lizzieLet5_4QNode_Int_8QNode_Int_d, t2a8p_destruct_d, lizzieLet5_4QNode_Int_9QNode_Int_d, t3a8q_destruct_d);
  assign {lizzieLet5_4QNode_Int_4QNode_Int_r,
          lizzieLet5_4QNode_Int_6QNode_Int_1_r,
          lizzieLet5_4QNode_Int_7QNode_Int_r,
          t1a8o_destruct_r,
          lizzieLet5_4QNode_Int_8QNode_Int_r,
          t2a8p_destruct_r,
          lizzieLet5_4QNode_Int_9QNode_Int_r,
          t3a8q_destruct_r} = {8 {(lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_r && lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_d[0])}};
  
  /* buf (Ty CT$wmAdd_Int) : (lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3,CT$wmAdd_Int) > (lizzieLet12_1_argbuf,CT$wmAdd_Int) */
  CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d;
  logic lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_r;
  assign lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_r = ((! lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d[0]) || lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d <= {115'd0,
                                                                                                                                                                                                                                     1'd0};
    else
      if (lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_r)
        lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d <= lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_d;
  CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf;
  assign lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_r = (! lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf[0] ? lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf :
                                   lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                       1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                         1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_buf <= lizzieLet5_4QNode_Int_4QNode_Int_1lizzieLet5_4QNode_Int_6QNode_Int_1lizzieLet5_4QNode_Int_7QNode_Int_1t1a8o_1lizzieLet5_4QNode_Int_8QNode_Int_1t2a8p_1lizzieLet5_4QNode_Int_9QNode_Int_1t3a8q_1Lcall_$wmAdd_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QNode_Int_4QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_4QNone_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_4QNone_Int_r = ((! lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QNode_Int_4QNone_Int_r)
        lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d <= lizzieLet5_4QNode_Int_4QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_4QNone_Int_bufchan_r = (! lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf :
                                                        lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_r && lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QNode_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_4QNone_Int_bufchan_buf <= lizzieLet5_4QNode_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QNode_Int_4QVal_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_4QVal_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_4QVal_Int_r = ((! lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QNode_Int_4QVal_Int_r)
        lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d <= lizzieLet5_4QNode_Int_4QVal_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_4QVal_Int_bufchan_r = (! lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf :
                                                       lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_r && lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QNode_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_4QVal_Int_bufchan_buf <= lizzieLet5_4QNode_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_5,QTree_Int) (lizzieLet5_6QNode_Int,Pointer_QTree_Int) > [(lizzieLet5_4QNode_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                                (_33,Pointer_QTree_Int),
                                                                                                                (_32,Pointer_QTree_Int),
                                                                                                                (_31,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet5_6QNode_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_5_d[0] && lizzieLet5_6QNode_Int_d[0]))
      unique case (lizzieLet5_4QNode_Int_5_d[2:1])
        2'd0: lizzieLet5_6QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_6QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_6QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_6QNode_Int_onehotd = 4'd8;
        default: lizzieLet5_6QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_6QNode_Int_onehotd = 4'd0;
  assign lizzieLet5_4QNode_Int_5QNone_Int_d = {lizzieLet5_6QNode_Int_d[16:1],
                                               lizzieLet5_6QNode_Int_onehotd[0]};
  assign _33_d = {lizzieLet5_6QNode_Int_d[16:1],
                  lizzieLet5_6QNode_Int_onehotd[1]};
  assign _32_d = {lizzieLet5_6QNode_Int_d[16:1],
                  lizzieLet5_6QNode_Int_onehotd[2]};
  assign _31_d = {lizzieLet5_6QNode_Int_d[16:1],
                  lizzieLet5_6QNode_Int_onehotd[3]};
  assign lizzieLet5_6QNode_Int_r = (| (lizzieLet5_6QNode_Int_onehotd & {_31_r,
                                                                        _32_r,
                                                                        _33_r,
                                                                        lizzieLet5_4QNode_Int_5QNone_Int_r}));
  assign lizzieLet5_4QNode_Int_5_r = lizzieLet5_6QNode_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d;
  logic lizzieLet5_4QNode_Int_5QNone_Int_bufchan_r;
  assign lizzieLet5_4QNode_Int_5QNone_Int_r = ((! lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d[0]) || lizzieLet5_4QNode_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QNode_Int_5QNone_Int_r)
        lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d <= lizzieLet5_4QNode_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet5_4QNode_Int_5QNone_Int_bufchan_r = (! lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_d = (lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf :
                                                        lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_r && lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QNode_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_5QNone_Int_bufchan_buf <= lizzieLet5_4QNode_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet5_4QNode_Int_6,QTree_Int) (lizzieLet5_8QNode_Int,MyDTInt_Int_Int) > [(_30,MyDTInt_Int_Int),
                                                                                                            (_29,MyDTInt_Int_Int),
                                                                                                            (lizzieLet5_4QNode_Int_6QNode_Int,MyDTInt_Int_Int),
                                                                                                            (_28,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet5_8QNode_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_6_d[0] && lizzieLet5_8QNode_Int_d[0]))
      unique case (lizzieLet5_4QNode_Int_6_d[2:1])
        2'd0: lizzieLet5_8QNode_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_8QNode_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_8QNode_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_8QNode_Int_onehotd = 4'd8;
        default: lizzieLet5_8QNode_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_8QNode_Int_onehotd = 4'd0;
  assign _30_d = lizzieLet5_8QNode_Int_onehotd[0];
  assign _29_d = lizzieLet5_8QNode_Int_onehotd[1];
  assign lizzieLet5_4QNode_Int_6QNode_Int_d = lizzieLet5_8QNode_Int_onehotd[2];
  assign _28_d = lizzieLet5_8QNode_Int_onehotd[3];
  assign lizzieLet5_8QNode_Int_r = (| (lizzieLet5_8QNode_Int_onehotd & {_28_r,
                                                                        lizzieLet5_4QNode_Int_6QNode_Int_r,
                                                                        _29_r,
                                                                        _30_r}));
  assign lizzieLet5_4QNode_Int_6_r = lizzieLet5_8QNode_Int_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet5_4QNode_Int_6QNode_Int,MyDTInt_Int_Int) > [(lizzieLet5_4QNode_Int_6QNode_Int_1,MyDTInt_Int_Int),
                                                                                  (lizzieLet5_4QNode_Int_6QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet5_4QNode_Int_6QNode_Int_emitted;
  logic [1:0] lizzieLet5_4QNode_Int_6QNode_Int_done;
  assign lizzieLet5_4QNode_Int_6QNode_Int_1_d = (lizzieLet5_4QNode_Int_6QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_6QNode_Int_emitted[0]));
  assign lizzieLet5_4QNode_Int_6QNode_Int_2_d = (lizzieLet5_4QNode_Int_6QNode_Int_d[0] && (! lizzieLet5_4QNode_Int_6QNode_Int_emitted[1]));
  assign lizzieLet5_4QNode_Int_6QNode_Int_done = (lizzieLet5_4QNode_Int_6QNode_Int_emitted | ({lizzieLet5_4QNode_Int_6QNode_Int_2_d[0],
                                                                                               lizzieLet5_4QNode_Int_6QNode_Int_1_d[0]} & {lizzieLet5_4QNode_Int_6QNode_Int_2_r,
                                                                                                                                           lizzieLet5_4QNode_Int_6QNode_Int_1_r}));
  assign lizzieLet5_4QNode_Int_6QNode_Int_r = (& lizzieLet5_4QNode_Int_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet5_4QNode_Int_6QNode_Int_emitted <= (lizzieLet5_4QNode_Int_6QNode_Int_r ? 2'd0 :
                                                   lizzieLet5_4QNode_Int_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet5_4QNode_Int_6QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d;
  logic lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_r;
  assign lizzieLet5_4QNode_Int_6QNode_Int_2_r = ((! lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d[0]) || lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QNode_Int_6QNode_Int_2_r)
        lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d <= lizzieLet5_4QNode_Int_6QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf;
  assign lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_r = (! lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_d = (lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf[0] ? lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf :
                                                        lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_r && lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QNode_Int_6QNode_Int_2_argbuf_r) && (! lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_buf <= lizzieLet5_4QNode_Int_6QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_7,QTree_Int) (q1a8j_destruct,Pointer_QTree_Int) > [(_27,Pointer_QTree_Int),
                                                                                                         (_26,Pointer_QTree_Int),
                                                                                                         (lizzieLet5_4QNode_Int_7QNode_Int,Pointer_QTree_Int),
                                                                                                         (_25,Pointer_QTree_Int)] */
  logic [3:0] q1a8j_destruct_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_7_d[0] && q1a8j_destruct_d[0]))
      unique case (lizzieLet5_4QNode_Int_7_d[2:1])
        2'd0: q1a8j_destruct_onehotd = 4'd1;
        2'd1: q1a8j_destruct_onehotd = 4'd2;
        2'd2: q1a8j_destruct_onehotd = 4'd4;
        2'd3: q1a8j_destruct_onehotd = 4'd8;
        default: q1a8j_destruct_onehotd = 4'd0;
      endcase
    else q1a8j_destruct_onehotd = 4'd0;
  assign _27_d = {q1a8j_destruct_d[16:1], q1a8j_destruct_onehotd[0]};
  assign _26_d = {q1a8j_destruct_d[16:1], q1a8j_destruct_onehotd[1]};
  assign lizzieLet5_4QNode_Int_7QNode_Int_d = {q1a8j_destruct_d[16:1],
                                               q1a8j_destruct_onehotd[2]};
  assign _25_d = {q1a8j_destruct_d[16:1], q1a8j_destruct_onehotd[3]};
  assign q1a8j_destruct_r = (| (q1a8j_destruct_onehotd & {_25_r,
                                                          lizzieLet5_4QNode_Int_7QNode_Int_r,
                                                          _26_r,
                                                          _27_r}));
  assign lizzieLet5_4QNode_Int_7_r = q1a8j_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_8,QTree_Int) (q2a8k_destruct,Pointer_QTree_Int) > [(_24,Pointer_QTree_Int),
                                                                                                         (_23,Pointer_QTree_Int),
                                                                                                         (lizzieLet5_4QNode_Int_8QNode_Int,Pointer_QTree_Int),
                                                                                                         (_22,Pointer_QTree_Int)] */
  logic [3:0] q2a8k_destruct_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_8_d[0] && q2a8k_destruct_d[0]))
      unique case (lizzieLet5_4QNode_Int_8_d[2:1])
        2'd0: q2a8k_destruct_onehotd = 4'd1;
        2'd1: q2a8k_destruct_onehotd = 4'd2;
        2'd2: q2a8k_destruct_onehotd = 4'd4;
        2'd3: q2a8k_destruct_onehotd = 4'd8;
        default: q2a8k_destruct_onehotd = 4'd0;
      endcase
    else q2a8k_destruct_onehotd = 4'd0;
  assign _24_d = {q2a8k_destruct_d[16:1], q2a8k_destruct_onehotd[0]};
  assign _23_d = {q2a8k_destruct_d[16:1], q2a8k_destruct_onehotd[1]};
  assign lizzieLet5_4QNode_Int_8QNode_Int_d = {q2a8k_destruct_d[16:1],
                                               q2a8k_destruct_onehotd[2]};
  assign _22_d = {q2a8k_destruct_d[16:1], q2a8k_destruct_onehotd[3]};
  assign q2a8k_destruct_r = (| (q2a8k_destruct_onehotd & {_22_r,
                                                          lizzieLet5_4QNode_Int_8QNode_Int_r,
                                                          _23_r,
                                                          _24_r}));
  assign lizzieLet5_4QNode_Int_8_r = q2a8k_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QNode_Int_9,QTree_Int) (q3a8l_destruct,Pointer_QTree_Int) > [(_21,Pointer_QTree_Int),
                                                                                                         (_20,Pointer_QTree_Int),
                                                                                                         (lizzieLet5_4QNode_Int_9QNode_Int,Pointer_QTree_Int),
                                                                                                         (_19,Pointer_QTree_Int)] */
  logic [3:0] q3a8l_destruct_onehotd;
  always_comb
    if ((lizzieLet5_4QNode_Int_9_d[0] && q3a8l_destruct_d[0]))
      unique case (lizzieLet5_4QNode_Int_9_d[2:1])
        2'd0: q3a8l_destruct_onehotd = 4'd1;
        2'd1: q3a8l_destruct_onehotd = 4'd2;
        2'd2: q3a8l_destruct_onehotd = 4'd4;
        2'd3: q3a8l_destruct_onehotd = 4'd8;
        default: q3a8l_destruct_onehotd = 4'd0;
      endcase
    else q3a8l_destruct_onehotd = 4'd0;
  assign _21_d = {q3a8l_destruct_d[16:1], q3a8l_destruct_onehotd[0]};
  assign _20_d = {q3a8l_destruct_d[16:1], q3a8l_destruct_onehotd[1]};
  assign lizzieLet5_4QNode_Int_9QNode_Int_d = {q3a8l_destruct_d[16:1],
                                               q3a8l_destruct_onehotd[2]};
  assign _19_d = {q3a8l_destruct_d[16:1], q3a8l_destruct_onehotd[3]};
  assign q3a8l_destruct_r = (| (q3a8l_destruct_onehotd & {_19_r,
                                                          lizzieLet5_4QNode_Int_9QNode_Int_r,
                                                          _20_r,
                                                          _21_r}));
  assign lizzieLet5_4QNode_Int_9_r = q3a8l_destruct_r;
  
  /* fork (Ty QTree_Int) : (lizzieLet5_4QVal_Int,QTree_Int) > [(lizzieLet5_4QVal_Int_1,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_2,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_3,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_4,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_5,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_6,QTree_Int),
                                                          (lizzieLet5_4QVal_Int_7,QTree_Int)] */
  logic [6:0] lizzieLet5_4QVal_Int_emitted;
  logic [6:0] lizzieLet5_4QVal_Int_done;
  assign lizzieLet5_4QVal_Int_1_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[0]))};
  assign lizzieLet5_4QVal_Int_2_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[1]))};
  assign lizzieLet5_4QVal_Int_3_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[2]))};
  assign lizzieLet5_4QVal_Int_4_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[3]))};
  assign lizzieLet5_4QVal_Int_5_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[4]))};
  assign lizzieLet5_4QVal_Int_6_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[5]))};
  assign lizzieLet5_4QVal_Int_7_d = {lizzieLet5_4QVal_Int_d[66:1],
                                     (lizzieLet5_4QVal_Int_d[0] && (! lizzieLet5_4QVal_Int_emitted[6]))};
  assign lizzieLet5_4QVal_Int_done = (lizzieLet5_4QVal_Int_emitted | ({lizzieLet5_4QVal_Int_7_d[0],
                                                                       lizzieLet5_4QVal_Int_6_d[0],
                                                                       lizzieLet5_4QVal_Int_5_d[0],
                                                                       lizzieLet5_4QVal_Int_4_d[0],
                                                                       lizzieLet5_4QVal_Int_3_d[0],
                                                                       lizzieLet5_4QVal_Int_2_d[0],
                                                                       lizzieLet5_4QVal_Int_1_d[0]} & {lizzieLet5_4QVal_Int_7_r,
                                                                                                       lizzieLet5_4QVal_Int_6_r,
                                                                                                       lizzieLet5_4QVal_Int_5_r,
                                                                                                       lizzieLet5_4QVal_Int_4_r,
                                                                                                       lizzieLet5_4QVal_Int_3_r,
                                                                                                       lizzieLet5_4QVal_Int_2_r,
                                                                                                       lizzieLet5_4QVal_Int_1_r}));
  assign lizzieLet5_4QVal_Int_r = (& lizzieLet5_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet5_4QVal_Int_emitted <= 7'd0;
    else
      lizzieLet5_4QVal_Int_emitted <= (lizzieLet5_4QVal_Int_r ? 7'd0 :
                                       lizzieLet5_4QVal_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet5_4QVal_Int_1QVal_Int,QTree_Int) > [(va8e_destruct,Int)] */
  assign va8e_destruct_d = {lizzieLet5_4QVal_Int_1QVal_Int_d[34:3],
                            lizzieLet5_4QVal_Int_1QVal_Int_d[0]};
  assign lizzieLet5_4QVal_Int_1QVal_Int_r = va8e_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet5_4QVal_Int_2,QTree_Int) (lizzieLet5_4QVal_Int_1,QTree_Int) > [(_18,QTree_Int),
                                                                                                (lizzieLet5_4QVal_Int_1QVal_Int,QTree_Int),
                                                                                                (_17,QTree_Int),
                                                                                                (_16,QTree_Int)] */
  logic [3:0] lizzieLet5_4QVal_Int_1_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_2_d[0] && lizzieLet5_4QVal_Int_1_d[0]))
      unique case (lizzieLet5_4QVal_Int_2_d[2:1])
        2'd0: lizzieLet5_4QVal_Int_1_onehotd = 4'd1;
        2'd1: lizzieLet5_4QVal_Int_1_onehotd = 4'd2;
        2'd2: lizzieLet5_4QVal_Int_1_onehotd = 4'd4;
        2'd3: lizzieLet5_4QVal_Int_1_onehotd = 4'd8;
        default: lizzieLet5_4QVal_Int_1_onehotd = 4'd0;
      endcase
    else lizzieLet5_4QVal_Int_1_onehotd = 4'd0;
  assign _18_d = {lizzieLet5_4QVal_Int_1_d[66:1],
                  lizzieLet5_4QVal_Int_1_onehotd[0]};
  assign lizzieLet5_4QVal_Int_1QVal_Int_d = {lizzieLet5_4QVal_Int_1_d[66:1],
                                             lizzieLet5_4QVal_Int_1_onehotd[1]};
  assign _17_d = {lizzieLet5_4QVal_Int_1_d[66:1],
                  lizzieLet5_4QVal_Int_1_onehotd[2]};
  assign _16_d = {lizzieLet5_4QVal_Int_1_d[66:1],
                  lizzieLet5_4QVal_Int_1_onehotd[3]};
  assign lizzieLet5_4QVal_Int_1_r = (| (lizzieLet5_4QVal_Int_1_onehotd & {_16_r,
                                                                          _17_r,
                                                                          lizzieLet5_4QVal_Int_1QVal_Int_r,
                                                                          _18_r}));
  assign lizzieLet5_4QVal_Int_2_r = lizzieLet5_4QVal_Int_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet5_4QVal_Int_3,QTree_Int) (lizzieLet5_3QVal_Int,Go) > [(lizzieLet5_4QVal_Int_3QNone_Int,Go),
                                                                                (lizzieLet5_4QVal_Int_3QVal_Int,Go),
                                                                                (lizzieLet5_4QVal_Int_3QNode_Int,Go),
                                                                                (lizzieLet5_4QVal_Int_3QError_Int,Go)] */
  logic [3:0] lizzieLet5_3QVal_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_3_d[0] && lizzieLet5_3QVal_Int_d[0]))
      unique case (lizzieLet5_4QVal_Int_3_d[2:1])
        2'd0: lizzieLet5_3QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_3QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_3QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_3QVal_Int_onehotd = 4'd8;
        default: lizzieLet5_3QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_3QVal_Int_onehotd = 4'd0;
  assign lizzieLet5_4QVal_Int_3QNone_Int_d = lizzieLet5_3QVal_Int_onehotd[0];
  assign lizzieLet5_4QVal_Int_3QVal_Int_d = lizzieLet5_3QVal_Int_onehotd[1];
  assign lizzieLet5_4QVal_Int_3QNode_Int_d = lizzieLet5_3QVal_Int_onehotd[2];
  assign lizzieLet5_4QVal_Int_3QError_Int_d = lizzieLet5_3QVal_Int_onehotd[3];
  assign lizzieLet5_3QVal_Int_r = (| (lizzieLet5_3QVal_Int_onehotd & {lizzieLet5_4QVal_Int_3QError_Int_r,
                                                                      lizzieLet5_4QVal_Int_3QNode_Int_r,
                                                                      lizzieLet5_4QVal_Int_3QVal_Int_r,
                                                                      lizzieLet5_4QVal_Int_3QNone_Int_r}));
  assign lizzieLet5_4QVal_Int_3_r = lizzieLet5_3QVal_Int_r;
  
  /* fork (Ty Go) : (lizzieLet5_4QVal_Int_3QError_Int,Go) > [(lizzieLet5_4QVal_Int_3QError_Int_1,Go),
                                                        (lizzieLet5_4QVal_Int_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet5_4QVal_Int_3QError_Int_emitted;
  logic [1:0] lizzieLet5_4QVal_Int_3QError_Int_done;
  assign lizzieLet5_4QVal_Int_3QError_Int_1_d = (lizzieLet5_4QVal_Int_3QError_Int_d[0] && (! lizzieLet5_4QVal_Int_3QError_Int_emitted[0]));
  assign lizzieLet5_4QVal_Int_3QError_Int_2_d = (lizzieLet5_4QVal_Int_3QError_Int_d[0] && (! lizzieLet5_4QVal_Int_3QError_Int_emitted[1]));
  assign lizzieLet5_4QVal_Int_3QError_Int_done = (lizzieLet5_4QVal_Int_3QError_Int_emitted | ({lizzieLet5_4QVal_Int_3QError_Int_2_d[0],
                                                                                               lizzieLet5_4QVal_Int_3QError_Int_1_d[0]} & {lizzieLet5_4QVal_Int_3QError_Int_2_r,
                                                                                                                                           lizzieLet5_4QVal_Int_3QError_Int_1_r}));
  assign lizzieLet5_4QVal_Int_3QError_Int_r = (& lizzieLet5_4QVal_Int_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet5_4QVal_Int_3QError_Int_emitted <= (lizzieLet5_4QVal_Int_3QError_Int_r ? 2'd0 :
                                                   lizzieLet5_4QVal_Int_3QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet5_4QVal_Int_3QError_Int_1,Go)] > (lizzieLet5_4QVal_Int_3QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet5_4QVal_Int_3QError_Int_1_d[0]}), lizzieLet5_4QVal_Int_3QError_Int_1_d);
  assign {lizzieLet5_4QVal_Int_3QError_Int_1_r} = {1 {(lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_r && lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet5_4QVal_Int_3QError_Int_1QError_Int,QTree_Int) > (lizzieLet9_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_r = ((! lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                 1'd0};
    else
      if (lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_r)
        lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d <= lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_r = (! lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf :
                                    lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                   1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                     1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_buf <= lizzieLet5_4QVal_Int_3QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QVal_Int_3QError_Int_2,Go) > (lizzieLet5_4QVal_Int_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QError_Int_2_r = ((! lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QVal_Int_3QError_Int_2_r)
        lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d <= lizzieLet5_4QVal_Int_3QError_Int_2_d;
  Go_t lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_r = (! lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_d = (lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf :
                                                        lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_r && lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QVal_Int_3QError_Int_2_argbuf_r) && (! lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_buf <= lizzieLet5_4QVal_Int_3QError_Int_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet5_4QVal_Int_3QNode_Int,Go) > [(lizzieLet5_4QVal_Int_3QNode_Int_1,Go),
                                                       (lizzieLet5_4QVal_Int_3QNode_Int_2,Go)] */
  logic [1:0] lizzieLet5_4QVal_Int_3QNode_Int_emitted;
  logic [1:0] lizzieLet5_4QVal_Int_3QNode_Int_done;
  assign lizzieLet5_4QVal_Int_3QNode_Int_1_d = (lizzieLet5_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet5_4QVal_Int_3QNode_Int_emitted[0]));
  assign lizzieLet5_4QVal_Int_3QNode_Int_2_d = (lizzieLet5_4QVal_Int_3QNode_Int_d[0] && (! lizzieLet5_4QVal_Int_3QNode_Int_emitted[1]));
  assign lizzieLet5_4QVal_Int_3QNode_Int_done = (lizzieLet5_4QVal_Int_3QNode_Int_emitted | ({lizzieLet5_4QVal_Int_3QNode_Int_2_d[0],
                                                                                             lizzieLet5_4QVal_Int_3QNode_Int_1_d[0]} & {lizzieLet5_4QVal_Int_3QNode_Int_2_r,
                                                                                                                                        lizzieLet5_4QVal_Int_3QNode_Int_1_r}));
  assign lizzieLet5_4QVal_Int_3QNode_Int_r = (& lizzieLet5_4QVal_Int_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet5_4QVal_Int_3QNode_Int_emitted <= (lizzieLet5_4QVal_Int_3QNode_Int_r ? 2'd0 :
                                                  lizzieLet5_4QVal_Int_3QNode_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet5_4QVal_Int_3QNode_Int_1,Go)] > (lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int,QTree_Int) */
  assign lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet5_4QVal_Int_3QNode_Int_1_d[0]}), lizzieLet5_4QVal_Int_3QNode_Int_1_d);
  assign {lizzieLet5_4QVal_Int_3QNode_Int_1_r} = {1 {(lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_r && lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int,QTree_Int) > (lizzieLet8_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_r = ((! lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= {66'd0,
                                                                1'd0};
    else
      if (lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_r)
        lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d <= lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_d;
  QTree_Int_t lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_r = (! lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf :
                                    lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                  1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= {66'd0,
                                                                    1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_buf <= lizzieLet5_4QVal_Int_3QNode_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QVal_Int_3QNode_Int_2,Go) > (lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf,Go) */
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QNode_Int_2_r = ((! lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QVal_Int_3QNode_Int_2_r)
        lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d <= lizzieLet5_4QVal_Int_3QNode_Int_2_d;
  Go_t lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_r = (! lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_d = (lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf :
                                                       lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_r && lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QVal_Int_3QNode_Int_2_argbuf_r) && (! lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_buf <= lizzieLet5_4QVal_Int_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QVal_Int_3QNone_Int,Go) > (lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QNone_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QNone_Int_r = ((! lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QVal_Int_3QNone_Int_r)
        lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d <= lizzieLet5_4QVal_Int_3QNone_Int_d;
  Go_t lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QNone_Int_bufchan_r = (! lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf :
                                                       lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_r && lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QVal_Int_3QNone_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QNone_Int_bufchan_buf <= lizzieLet5_4QVal_Int_3QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet5_4QVal_Int_3QVal_Int,Go) > (lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_3QVal_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_3QVal_Int_r = ((! lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QVal_Int_3QVal_Int_r)
        lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d <= lizzieLet5_4QVal_Int_3QVal_Int_d;
  Go_t lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_3QVal_Int_bufchan_r = (! lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf :
                                                      lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_r && lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QVal_Int_3QVal_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_3QVal_Int_bufchan_buf <= lizzieLet5_4QVal_Int_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QVal_Int_4,QTree_Int) (lizzieLet5_5QVal_Int,Pointer_CT$wmAdd_Int) > [(lizzieLet5_4QVal_Int_4QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet5_4QVal_Int_4QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet5_4QVal_Int_4QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                                    (lizzieLet5_4QVal_Int_4QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] lizzieLet5_5QVal_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_4_d[0] && lizzieLet5_5QVal_Int_d[0]))
      unique case (lizzieLet5_4QVal_Int_4_d[2:1])
        2'd0: lizzieLet5_5QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_5QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_5QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_5QVal_Int_onehotd = 4'd8;
        default: lizzieLet5_5QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_5QVal_Int_onehotd = 4'd0;
  assign lizzieLet5_4QVal_Int_4QNone_Int_d = {lizzieLet5_5QVal_Int_d[16:1],
                                              lizzieLet5_5QVal_Int_onehotd[0]};
  assign lizzieLet5_4QVal_Int_4QVal_Int_d = {lizzieLet5_5QVal_Int_d[16:1],
                                             lizzieLet5_5QVal_Int_onehotd[1]};
  assign lizzieLet5_4QVal_Int_4QNode_Int_d = {lizzieLet5_5QVal_Int_d[16:1],
                                              lizzieLet5_5QVal_Int_onehotd[2]};
  assign lizzieLet5_4QVal_Int_4QError_Int_d = {lizzieLet5_5QVal_Int_d[16:1],
                                               lizzieLet5_5QVal_Int_onehotd[3]};
  assign lizzieLet5_5QVal_Int_r = (| (lizzieLet5_5QVal_Int_onehotd & {lizzieLet5_4QVal_Int_4QError_Int_r,
                                                                      lizzieLet5_4QVal_Int_4QNode_Int_r,
                                                                      lizzieLet5_4QVal_Int_4QVal_Int_r,
                                                                      lizzieLet5_4QVal_Int_4QNone_Int_r}));
  assign lizzieLet5_4QVal_Int_4_r = lizzieLet5_5QVal_Int_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QVal_Int_4QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QVal_Int_4QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QError_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_4QError_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_4QError_Int_r = ((! lizzieLet5_4QVal_Int_4QError_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_4QError_Int_r)
        lizzieLet5_4QVal_Int_4QError_Int_bufchan_d <= lizzieLet5_4QVal_Int_4QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_4QError_Int_bufchan_r = (! lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf :
                                                        lizzieLet5_4QVal_Int_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_r && lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_4QError_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_4QError_Int_bufchan_buf <= lizzieLet5_4QVal_Int_4QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QVal_Int_4QNode_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_4QNode_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_4QNode_Int_r = ((! lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_4QNode_Int_r)
        lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d <= lizzieLet5_4QVal_Int_4QNode_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_4QNode_Int_bufchan_r = (! lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf :
                                                       lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_r && lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_4QNode_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_4QNode_Int_bufchan_buf <= lizzieLet5_4QVal_Int_4QNode_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QVal_Int_4QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_4QNone_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_4QNone_Int_r = ((! lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_4QNone_Int_r)
        lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d <= lizzieLet5_4QVal_Int_4QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_4QNone_Int_bufchan_r = (! lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf :
                                                       lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_r && lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_4QNone_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_4QNone_Int_bufchan_buf <= lizzieLet5_4QVal_Int_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_4QVal_Int_4QVal_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_4QVal_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_4QVal_Int_r = ((! lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_4QVal_Int_r)
        lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d <= lizzieLet5_4QVal_Int_4QVal_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_4QVal_Int_bufchan_r = (! lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf :
                                                      lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_r && lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_4QVal_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_4QVal_Int_bufchan_buf <= lizzieLet5_4QVal_Int_4QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_4QVal_Int_5,QTree_Int) (lizzieLet5_6QVal_Int,Pointer_QTree_Int) > [(lizzieLet5_4QVal_Int_5QNone_Int,Pointer_QTree_Int),
                                                                                                              (_15,Pointer_QTree_Int),
                                                                                                              (_14,Pointer_QTree_Int),
                                                                                                              (_13,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet5_6QVal_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_5_d[0] && lizzieLet5_6QVal_Int_d[0]))
      unique case (lizzieLet5_4QVal_Int_5_d[2:1])
        2'd0: lizzieLet5_6QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_6QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_6QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_6QVal_Int_onehotd = 4'd8;
        default: lizzieLet5_6QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_6QVal_Int_onehotd = 4'd0;
  assign lizzieLet5_4QVal_Int_5QNone_Int_d = {lizzieLet5_6QVal_Int_d[16:1],
                                              lizzieLet5_6QVal_Int_onehotd[0]};
  assign _15_d = {lizzieLet5_6QVal_Int_d[16:1],
                  lizzieLet5_6QVal_Int_onehotd[1]};
  assign _14_d = {lizzieLet5_6QVal_Int_d[16:1],
                  lizzieLet5_6QVal_Int_onehotd[2]};
  assign _13_d = {lizzieLet5_6QVal_Int_d[16:1],
                  lizzieLet5_6QVal_Int_onehotd[3]};
  assign lizzieLet5_6QVal_Int_r = (| (lizzieLet5_6QVal_Int_onehotd & {_13_r,
                                                                      _14_r,
                                                                      _15_r,
                                                                      lizzieLet5_4QVal_Int_5QNone_Int_r}));
  assign lizzieLet5_4QVal_Int_5_r = lizzieLet5_6QVal_Int_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet5_4QVal_Int_5QNone_Int,Pointer_QTree_Int) > (lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_5QNone_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_5QNone_Int_r = ((! lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_5QNone_Int_r)
        lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d <= lizzieLet5_4QVal_Int_5QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_5QNone_Int_bufchan_r = (! lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf :
                                                       lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_r && lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_5QNone_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_5QNone_Int_bufchan_buf <= lizzieLet5_4QVal_Int_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet5_4QVal_Int_6,QTree_Int) (lizzieLet5_8QVal_Int,MyDTInt_Int_Int) > [(_12,MyDTInt_Int_Int),
                                                                                                          (lizzieLet5_4QVal_Int_6QVal_Int,MyDTInt_Int_Int),
                                                                                                          (_11,MyDTInt_Int_Int),
                                                                                                          (_10,MyDTInt_Int_Int)] */
  logic [3:0] lizzieLet5_8QVal_Int_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_6_d[0] && lizzieLet5_8QVal_Int_d[0]))
      unique case (lizzieLet5_4QVal_Int_6_d[2:1])
        2'd0: lizzieLet5_8QVal_Int_onehotd = 4'd1;
        2'd1: lizzieLet5_8QVal_Int_onehotd = 4'd2;
        2'd2: lizzieLet5_8QVal_Int_onehotd = 4'd4;
        2'd3: lizzieLet5_8QVal_Int_onehotd = 4'd8;
        default: lizzieLet5_8QVal_Int_onehotd = 4'd0;
      endcase
    else lizzieLet5_8QVal_Int_onehotd = 4'd0;
  assign _12_d = lizzieLet5_8QVal_Int_onehotd[0];
  assign lizzieLet5_4QVal_Int_6QVal_Int_d = lizzieLet5_8QVal_Int_onehotd[1];
  assign _11_d = lizzieLet5_8QVal_Int_onehotd[2];
  assign _10_d = lizzieLet5_8QVal_Int_onehotd[3];
  assign lizzieLet5_8QVal_Int_r = (| (lizzieLet5_8QVal_Int_onehotd & {_10_r,
                                                                      _11_r,
                                                                      lizzieLet5_4QVal_Int_6QVal_Int_r,
                                                                      _12_r}));
  assign lizzieLet5_4QVal_Int_6_r = lizzieLet5_8QVal_Int_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet5_4QVal_Int_6QVal_Int,MyDTInt_Int_Int) > (lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_6QVal_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_6QVal_Int_r = ((! lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet5_4QVal_Int_6QVal_Int_r)
        lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d <= lizzieLet5_4QVal_Int_6QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_6QVal_Int_bufchan_r = (! lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf :
                                                      lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_r && lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_6QVal_Int_bufchan_buf <= lizzieLet5_4QVal_Int_6QVal_Int_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf,Int),
                                              (va8e_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_d[0],
                                                                                                        va8e_1_argbuf_d[0]}), lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_d, lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_d, va8e_1_argbuf_d);
  assign {lizzieLet5_4QVal_Int_6QVal_Int_1_argbuf_r,
          lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_r,
          va8e_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet5_4QVal_Int_7,QTree_Int) (v1a8d_destruct,Int) > [(_9,Int),
                                                                            (lizzieLet5_4QVal_Int_7QVal_Int,Int),
                                                                            (_8,Int),
                                                                            (_7,Int)] */
  logic [3:0] v1a8d_destruct_onehotd;
  always_comb
    if ((lizzieLet5_4QVal_Int_7_d[0] && v1a8d_destruct_d[0]))
      unique case (lizzieLet5_4QVal_Int_7_d[2:1])
        2'd0: v1a8d_destruct_onehotd = 4'd1;
        2'd1: v1a8d_destruct_onehotd = 4'd2;
        2'd2: v1a8d_destruct_onehotd = 4'd4;
        2'd3: v1a8d_destruct_onehotd = 4'd8;
        default: v1a8d_destruct_onehotd = 4'd0;
      endcase
    else v1a8d_destruct_onehotd = 4'd0;
  assign _9_d = {v1a8d_destruct_d[32:1], v1a8d_destruct_onehotd[0]};
  assign lizzieLet5_4QVal_Int_7QVal_Int_d = {v1a8d_destruct_d[32:1],
                                             v1a8d_destruct_onehotd[1]};
  assign _8_d = {v1a8d_destruct_d[32:1], v1a8d_destruct_onehotd[2]};
  assign _7_d = {v1a8d_destruct_d[32:1], v1a8d_destruct_onehotd[3]};
  assign v1a8d_destruct_r = (| (v1a8d_destruct_onehotd & {_7_r,
                                                          _8_r,
                                                          lizzieLet5_4QVal_Int_7QVal_Int_r,
                                                          _9_r}));
  assign lizzieLet5_4QVal_Int_7_r = v1a8d_destruct_r;
  
  /* buf (Ty Int) : (lizzieLet5_4QVal_Int_7QVal_Int,Int) > (lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d;
  logic lizzieLet5_4QVal_Int_7QVal_Int_bufchan_r;
  assign lizzieLet5_4QVal_Int_7QVal_Int_r = ((! lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d[0]) || lizzieLet5_4QVal_Int_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet5_4QVal_Int_7QVal_Int_r)
        lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d <= lizzieLet5_4QVal_Int_7QVal_Int_d;
  Int_t lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf;
  assign lizzieLet5_4QVal_Int_7QVal_Int_bufchan_r = (! lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_d = (lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf[0] ? lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf :
                                                      lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_r && lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf[0]))
        lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet5_4QVal_Int_7QVal_Int_1_argbuf_r) && (! lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf[0])))
        lizzieLet5_4QVal_Int_7QVal_Int_bufchan_buf <= lizzieLet5_4QVal_Int_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_5,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wmAdd_Int) > [(lizzieLet5_5QNone_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet5_5QVal_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet5_5QNode_Int,Pointer_CT$wmAdd_Int),
                                                                                                    (lizzieLet5_5QError_Int,Pointer_CT$wmAdd_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet5_5_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet5_5_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet5_5QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet5_5QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet5_5QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet5_5QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet5_5QError_Int_r,
                                                          lizzieLet5_5QNode_Int_r,
                                                          lizzieLet5_5QVal_Int_r,
                                                          lizzieLet5_5QNone_Int_r}));
  assign lizzieLet5_5_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_5QError_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_5QError_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QError_Int_bufchan_d;
  logic lizzieLet5_5QError_Int_bufchan_r;
  assign lizzieLet5_5QError_Int_r = ((! lizzieLet5_5QError_Int_bufchan_d[0]) || lizzieLet5_5QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_5QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_5QError_Int_r)
        lizzieLet5_5QError_Int_bufchan_d <= lizzieLet5_5QError_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QError_Int_bufchan_buf;
  assign lizzieLet5_5QError_Int_bufchan_r = (! lizzieLet5_5QError_Int_bufchan_buf[0]);
  assign lizzieLet5_5QError_Int_1_argbuf_d = (lizzieLet5_5QError_Int_bufchan_buf[0] ? lizzieLet5_5QError_Int_bufchan_buf :
                                              lizzieLet5_5QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_5QError_Int_1_argbuf_r && lizzieLet5_5QError_Int_bufchan_buf[0]))
        lizzieLet5_5QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_5QError_Int_1_argbuf_r) && (! lizzieLet5_5QError_Int_bufchan_buf[0])))
        lizzieLet5_5QError_Int_bufchan_buf <= lizzieLet5_5QError_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (lizzieLet5_5QNone_Int,Pointer_CT$wmAdd_Int) > (lizzieLet5_5QNone_Int_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QNone_Int_bufchan_d;
  logic lizzieLet5_5QNone_Int_bufchan_r;
  assign lizzieLet5_5QNone_Int_r = ((! lizzieLet5_5QNone_Int_bufchan_d[0]) || lizzieLet5_5QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_5QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_5QNone_Int_r)
        lizzieLet5_5QNone_Int_bufchan_d <= lizzieLet5_5QNone_Int_d;
  Pointer_CT$wmAdd_Int_t lizzieLet5_5QNone_Int_bufchan_buf;
  assign lizzieLet5_5QNone_Int_bufchan_r = (! lizzieLet5_5QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_5QNone_Int_1_argbuf_d = (lizzieLet5_5QNone_Int_bufchan_buf[0] ? lizzieLet5_5QNone_Int_bufchan_buf :
                                             lizzieLet5_5QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_5QNone_Int_1_argbuf_r && lizzieLet5_5QNone_Int_bufchan_buf[0]))
        lizzieLet5_5QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_5QNone_Int_1_argbuf_r) && (! lizzieLet5_5QNone_Int_bufchan_buf[0])))
        lizzieLet5_5QNone_Int_bufchan_buf <= lizzieLet5_5QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_6,QTree_Int) (w1slS_1_2,Pointer_QTree_Int) > [(_6,Pointer_QTree_Int),
                                                                                         (lizzieLet5_6QVal_Int,Pointer_QTree_Int),
                                                                                         (lizzieLet5_6QNode_Int,Pointer_QTree_Int),
                                                                                         (_5,Pointer_QTree_Int)] */
  logic [3:0] w1slS_1_2_onehotd;
  always_comb
    if ((lizzieLet5_6_d[0] && w1slS_1_2_d[0]))
      unique case (lizzieLet5_6_d[2:1])
        2'd0: w1slS_1_2_onehotd = 4'd1;
        2'd1: w1slS_1_2_onehotd = 4'd2;
        2'd2: w1slS_1_2_onehotd = 4'd4;
        2'd3: w1slS_1_2_onehotd = 4'd8;
        default: w1slS_1_2_onehotd = 4'd0;
      endcase
    else w1slS_1_2_onehotd = 4'd0;
  assign _6_d = {w1slS_1_2_d[16:1], w1slS_1_2_onehotd[0]};
  assign lizzieLet5_6QVal_Int_d = {w1slS_1_2_d[16:1],
                                   w1slS_1_2_onehotd[1]};
  assign lizzieLet5_6QNode_Int_d = {w1slS_1_2_d[16:1],
                                    w1slS_1_2_onehotd[2]};
  assign _5_d = {w1slS_1_2_d[16:1], w1slS_1_2_onehotd[3]};
  assign w1slS_1_2_r = (| (w1slS_1_2_onehotd & {_5_r,
                                                lizzieLet5_6QNode_Int_r,
                                                lizzieLet5_6QVal_Int_r,
                                                _6_r}));
  assign lizzieLet5_6_r = w1slS_1_2_r;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet5_7,QTree_Int) (w2slT_1_2,Pointer_QTree_Int) > [(lizzieLet5_7QNone_Int,Pointer_QTree_Int),
                                                                                         (_4,Pointer_QTree_Int),
                                                                                         (_3,Pointer_QTree_Int),
                                                                                         (_2,Pointer_QTree_Int)] */
  logic [3:0] w2slT_1_2_onehotd;
  always_comb
    if ((lizzieLet5_7_d[0] && w2slT_1_2_d[0]))
      unique case (lizzieLet5_7_d[2:1])
        2'd0: w2slT_1_2_onehotd = 4'd1;
        2'd1: w2slT_1_2_onehotd = 4'd2;
        2'd2: w2slT_1_2_onehotd = 4'd4;
        2'd3: w2slT_1_2_onehotd = 4'd8;
        default: w2slT_1_2_onehotd = 4'd0;
      endcase
    else w2slT_1_2_onehotd = 4'd0;
  assign lizzieLet5_7QNone_Int_d = {w2slT_1_2_d[16:1],
                                    w2slT_1_2_onehotd[0]};
  assign _4_d = {w2slT_1_2_d[16:1], w2slT_1_2_onehotd[1]};
  assign _3_d = {w2slT_1_2_d[16:1], w2slT_1_2_onehotd[2]};
  assign _2_d = {w2slT_1_2_d[16:1], w2slT_1_2_onehotd[3]};
  assign w2slT_1_2_r = (| (w2slT_1_2_onehotd & {_2_r,
                                                _3_r,
                                                _4_r,
                                                lizzieLet5_7QNone_Int_r}));
  assign lizzieLet5_7_r = w2slT_1_2_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet5_7QNone_Int,Pointer_QTree_Int) > (lizzieLet5_7QNone_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet5_7QNone_Int_bufchan_d;
  logic lizzieLet5_7QNone_Int_bufchan_r;
  assign lizzieLet5_7QNone_Int_r = ((! lizzieLet5_7QNone_Int_bufchan_d[0]) || lizzieLet5_7QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_7QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet5_7QNone_Int_r)
        lizzieLet5_7QNone_Int_bufchan_d <= lizzieLet5_7QNone_Int_d;
  Pointer_QTree_Int_t lizzieLet5_7QNone_Int_bufchan_buf;
  assign lizzieLet5_7QNone_Int_bufchan_r = (! lizzieLet5_7QNone_Int_bufchan_buf[0]);
  assign lizzieLet5_7QNone_Int_1_argbuf_d = (lizzieLet5_7QNone_Int_bufchan_buf[0] ? lizzieLet5_7QNone_Int_bufchan_buf :
                                             lizzieLet5_7QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet5_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet5_7QNone_Int_1_argbuf_r && lizzieLet5_7QNone_Int_bufchan_buf[0]))
        lizzieLet5_7QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet5_7QNone_Int_1_argbuf_r) && (! lizzieLet5_7QNone_Int_bufchan_buf[0])))
        lizzieLet5_7QNone_Int_bufchan_buf <= lizzieLet5_7QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet5_8,QTree_Int) (wslR_1_goMux_mux,MyDTInt_Int_Int) > [(_1,MyDTInt_Int_Int),
                                                                                            (lizzieLet5_8QVal_Int,MyDTInt_Int_Int),
                                                                                            (lizzieLet5_8QNode_Int,MyDTInt_Int_Int),
                                                                                            (_0,MyDTInt_Int_Int)] */
  logic [3:0] wslR_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet5_8_d[0] && wslR_1_goMux_mux_d[0]))
      unique case (lizzieLet5_8_d[2:1])
        2'd0: wslR_1_goMux_mux_onehotd = 4'd1;
        2'd1: wslR_1_goMux_mux_onehotd = 4'd2;
        2'd2: wslR_1_goMux_mux_onehotd = 4'd4;
        2'd3: wslR_1_goMux_mux_onehotd = 4'd8;
        default: wslR_1_goMux_mux_onehotd = 4'd0;
      endcase
    else wslR_1_goMux_mux_onehotd = 4'd0;
  assign _1_d = wslR_1_goMux_mux_onehotd[0];
  assign lizzieLet5_8QVal_Int_d = wslR_1_goMux_mux_onehotd[1];
  assign lizzieLet5_8QNode_Int_d = wslR_1_goMux_mux_onehotd[2];
  assign _0_d = wslR_1_goMux_mux_onehotd[3];
  assign wslR_1_goMux_mux_r = (| (wslR_1_goMux_mux_onehotd & {_0_r,
                                                              lizzieLet5_8QNode_Int_r,
                                                              lizzieLet5_8QVal_Int_r,
                                                              _1_r}));
  assign lizzieLet5_8_r = wslR_1_goMux_mux_r;
  
  /* buf (Ty Pointer_QTree_Int) : (ma8M_goMux_mux,Pointer_QTree_Int) > (ma8M_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t ma8M_goMux_mux_bufchan_d;
  logic ma8M_goMux_mux_bufchan_r;
  assign ma8M_goMux_mux_r = ((! ma8M_goMux_mux_bufchan_d[0]) || ma8M_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8M_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (ma8M_goMux_mux_r) ma8M_goMux_mux_bufchan_d <= ma8M_goMux_mux_d;
  Pointer_QTree_Int_t ma8M_goMux_mux_bufchan_buf;
  assign ma8M_goMux_mux_bufchan_r = (! ma8M_goMux_mux_bufchan_buf[0]);
  assign ma8M_1_argbuf_d = (ma8M_goMux_mux_bufchan_buf[0] ? ma8M_goMux_mux_bufchan_buf :
                            ma8M_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8M_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((ma8M_1_argbuf_r && ma8M_goMux_mux_bufchan_buf[0]))
        ma8M_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! ma8M_1_argbuf_r) && (! ma8M_goMux_mux_bufchan_buf[0])))
        ma8M_goMux_mux_bufchan_buf <= ma8M_goMux_mux_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int,
          Dcon TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int) : (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1,TupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int) > [(main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14,Go),
                                                                                                                                                                                                                      (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1,MyDTBool_Bool),
                                                                                                                                                                                                                      (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1,MyDTInt_Bool),
                                                                                                                                                                                                                      (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1,Pointer_QTree_Int)] */
  logic [3:0] \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted ;
  logic [3:0] \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_done ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_d  = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted [0]));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_d  = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted [1]));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_d  = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted [2]));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_d  = {\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [16:1],
                                                                                                 (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted [3]))};
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_done  = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted  | ({\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_d [0],
                                                                                                                                                                                           \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_d [0],
                                                                                                                                                                                           \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_d [0],
                                                                                                                                                                                           \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_d [0]} & {\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_r }));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_r  = (& \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted  <= 4'd0;
    else
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_emitted  <= (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_r  ? 4'd0 :
                                                                                                 \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Int_1_done );
  
  /* buf (Ty MyDTInt_Bool) : (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1,MyDTInt_Bool) > (ga8L_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_r ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_r  = ((! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d [0]) || \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_r )
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_d ;
  MyDTInt_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_r  = (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf [0]);
  assign ga8L_1_1_argbuf_d = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf [0] ? \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf  :
                              \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf  <= 1'd0;
    else
      if ((ga8L_1_1_argbuf_r && \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf [0]))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf  <= 1'd0;
      else if (((! ga8L_1_1_argbuf_r) && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf [0])))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_buf  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intga8L_1_bufchan_d ;
  
  /* fork (Ty Go) : (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14,Go) > [(go_14_1,Go),
                                                                                                       (go_14_2,Go)] */
  logic [1:0] \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted ;
  logic [1:0] \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_done ;
  assign go_14_1_d = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted [0]));
  assign go_14_2_d = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_d [0] && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted [1]));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_done  = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted  | ({go_14_2_d[0],
                                                                                                                                                                                                 go_14_1_d[0]} & {go_14_2_r,
                                                                                                                                                                                                                  go_14_1_r}));
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_r  = (& \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted  <= 2'd0;
    else
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_emitted  <= (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_r  ? 2'd0 :
                                                                                                    \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intgo_14_done );
  
  /* buf (Ty MyDTBool_Bool) : (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1,MyDTBool_Bool) > (isZa8K_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_r ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_r  = ((! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d [0]) || \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_r )
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_d ;
  MyDTBool_Bool_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_r  = (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf [0]);
  assign isZa8K_1_1_argbuf_d = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf [0] ? \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf  :
                                \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf  <= 1'd0;
    else
      if ((isZa8K_1_1_argbuf_r && \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf [0]))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf  <= 1'd0;
      else if (((! isZa8K_1_1_argbuf_r) && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf [0])))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_buf  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_IntisZa8K_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1,Pointer_QTree_Int) > (ma8M_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d ;
  logic \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_r ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_r  = ((! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d [0]) || \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d  <= {16'd0,
                                                                                                       1'd0};
    else
      if (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_r )
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_d ;
  Pointer_QTree_Int_t \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf ;
  assign \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_r  = (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf [0]);
  assign ma8M_1_1_argbuf_d = (\main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf [0] ? \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf  :
                              \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
    else
      if ((ma8M_1_1_argbuf_r && \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf [0]))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf  <= {16'd0,
                                                                                                           1'd0};
      else if (((! ma8M_1_1_argbuf_r) && (! \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf [0])))
        \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_buf  <= \main_map'_Int_BoolTupGo___MyDTBool_Bool___MyDTInt_Bool___Pointer_QTree_Intma8M_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (main_map'_Int_Bool_resbuf,Pointer_QTree_Bool) > (es_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \main_map'_Int_Bool_resbuf_bufchan_d ;
  logic \main_map'_Int_Bool_resbuf_bufchan_r ;
  assign \main_map'_Int_Bool_resbuf_r  = ((! \main_map'_Int_Bool_resbuf_bufchan_d [0]) || \main_map'_Int_Bool_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_Bool_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\main_map'_Int_Bool_resbuf_r )
        \main_map'_Int_Bool_resbuf_bufchan_d  <= \main_map'_Int_Bool_resbuf_d ;
  Pointer_QTree_Bool_t \main_map'_Int_Bool_resbuf_bufchan_buf ;
  assign \main_map'_Int_Bool_resbuf_bufchan_r  = (! \main_map'_Int_Bool_resbuf_bufchan_buf [0]);
  assign es_0_1_1_argbuf_d = (\main_map'_Int_Bool_resbuf_bufchan_buf [0] ? \main_map'_Int_Bool_resbuf_bufchan_buf  :
                              \main_map'_Int_Bool_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Int_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((es_0_1_1_argbuf_r && \main_map'_Int_Bool_resbuf_bufchan_buf [0]))
        \main_map'_Int_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! es_0_1_1_argbuf_r) && (! \main_map'_Int_Bool_resbuf_bufchan_buf [0])))
        \main_map'_Int_Bool_resbuf_bufchan_buf  <= \main_map'_Int_Bool_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8O_3_destruct,Pointer_QTree_Int) > (q1a8O_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8O_3_destruct_bufchan_d;
  logic q1a8O_3_destruct_bufchan_r;
  assign q1a8O_3_destruct_r = ((! q1a8O_3_destruct_bufchan_d[0]) || q1a8O_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8O_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8O_3_destruct_r)
        q1a8O_3_destruct_bufchan_d <= q1a8O_3_destruct_d;
  Pointer_QTree_Int_t q1a8O_3_destruct_bufchan_buf;
  assign q1a8O_3_destruct_bufchan_r = (! q1a8O_3_destruct_bufchan_buf[0]);
  assign q1a8O_3_1_argbuf_d = (q1a8O_3_destruct_bufchan_buf[0] ? q1a8O_3_destruct_bufchan_buf :
                               q1a8O_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8O_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8O_3_1_argbuf_r && q1a8O_3_destruct_bufchan_buf[0]))
        q1a8O_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8O_3_1_argbuf_r) && (! q1a8O_3_destruct_bufchan_buf[0])))
        q1a8O_3_destruct_bufchan_buf <= q1a8O_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1a8j_3_destruct,Pointer_QTree_Int) > (q1a8j_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1a8j_3_destruct_bufchan_d;
  logic q1a8j_3_destruct_bufchan_r;
  assign q1a8j_3_destruct_r = ((! q1a8j_3_destruct_bufchan_d[0]) || q1a8j_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8j_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8j_3_destruct_r)
        q1a8j_3_destruct_bufchan_d <= q1a8j_3_destruct_d;
  Pointer_QTree_Int_t q1a8j_3_destruct_bufchan_buf;
  assign q1a8j_3_destruct_bufchan_r = (! q1a8j_3_destruct_bufchan_buf[0]);
  assign q1a8j_3_1_argbuf_d = (q1a8j_3_destruct_bufchan_buf[0] ? q1a8j_3_destruct_bufchan_buf :
                               q1a8j_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8j_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8j_3_1_argbuf_r && q1a8j_3_destruct_bufchan_buf[0]))
        q1a8j_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8j_3_1_argbuf_r) && (! q1a8j_3_destruct_bufchan_buf[0])))
        q1a8j_3_destruct_bufchan_buf <= q1a8j_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a92_destruct,Pointer_QTree_Bool) > (q1a92_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a92_destruct_bufchan_d;
  logic q1a92_destruct_bufchan_r;
  assign q1a92_destruct_r = ((! q1a92_destruct_bufchan_d[0]) || q1a92_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a92_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a92_destruct_r) q1a92_destruct_bufchan_d <= q1a92_destruct_d;
  Pointer_QTree_Bool_t q1a92_destruct_bufchan_buf;
  assign q1a92_destruct_bufchan_r = (! q1a92_destruct_bufchan_buf[0]);
  assign q1a92_1_argbuf_d = (q1a92_destruct_bufchan_buf[0] ? q1a92_destruct_bufchan_buf :
                             q1a92_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a92_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a92_1_argbuf_r && q1a92_destruct_bufchan_buf[0]))
        q1a92_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a92_1_argbuf_r) && (! q1a92_destruct_bufchan_buf[0])))
        q1a92_destruct_bufchan_buf <= q1a92_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8P_2_destruct,Pointer_QTree_Int) > (q2a8P_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8P_2_destruct_bufchan_d;
  logic q2a8P_2_destruct_bufchan_r;
  assign q2a8P_2_destruct_r = ((! q2a8P_2_destruct_bufchan_d[0]) || q2a8P_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8P_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8P_2_destruct_r)
        q2a8P_2_destruct_bufchan_d <= q2a8P_2_destruct_d;
  Pointer_QTree_Int_t q2a8P_2_destruct_bufchan_buf;
  assign q2a8P_2_destruct_bufchan_r = (! q2a8P_2_destruct_bufchan_buf[0]);
  assign q2a8P_2_1_argbuf_d = (q2a8P_2_destruct_bufchan_buf[0] ? q2a8P_2_destruct_bufchan_buf :
                               q2a8P_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8P_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8P_2_1_argbuf_r && q2a8P_2_destruct_bufchan_buf[0]))
        q2a8P_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8P_2_1_argbuf_r) && (! q2a8P_2_destruct_bufchan_buf[0])))
        q2a8P_2_destruct_bufchan_buf <= q2a8P_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2a8k_2_destruct,Pointer_QTree_Int) > (q2a8k_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2a8k_2_destruct_bufchan_d;
  logic q2a8k_2_destruct_bufchan_r;
  assign q2a8k_2_destruct_r = ((! q2a8k_2_destruct_bufchan_d[0]) || q2a8k_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8k_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8k_2_destruct_r)
        q2a8k_2_destruct_bufchan_d <= q2a8k_2_destruct_d;
  Pointer_QTree_Int_t q2a8k_2_destruct_bufchan_buf;
  assign q2a8k_2_destruct_bufchan_r = (! q2a8k_2_destruct_bufchan_buf[0]);
  assign q2a8k_2_1_argbuf_d = (q2a8k_2_destruct_bufchan_buf[0] ? q2a8k_2_destruct_bufchan_buf :
                               q2a8k_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8k_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8k_2_1_argbuf_r && q2a8k_2_destruct_bufchan_buf[0]))
        q2a8k_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8k_2_1_argbuf_r) && (! q2a8k_2_destruct_bufchan_buf[0])))
        q2a8k_2_destruct_bufchan_buf <= q2a8k_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a93_1_destruct,Pointer_QTree_Bool) > (q2a93_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a93_1_destruct_bufchan_d;
  logic q2a93_1_destruct_bufchan_r;
  assign q2a93_1_destruct_r = ((! q2a93_1_destruct_bufchan_d[0]) || q2a93_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a93_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a93_1_destruct_r)
        q2a93_1_destruct_bufchan_d <= q2a93_1_destruct_d;
  Pointer_QTree_Bool_t q2a93_1_destruct_bufchan_buf;
  assign q2a93_1_destruct_bufchan_r = (! q2a93_1_destruct_bufchan_buf[0]);
  assign q2a93_1_1_argbuf_d = (q2a93_1_destruct_bufchan_buf[0] ? q2a93_1_destruct_bufchan_buf :
                               q2a93_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a93_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a93_1_1_argbuf_r && q2a93_1_destruct_bufchan_buf[0]))
        q2a93_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a93_1_1_argbuf_r) && (! q2a93_1_destruct_bufchan_buf[0])))
        q2a93_1_destruct_bufchan_buf <= q2a93_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8Q_1_destruct,Pointer_QTree_Int) > (q3a8Q_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8Q_1_destruct_bufchan_d;
  logic q3a8Q_1_destruct_bufchan_r;
  assign q3a8Q_1_destruct_r = ((! q3a8Q_1_destruct_bufchan_d[0]) || q3a8Q_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8Q_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8Q_1_destruct_r)
        q3a8Q_1_destruct_bufchan_d <= q3a8Q_1_destruct_d;
  Pointer_QTree_Int_t q3a8Q_1_destruct_bufchan_buf;
  assign q3a8Q_1_destruct_bufchan_r = (! q3a8Q_1_destruct_bufchan_buf[0]);
  assign q3a8Q_1_1_argbuf_d = (q3a8Q_1_destruct_bufchan_buf[0] ? q3a8Q_1_destruct_bufchan_buf :
                               q3a8Q_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8Q_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8Q_1_1_argbuf_r && q3a8Q_1_destruct_bufchan_buf[0]))
        q3a8Q_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8Q_1_1_argbuf_r) && (! q3a8Q_1_destruct_bufchan_buf[0])))
        q3a8Q_1_destruct_bufchan_buf <= q3a8Q_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3a8l_1_destruct,Pointer_QTree_Int) > (q3a8l_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3a8l_1_destruct_bufchan_d;
  logic q3a8l_1_destruct_bufchan_r;
  assign q3a8l_1_destruct_r = ((! q3a8l_1_destruct_bufchan_d[0]) || q3a8l_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8l_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8l_1_destruct_r)
        q3a8l_1_destruct_bufchan_d <= q3a8l_1_destruct_d;
  Pointer_QTree_Int_t q3a8l_1_destruct_bufchan_buf;
  assign q3a8l_1_destruct_bufchan_r = (! q3a8l_1_destruct_bufchan_buf[0]);
  assign q3a8l_1_1_argbuf_d = (q3a8l_1_destruct_bufchan_buf[0] ? q3a8l_1_destruct_bufchan_buf :
                               q3a8l_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8l_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8l_1_1_argbuf_r && q3a8l_1_destruct_bufchan_buf[0]))
        q3a8l_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8l_1_1_argbuf_r) && (! q3a8l_1_destruct_bufchan_buf[0])))
        q3a8l_1_destruct_bufchan_buf <= q3a8l_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a94_2_destruct,Pointer_QTree_Bool) > (q3a94_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a94_2_destruct_bufchan_d;
  logic q3a94_2_destruct_bufchan_r;
  assign q3a94_2_destruct_r = ((! q3a94_2_destruct_bufchan_d[0]) || q3a94_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a94_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a94_2_destruct_r)
        q3a94_2_destruct_bufchan_d <= q3a94_2_destruct_d;
  Pointer_QTree_Bool_t q3a94_2_destruct_bufchan_buf;
  assign q3a94_2_destruct_bufchan_r = (! q3a94_2_destruct_bufchan_buf[0]);
  assign q3a94_2_1_argbuf_d = (q3a94_2_destruct_bufchan_buf[0] ? q3a94_2_destruct_bufchan_buf :
                               q3a94_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a94_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a94_2_1_argbuf_r && q3a94_2_destruct_bufchan_buf[0]))
        q3a94_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a94_2_1_argbuf_r) && (! q3a94_2_destruct_bufchan_buf[0])))
        q3a94_2_destruct_bufchan_buf <= q3a94_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4a8R_destruct,Pointer_QTree_Int) > (q4a8R_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4a8R_destruct_bufchan_d;
  logic q4a8R_destruct_bufchan_r;
  assign q4a8R_destruct_r = ((! q4a8R_destruct_bufchan_d[0]) || q4a8R_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8R_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a8R_destruct_r) q4a8R_destruct_bufchan_d <= q4a8R_destruct_d;
  Pointer_QTree_Int_t q4a8R_destruct_bufchan_buf;
  assign q4a8R_destruct_bufchan_r = (! q4a8R_destruct_bufchan_buf[0]);
  assign q4a8R_1_argbuf_d = (q4a8R_destruct_bufchan_buf[0] ? q4a8R_destruct_bufchan_buf :
                             q4a8R_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a8R_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a8R_1_argbuf_r && q4a8R_destruct_bufchan_buf[0]))
        q4a8R_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a8R_1_argbuf_r) && (! q4a8R_destruct_bufchan_buf[0])))
        q4a8R_destruct_bufchan_buf <= q4a8R_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4a95_3_destruct,Pointer_QTree_Bool) > (q4a95_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4a95_3_destruct_bufchan_d;
  logic q4a95_3_destruct_bufchan_r;
  assign q4a95_3_destruct_r = ((! q4a95_3_destruct_bufchan_d[0]) || q4a95_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a95_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4a95_3_destruct_r)
        q4a95_3_destruct_bufchan_d <= q4a95_3_destruct_d;
  Pointer_QTree_Bool_t q4a95_3_destruct_bufchan_buf;
  assign q4a95_3_destruct_bufchan_r = (! q4a95_3_destruct_bufchan_buf[0]);
  assign q4a95_3_1_argbuf_d = (q4a95_3_destruct_bufchan_buf[0] ? q4a95_3_destruct_bufchan_buf :
                               q4a95_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4a95_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4a95_3_1_argbuf_r && q4a95_3_destruct_bufchan_buf[0]))
        q4a95_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4a95_3_1_argbuf_r) && (! q4a95_3_destruct_bufchan_buf[0])))
        q4a95_3_destruct_bufchan_buf <= q4a95_3_destruct_bufchan_d;
  
  /* buf (Ty CT$wmAdd_Int) : (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf,CT$wmAdd_Int) > (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb,CT$wmAdd_Int) */
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                              1'd0};
    else
      if (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_d;
  CT$wmAdd_Int_t readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf :
                                                            readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                1'd0};
    else
      if ((readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                  1'd0};
      else if (((! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wmAdd_Int) : (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb,CT$wmAdd_Int) > [(lizzieLet24_1,CT$wmAdd_Int),
                                                                                         (lizzieLet24_2,CT$wmAdd_Int),
                                                                                         (lizzieLet24_3,CT$wmAdd_Int),
                                                                                         (lizzieLet24_4,CT$wmAdd_Int)] */
  logic [3:0] readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet24_1_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet24_2_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet24_3_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet24_4_d = {readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet24_4_d[0],
                                                                                                                         lizzieLet24_3_d[0],
                                                                                                                         lizzieLet24_2_d[0],
                                                                                                                         lizzieLet24_1_d[0]} & {lizzieLet24_4_r,
                                                                                                                                                lizzieLet24_3_r,
                                                                                                                                                lizzieLet24_2_r,
                                                                                                                                                lizzieLet24_1_r}));
  assign readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                                readPointer_CT$wmAdd_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_1_argbuf,CT$wnnz) > (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb,CT$wnnz) */
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_r = ((! readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d <= {115'd0, 1'd0};
    else
      if (readPointer_CT$wnnzscfarg_0_1_1_argbuf_r)
        readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CT$wnnzscfarg_0_1_1_argbuf_d;
  CT$wnnz_t readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d = (readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf :
                                                         readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                             1'd0};
    else
      if ((readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_r && readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                               1'd0};
      else if (((! readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CT$wnnzscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz) : (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb,CT$wnnz) > [(lizzieLet29_1,CT$wnnz),
                                                                            (lizzieLet29_2,CT$wnnz),
                                                                            (lizzieLet29_3,CT$wnnz),
                                                                            (lizzieLet29_4,CT$wnnz)] */
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet29_1_d = {readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet29_2_d = {readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet29_3_d = {readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet29_4_d = {readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_done = (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet29_4_d[0],
                                                                                                                   lizzieLet29_3_d[0],
                                                                                                                   lizzieLet29_2_d[0],
                                                                                                                   lizzieLet29_1_d[0]} & {lizzieLet29_4_r,
                                                                                                                                          lizzieLet29_3_r,
                                                                                                                                          lizzieLet29_2_r,
                                                                                                                                          lizzieLet29_1_r}));
  assign readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                             readPointer_CT$wnnzscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_map'_Int_Bool) : (readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf,CTmain_map'_Int_Bool) > (readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb,CTmain_map'_Int_Bool) */
  \CTmain_map'_Int_Bool_t  \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d  <= {67'd0,
                                                                          1'd0};
    else
      if (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_r )
        \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_d ;
  \CTmain_map'_Int_Bool_t  \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf  :
                                                                        \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {67'd0,
                                                                            1'd0};
    else
      if ((\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {67'd0,
                                                                              1'd0};
      else if (((! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmain_map'_Int_Bool) : (readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb,CTmain_map'_Int_Bool) > [(lizzieLet33_1,CTmain_map'_Int_Bool),
                                                                                                                   (lizzieLet33_2,CTmain_map'_Int_Bool),
                                                                                                                   (lizzieLet33_3,CTmain_map'_Int_Bool),
                                                                                                                   (lizzieLet33_4,CTmain_map'_Int_Bool)] */
  logic [3:0] \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet33_1_d = {\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet33_2_d = {\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet33_3_d = {\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet33_4_d = {\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet33_4_d[0],
                                                                                                                                                 lizzieLet33_3_d[0],
                                                                                                                                                 lizzieLet33_2_d[0],
                                                                                                                                                 lizzieLet33_1_d[0]} & {lizzieLet33_4_r,
                                                                                                                                                                        lizzieLet33_3_r,
                                                                                                                                                                        lizzieLet33_2_r,
                                                                                                                                                                        lizzieLet33_1_r}));
  assign \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                            \readPointer_CTmain_map'_Int_Boolscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_BoolwslW_1_1_argbuf,QTree_Bool) > (readPointer_QTree_BoolwslW_1_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_BoolwslW_1_1_argbuf_r = ((! readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_BoolwslW_1_1_argbuf_r)
        readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d <= readPointer_QTree_BoolwslW_1_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_r = (! readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d = (readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_BoolwslW_1_1_argbuf_rwb_r && readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_BoolwslW_1_1_argbuf_rwb_r) && (! readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_buf <= readPointer_QTree_BoolwslW_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_BoolwslW_1_1_argbuf_rwb,QTree_Bool) > [(lizzieLet15_1,QTree_Bool),
                                                                                 (lizzieLet15_2,QTree_Bool),
                                                                                 (lizzieLet15_3,QTree_Bool),
                                                                                 (lizzieLet15_4,QTree_Bool)] */
  logic [3:0] readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_BoolwslW_1_1_argbuf_rwb_done;
  assign lizzieLet15_1_d = {readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet15_2_d = {readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet15_3_d = {readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet15_4_d = {readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_BoolwslW_1_1_argbuf_rwb_done = (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted | ({lizzieLet15_4_d[0],
                                                                                                                 lizzieLet15_3_d[0],
                                                                                                                 lizzieLet15_2_d[0],
                                                                                                                 lizzieLet15_1_d[0]} & {lizzieLet15_4_r,
                                                                                                                                        lizzieLet15_3_r,
                                                                                                                                        lizzieLet15_2_r,
                                                                                                                                        lizzieLet15_1_r}));
  assign readPointer_QTree_BoolwslW_1_1_argbuf_rwb_r = (& readPointer_QTree_BoolwslW_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_BoolwslW_1_1_argbuf_rwb_emitted <= (readPointer_QTree_BoolwslW_1_1_argbuf_rwb_r ? 4'd0 :
                                                            readPointer_QTree_BoolwslW_1_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intma8M_1_argbuf,QTree_Int) > (readPointer_QTree_Intma8M_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intma8M_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intma8M_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intma8M_1_argbuf_r = ((! readPointer_QTree_Intma8M_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intma8M_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intma8M_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intma8M_1_argbuf_r)
        readPointer_QTree_Intma8M_1_argbuf_bufchan_d <= readPointer_QTree_Intma8M_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intma8M_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intma8M_1_argbuf_bufchan_r = (! readPointer_QTree_Intma8M_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intma8M_1_argbuf_rwb_d = (readPointer_QTree_Intma8M_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intma8M_1_argbuf_bufchan_buf :
                                                     readPointer_QTree_Intma8M_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intma8M_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intma8M_1_argbuf_rwb_r && readPointer_QTree_Intma8M_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intma8M_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intma8M_1_argbuf_rwb_r) && (! readPointer_QTree_Intma8M_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intma8M_1_argbuf_bufchan_buf <= readPointer_QTree_Intma8M_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intma8M_1_argbuf_rwb,QTree_Int) > [(lizzieLet17_1,QTree_Int),
                                                                            (lizzieLet17_2,QTree_Int),
                                                                            (lizzieLet17_3,QTree_Int),
                                                                            (lizzieLet17_4,QTree_Int),
                                                                            (lizzieLet17_5,QTree_Int),
                                                                            (lizzieLet17_6,QTree_Int)] */
  logic [5:0] readPointer_QTree_Intma8M_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_QTree_Intma8M_1_argbuf_rwb_done;
  assign lizzieLet17_1_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet17_2_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet17_3_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet17_4_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet17_5_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet17_6_d = {readPointer_QTree_Intma8M_1_argbuf_rwb_d[66:1],
                            (readPointer_QTree_Intma8M_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intma8M_1_argbuf_rwb_emitted[5]))};
  assign readPointer_QTree_Intma8M_1_argbuf_rwb_done = (readPointer_QTree_Intma8M_1_argbuf_rwb_emitted | ({lizzieLet17_6_d[0],
                                                                                                           lizzieLet17_5_d[0],
                                                                                                           lizzieLet17_4_d[0],
                                                                                                           lizzieLet17_3_d[0],
                                                                                                           lizzieLet17_2_d[0],
                                                                                                           lizzieLet17_1_d[0]} & {lizzieLet17_6_r,
                                                                                                                                  lizzieLet17_5_r,
                                                                                                                                  lizzieLet17_4_r,
                                                                                                                                  lizzieLet17_3_r,
                                                                                                                                  lizzieLet17_2_r,
                                                                                                                                  lizzieLet17_1_r}));
  assign readPointer_QTree_Intma8M_1_argbuf_rwb_r = (& readPointer_QTree_Intma8M_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intma8M_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_QTree_Intma8M_1_argbuf_rwb_emitted <= (readPointer_QTree_Intma8M_1_argbuf_rwb_r ? 6'd0 :
                                                         readPointer_QTree_Intma8M_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intw1slS_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intw1slS_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intw1slS_1_1_argbuf_r = ((! readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intw1slS_1_1_argbuf_r)
        readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d <= readPointer_QTree_Intw1slS_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d = (readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intw1slS_1_1_argbuf_rwb_r && readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intw1slS_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intw1slS_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet5_1,QTree_Int),
                                                                               (lizzieLet5_2,QTree_Int),
                                                                               (lizzieLet5_3,QTree_Int),
                                                                               (lizzieLet5_4,QTree_Int),
                                                                               (lizzieLet5_5,QTree_Int),
                                                                               (lizzieLet5_6,QTree_Int),
                                                                               (lizzieLet5_7,QTree_Int),
                                                                               (lizzieLet5_8,QTree_Int)] */
  logic [7:0] readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted;
  logic [7:0] readPointer_QTree_Intw1slS_1_1_argbuf_rwb_done;
  assign lizzieLet5_1_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet5_2_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet5_3_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet5_4_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet5_5_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet5_6_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet5_7_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet5_8_d = {readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted[7]))};
  assign readPointer_QTree_Intw1slS_1_1_argbuf_rwb_done = (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted | ({lizzieLet5_8_d[0],
                                                                                                                 lizzieLet5_7_d[0],
                                                                                                                 lizzieLet5_6_d[0],
                                                                                                                 lizzieLet5_5_d[0],
                                                                                                                 lizzieLet5_4_d[0],
                                                                                                                 lizzieLet5_3_d[0],
                                                                                                                 lizzieLet5_2_d[0],
                                                                                                                 lizzieLet5_1_d[0]} & {lizzieLet5_8_r,
                                                                                                                                       lizzieLet5_7_r,
                                                                                                                                       lizzieLet5_6_r,
                                                                                                                                       lizzieLet5_5_r,
                                                                                                                                       lizzieLet5_4_r,
                                                                                                                                       lizzieLet5_3_r,
                                                                                                                                       lizzieLet5_2_r,
                                                                                                                                       lizzieLet5_1_r}));
  assign readPointer_QTree_Intw1slS_1_1_argbuf_rwb_r = (& readPointer_QTree_Intw1slS_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted <= 8'd0;
    else
      readPointer_QTree_Intw1slS_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Intw1slS_1_1_argbuf_rwb_r ? 8'd0 :
                                                            readPointer_QTree_Intw1slS_1_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intw2slT_1_1_argbuf,QTree_Int) > (readPointer_QTree_Intw2slT_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intw2slT_1_1_argbuf_r = ((! readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intw2slT_1_1_argbuf_r)
        readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d <= readPointer_QTree_Intw2slT_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_r = (! readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intw2slT_1_1_argbuf_rwb_d = (readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf :
                                                        readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intw2slT_1_1_argbuf_rwb_r && readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intw2slT_1_1_argbuf_rwb_r) && (! readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_buf <= readPointer_QTree_Intw2slT_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (sc_0_10_destruct,Pointer_CT$wnnz) > (sc_0_10_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  Pointer_CT$wnnz_t sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (sc_0_14_destruct,Pointer_CTmain_map'_Int_Bool) > (sc_0_14_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  \Pointer_CTmain_map'_Int_Bool_t  sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (sc_0_6_destruct,Pointer_CT$wmAdd_Int) > (sc_0_6_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wmAdd_Int_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (scfarg_0_1_goMux_mux,Pointer_CT$wnnz) > (scfarg_0_1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CT$wnnz_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (scfarg_0_2_goMux_mux,Pointer_CTmain_map'_Int_Bool) > (scfarg_0_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTmain_map'_Int_Bool_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Int) > (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wmAdd_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t1a8o_3_destruct,Pointer_QTree_Int) > (t1a8o_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t1a8o_3_destruct_bufchan_d;
  logic t1a8o_3_destruct_bufchan_r;
  assign t1a8o_3_destruct_r = ((! t1a8o_3_destruct_bufchan_d[0]) || t1a8o_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8o_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8o_3_destruct_r)
        t1a8o_3_destruct_bufchan_d <= t1a8o_3_destruct_d;
  Pointer_QTree_Int_t t1a8o_3_destruct_bufchan_buf;
  assign t1a8o_3_destruct_bufchan_r = (! t1a8o_3_destruct_bufchan_buf[0]);
  assign t1a8o_3_1_argbuf_d = (t1a8o_3_destruct_bufchan_buf[0] ? t1a8o_3_destruct_bufchan_buf :
                               t1a8o_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8o_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8o_3_1_argbuf_r && t1a8o_3_destruct_bufchan_buf[0]))
        t1a8o_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8o_3_1_argbuf_r) && (! t1a8o_3_destruct_bufchan_buf[0])))
        t1a8o_3_destruct_bufchan_buf <= t1a8o_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t2a8p_2_destruct,Pointer_QTree_Int) > (t2a8p_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t2a8p_2_destruct_bufchan_d;
  logic t2a8p_2_destruct_bufchan_r;
  assign t2a8p_2_destruct_r = ((! t2a8p_2_destruct_bufchan_d[0]) || t2a8p_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8p_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8p_2_destruct_r)
        t2a8p_2_destruct_bufchan_d <= t2a8p_2_destruct_d;
  Pointer_QTree_Int_t t2a8p_2_destruct_bufchan_buf;
  assign t2a8p_2_destruct_bufchan_r = (! t2a8p_2_destruct_bufchan_buf[0]);
  assign t2a8p_2_1_argbuf_d = (t2a8p_2_destruct_bufchan_buf[0] ? t2a8p_2_destruct_bufchan_buf :
                               t2a8p_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8p_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8p_2_1_argbuf_r && t2a8p_2_destruct_bufchan_buf[0]))
        t2a8p_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8p_2_1_argbuf_r) && (! t2a8p_2_destruct_bufchan_buf[0])))
        t2a8p_2_destruct_bufchan_buf <= t2a8p_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t3a8q_1_destruct,Pointer_QTree_Int) > (t3a8q_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t3a8q_1_destruct_bufchan_d;
  logic t3a8q_1_destruct_bufchan_r;
  assign t3a8q_1_destruct_r = ((! t3a8q_1_destruct_bufchan_d[0]) || t3a8q_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8q_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8q_1_destruct_r)
        t3a8q_1_destruct_bufchan_d <= t3a8q_1_destruct_d;
  Pointer_QTree_Int_t t3a8q_1_destruct_bufchan_buf;
  assign t3a8q_1_destruct_bufchan_r = (! t3a8q_1_destruct_bufchan_buf[0]);
  assign t3a8q_1_1_argbuf_d = (t3a8q_1_destruct_bufchan_buf[0] ? t3a8q_1_destruct_bufchan_buf :
                               t3a8q_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8q_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8q_1_1_argbuf_r && t3a8q_1_destruct_bufchan_buf[0]))
        t3a8q_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8q_1_1_argbuf_r) && (! t3a8q_1_destruct_bufchan_buf[0])))
        t3a8q_1_destruct_bufchan_buf <= t3a8q_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (t4a8r_destruct,Pointer_QTree_Int) > (t4a8r_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t t4a8r_destruct_bufchan_d;
  logic t4a8r_destruct_bufchan_r;
  assign t4a8r_destruct_r = ((! t4a8r_destruct_bufchan_d[0]) || t4a8r_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8r_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8r_destruct_r) t4a8r_destruct_bufchan_d <= t4a8r_destruct_d;
  Pointer_QTree_Int_t t4a8r_destruct_bufchan_buf;
  assign t4a8r_destruct_bufchan_r = (! t4a8r_destruct_bufchan_buf[0]);
  assign t4a8r_1_argbuf_d = (t4a8r_destruct_bufchan_buf[0] ? t4a8r_destruct_bufchan_buf :
                             t4a8r_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8r_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8r_1_argbuf_r && t4a8r_destruct_bufchan_buf[0]))
        t4a8r_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8r_1_argbuf_r) && (! t4a8r_destruct_bufchan_buf[0])))
        t4a8r_destruct_bufchan_buf <= t4a8r_destruct_bufchan_d;
  
  /* buf (Ty Int) : (va8N_destruct,Int) > (va8N_1_argbuf,Int) */
  Int_t va8N_destruct_bufchan_d;
  logic va8N_destruct_bufchan_r;
  assign va8N_destruct_r = ((! va8N_destruct_bufchan_d[0]) || va8N_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8N_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (va8N_destruct_r) va8N_destruct_bufchan_d <= va8N_destruct_d;
  Int_t va8N_destruct_bufchan_buf;
  assign va8N_destruct_bufchan_r = (! va8N_destruct_bufchan_buf[0]);
  assign va8N_1_argbuf_d = (va8N_destruct_bufchan_buf[0] ? va8N_destruct_bufchan_buf :
                            va8N_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8N_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8N_1_argbuf_r && va8N_destruct_bufchan_buf[0]))
        va8N_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8N_1_argbuf_r) && (! va8N_destruct_bufchan_buf[0])))
        va8N_destruct_bufchan_buf <= va8N_destruct_bufchan_d;
  
  /* buf (Ty Int) : (va8e_destruct,Int) > (va8e_1_argbuf,Int) */
  Int_t va8e_destruct_bufchan_d;
  logic va8e_destruct_bufchan_r;
  assign va8e_destruct_r = ((! va8e_destruct_bufchan_d[0]) || va8e_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8e_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (va8e_destruct_r) va8e_destruct_bufchan_d <= va8e_destruct_d;
  Int_t va8e_destruct_bufchan_buf;
  assign va8e_destruct_bufchan_r = (! va8e_destruct_bufchan_buf[0]);
  assign va8e_1_argbuf_d = (va8e_destruct_bufchan_buf[0] ? va8e_destruct_bufchan_buf :
                            va8e_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8e_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((va8e_1_argbuf_r && va8e_destruct_bufchan_buf[0]))
        va8e_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! va8e_1_argbuf_r) && (! va8e_destruct_bufchan_buf[0])))
        va8e_destruct_bufchan_buf <= va8e_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (w1slS_1_1,Pointer_QTree_Int) > (w1slS_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t w1slS_1_1_bufchan_d;
  logic w1slS_1_1_bufchan_r;
  assign w1slS_1_1_r = ((! w1slS_1_1_bufchan_d[0]) || w1slS_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1slS_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w1slS_1_1_r) w1slS_1_1_bufchan_d <= w1slS_1_1_d;
  Pointer_QTree_Int_t w1slS_1_1_bufchan_buf;
  assign w1slS_1_1_bufchan_r = (! w1slS_1_1_bufchan_buf[0]);
  assign w1slS_1_1_argbuf_d = (w1slS_1_1_bufchan_buf[0] ? w1slS_1_1_bufchan_buf :
                               w1slS_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1slS_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w1slS_1_1_argbuf_r && w1slS_1_1_bufchan_buf[0]))
        w1slS_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w1slS_1_1_argbuf_r) && (! w1slS_1_1_bufchan_buf[0])))
        w1slS_1_1_bufchan_buf <= w1slS_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (w1slS_1_goMux_mux,Pointer_QTree_Int) > [(w1slS_1_1,Pointer_QTree_Int),
                                                                       (w1slS_1_2,Pointer_QTree_Int)] */
  logic [1:0] w1slS_1_goMux_mux_emitted;
  logic [1:0] w1slS_1_goMux_mux_done;
  assign w1slS_1_1_d = {w1slS_1_goMux_mux_d[16:1],
                        (w1slS_1_goMux_mux_d[0] && (! w1slS_1_goMux_mux_emitted[0]))};
  assign w1slS_1_2_d = {w1slS_1_goMux_mux_d[16:1],
                        (w1slS_1_goMux_mux_d[0] && (! w1slS_1_goMux_mux_emitted[1]))};
  assign w1slS_1_goMux_mux_done = (w1slS_1_goMux_mux_emitted | ({w1slS_1_2_d[0],
                                                                 w1slS_1_1_d[0]} & {w1slS_1_2_r,
                                                                                    w1slS_1_1_r}));
  assign w1slS_1_goMux_mux_r = (& w1slS_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1slS_1_goMux_mux_emitted <= 2'd0;
    else
      w1slS_1_goMux_mux_emitted <= (w1slS_1_goMux_mux_r ? 2'd0 :
                                    w1slS_1_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Int) : (w2slT_1_1,Pointer_QTree_Int) > (w2slT_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t w2slT_1_1_bufchan_d;
  logic w2slT_1_1_bufchan_r;
  assign w2slT_1_1_r = ((! w2slT_1_1_bufchan_d[0]) || w2slT_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2slT_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w2slT_1_1_r) w2slT_1_1_bufchan_d <= w2slT_1_1_d;
  Pointer_QTree_Int_t w2slT_1_1_bufchan_buf;
  assign w2slT_1_1_bufchan_r = (! w2slT_1_1_bufchan_buf[0]);
  assign w2slT_1_1_argbuf_d = (w2slT_1_1_bufchan_buf[0] ? w2slT_1_1_bufchan_buf :
                               w2slT_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2slT_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w2slT_1_1_argbuf_r && w2slT_1_1_bufchan_buf[0]))
        w2slT_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w2slT_1_1_argbuf_r) && (! w2slT_1_1_bufchan_buf[0])))
        w2slT_1_1_bufchan_buf <= w2slT_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (w2slT_1_goMux_mux,Pointer_QTree_Int) > [(w2slT_1_1,Pointer_QTree_Int),
                                                                       (w2slT_1_2,Pointer_QTree_Int)] */
  logic [1:0] w2slT_1_goMux_mux_emitted;
  logic [1:0] w2slT_1_goMux_mux_done;
  assign w2slT_1_1_d = {w2slT_1_goMux_mux_d[16:1],
                        (w2slT_1_goMux_mux_d[0] && (! w2slT_1_goMux_mux_emitted[0]))};
  assign w2slT_1_2_d = {w2slT_1_goMux_mux_d[16:1],
                        (w2slT_1_goMux_mux_d[0] && (! w2slT_1_goMux_mux_emitted[1]))};
  assign w2slT_1_goMux_mux_done = (w2slT_1_goMux_mux_emitted | ({w2slT_1_2_d[0],
                                                                 w2slT_1_1_d[0]} & {w2slT_1_2_r,
                                                                                    w2slT_1_1_r}));
  assign w2slT_1_goMux_mux_r = (& w2slT_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2slT_1_goMux_mux_emitted <= 2'd0;
    else
      w2slT_1_goMux_mux_emitted <= (w2slT_1_goMux_mux_r ? 2'd0 :
                                    w2slT_1_goMux_mux_done);
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet0_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet0_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                       writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (lizzieLet14_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet12_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet12_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet12_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet12_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca3_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet12_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet25_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet25_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca2_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet26_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet26_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet26_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca1_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet27_1_argbuf,Pointer_CT$wmAdd_Int) > (writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_r = ((! writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet27_1_argbuf_r)
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d <= writeCT$wmAdd_IntlizzieLet27_1_argbuf_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_r = (! writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_d = (writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_r && writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_r) && (! writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_buf <= writeCT$wmAdd_IntlizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Int) : (writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb,Pointer_CT$wmAdd_Int) > (sca0_1_argbuf,Pointer_CT$wmAdd_Int) */
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_r = ((! writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_r)
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Int_t writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet16_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet16_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet16_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet16_1_argbuf_r = ((! writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet16_1_argbuf_r)
        writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet16_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet16_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet16_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet16_1_argbuf_rwb_r && writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet16_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet16_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet16_1_argbuf_rwb,Pointer_CT$wnnz) > (sca3_1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet16_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet16_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet16_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet1_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet1_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet1_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet1_1_argbuf_r = ((! writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet1_1_argbuf_r)
        writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet1_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet1_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet1_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf :
                                                  writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet1_1_argbuf_rwb_r && writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet1_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet1_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet1_1_argbuf_rwb,Pointer_CT$wnnz) > (lizzieLet7_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet1_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet1_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet1_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf :
                                  writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet30_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet30_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet30_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet30_1_argbuf_r = ((! writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet30_1_argbuf_r)
        writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet30_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet30_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet30_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet30_1_argbuf_rwb_r && writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet30_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet30_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet30_1_argbuf_rwb,Pointer_CT$wnnz) > (sca2_1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet30_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet30_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet30_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet31_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet31_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet31_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet31_1_argbuf_r = ((! writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet31_1_argbuf_r)
        writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet31_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet31_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet31_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet31_1_argbuf_rwb_r && writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet31_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet31_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet31_1_argbuf_rwb,Pointer_CT$wnnz) > (sca1_1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet31_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet31_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet31_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet32_1_argbuf,Pointer_CT$wnnz) > (writeCT$wnnzlizzieLet32_1_argbuf_rwb,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d;
  logic writeCT$wnnzlizzieLet32_1_argbuf_bufchan_r;
  assign writeCT$wnnzlizzieLet32_1_argbuf_r = ((! writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d[0]) || writeCT$wnnzlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet32_1_argbuf_r)
        writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d <= writeCT$wnnzlizzieLet32_1_argbuf_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf;
  assign writeCT$wnnzlizzieLet32_1_argbuf_bufchan_r = (! writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnzlizzieLet32_1_argbuf_rwb_d = (writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf[0] ? writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf :
                                                   writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnzlizzieLet32_1_argbuf_rwb_r && writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnzlizzieLet32_1_argbuf_rwb_r) && (! writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeCT$wnnzlizzieLet32_1_argbuf_bufchan_buf <= writeCT$wnnzlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz) : (writeCT$wnnzlizzieLet32_1_argbuf_rwb,Pointer_CT$wnnz) > (sca0_1_1_argbuf,Pointer_CT$wnnz) */
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnzlizzieLet32_1_argbuf_rwb_r = ((! writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnzlizzieLet32_1_argbuf_rwb_r)
        writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d <= writeCT$wnnzlizzieLet32_1_argbuf_rwb_d;
  Pointer_CT$wnnz_t writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf :
                              writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeCT$wnnzlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet21_1_argbuf,Pointer_CTmain_map'_Int_Bool) > (writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_r  = ((! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_r )
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_r  && \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) > (sca3_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet21_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet23_1_argbuf,Pointer_CTmain_map'_Int_Bool) > (writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_r  = ((! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_r )
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_r  && \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) > (lizzieLet4_1_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet4_1_1_argbuf_d = (\writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet23_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet34_1_argbuf,Pointer_CTmain_map'_Int_Bool) > (writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_r  = ((! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_r )
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_r  && \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) > (sca2_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet34_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet35_1_argbuf,Pointer_CTmain_map'_Int_Bool) > (writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_r  = ((! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_r )
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_r  && \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) > (sca1_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet35_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet36_1_argbuf,Pointer_CTmain_map'_Int_Bool) > (writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_r  = ((! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_r )
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_d  = (\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_r  && \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Int_Bool) : (writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb,Pointer_CTmain_map'_Int_Bool) > (sca0_2_1_argbuf,Pointer_CTmain_map'_Int_Bool) */
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_r )
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Int_Bool_t  \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Int_BoollizzieLet36_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet18_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_argbuf_r = ((! writeQTree_BoollizzieLet18_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_argbuf_r)
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet18_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_d = (writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet18_1_argbuf_rwb_r && writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet18_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet18_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet18_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet18_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet19_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_argbuf_r = ((! writeQTree_BoollizzieLet19_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_argbuf_r)
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet19_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_d = (writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet19_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet19_1_argbuf_rwb_r && writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet19_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet19_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet19_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet19_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet19_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet19_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet20_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet20_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet20_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet20_1_argbuf_r = ((! writeQTree_BoollizzieLet20_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet20_1_argbuf_r)
        writeQTree_BoollizzieLet20_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet20_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet20_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet20_1_argbuf_rwb_d = (writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet20_1_argbuf_rwb_r && writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet20_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet20_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet20_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet20_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet20_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet20_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet22_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet22_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet22_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet22_1_argbuf_r = ((! writeQTree_BoollizzieLet22_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet22_1_argbuf_r)
        writeQTree_BoollizzieLet22_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet22_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet22_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet22_1_argbuf_rwb_d = (writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet22_1_argbuf_rwb_r && writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet22_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet22_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet22_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet22_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet22_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet22_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_r = ((! writeQTree_BoollizzieLet37_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_r)
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_d = (writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet37_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet37_1_argbuf_rwb_r && writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet37_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet37_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet37_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet37_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet37_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet11_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_r = ((! writeQTree_IntlizzieLet13_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_r)
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_d = (writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet13_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet13_1_argbuf_rwb_r && writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet13_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet13_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet12_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet13_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet13_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet13_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet14_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_1_argbuf_r = ((! writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_1_argbuf_r)
        writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet14_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet14_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet14_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet14_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet14_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet13_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet14_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf :
                                     writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet14_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_r = ((! writeQTree_IntlizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_r)
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_d = (writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet28_1_argbuf_rwb_r && writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet28_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet28_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet28_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf :
                                                      writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet8_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet8_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_r = ((! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_1_argbuf_r)
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet8_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf :
                                                      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet8_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet8_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet8_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf :
                                                      writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet10_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (wslR_2_2,MyDTInt_Int_Int) > (wslR_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wslR_2_2_bufchan_d;
  logic wslR_2_2_bufchan_r;
  assign wslR_2_2_r = ((! wslR_2_2_bufchan_d[0]) || wslR_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_2_2_bufchan_d <= 1'd0;
    else if (wslR_2_2_r) wslR_2_2_bufchan_d <= wslR_2_2_d;
  MyDTInt_Int_Int_t wslR_2_2_bufchan_buf;
  assign wslR_2_2_bufchan_r = (! wslR_2_2_bufchan_buf[0]);
  assign wslR_2_2_argbuf_d = (wslR_2_2_bufchan_buf[0] ? wslR_2_2_bufchan_buf :
                              wslR_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_2_2_bufchan_buf <= 1'd0;
    else
      if ((wslR_2_2_argbuf_r && wslR_2_2_bufchan_buf[0]))
        wslR_2_2_bufchan_buf <= 1'd0;
      else if (((! wslR_2_2_argbuf_r) && (! wslR_2_2_bufchan_buf[0])))
        wslR_2_2_bufchan_buf <= wslR_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (wslR_2_destruct,MyDTInt_Int_Int) > [(wslR_2_1,MyDTInt_Int_Int),
                                                                 (wslR_2_2,MyDTInt_Int_Int)] */
  logic [1:0] wslR_2_destruct_emitted;
  logic [1:0] wslR_2_destruct_done;
  assign wslR_2_1_d = (wslR_2_destruct_d[0] && (! wslR_2_destruct_emitted[0]));
  assign wslR_2_2_d = (wslR_2_destruct_d[0] && (! wslR_2_destruct_emitted[1]));
  assign wslR_2_destruct_done = (wslR_2_destruct_emitted | ({wslR_2_2_d[0],
                                                             wslR_2_1_d[0]} & {wslR_2_2_r,
                                                                               wslR_2_1_r}));
  assign wslR_2_destruct_r = (& wslR_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_2_destruct_emitted <= 2'd0;
    else
      wslR_2_destruct_emitted <= (wslR_2_destruct_r ? 2'd0 :
                                  wslR_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (wslR_3_2,MyDTInt_Int_Int) > (wslR_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wslR_3_2_bufchan_d;
  logic wslR_3_2_bufchan_r;
  assign wslR_3_2_r = ((! wslR_3_2_bufchan_d[0]) || wslR_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_3_2_bufchan_d <= 1'd0;
    else if (wslR_3_2_r) wslR_3_2_bufchan_d <= wslR_3_2_d;
  MyDTInt_Int_Int_t wslR_3_2_bufchan_buf;
  assign wslR_3_2_bufchan_r = (! wslR_3_2_bufchan_buf[0]);
  assign wslR_3_2_argbuf_d = (wslR_3_2_bufchan_buf[0] ? wslR_3_2_bufchan_buf :
                              wslR_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_3_2_bufchan_buf <= 1'd0;
    else
      if ((wslR_3_2_argbuf_r && wslR_3_2_bufchan_buf[0]))
        wslR_3_2_bufchan_buf <= 1'd0;
      else if (((! wslR_3_2_argbuf_r) && (! wslR_3_2_bufchan_buf[0])))
        wslR_3_2_bufchan_buf <= wslR_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (wslR_3_destruct,MyDTInt_Int_Int) > [(wslR_3_1,MyDTInt_Int_Int),
                                                                 (wslR_3_2,MyDTInt_Int_Int)] */
  logic [1:0] wslR_3_destruct_emitted;
  logic [1:0] wslR_3_destruct_done;
  assign wslR_3_1_d = (wslR_3_destruct_d[0] && (! wslR_3_destruct_emitted[0]));
  assign wslR_3_2_d = (wslR_3_destruct_d[0] && (! wslR_3_destruct_emitted[1]));
  assign wslR_3_destruct_done = (wslR_3_destruct_emitted | ({wslR_3_2_d[0],
                                                             wslR_3_1_d[0]} & {wslR_3_2_r,
                                                                               wslR_3_1_r}));
  assign wslR_3_destruct_r = (& wslR_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_3_destruct_emitted <= 2'd0;
    else
      wslR_3_destruct_emitted <= (wslR_3_destruct_r ? 2'd0 :
                                  wslR_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (wslR_4_destruct,MyDTInt_Int_Int) > (wslR_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t wslR_4_destruct_bufchan_d;
  logic wslR_4_destruct_bufchan_r;
  assign wslR_4_destruct_r = ((! wslR_4_destruct_bufchan_d[0]) || wslR_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_4_destruct_bufchan_d <= 1'd0;
    else
      if (wslR_4_destruct_r)
        wslR_4_destruct_bufchan_d <= wslR_4_destruct_d;
  MyDTInt_Int_Int_t wslR_4_destruct_bufchan_buf;
  assign wslR_4_destruct_bufchan_r = (! wslR_4_destruct_bufchan_buf[0]);
  assign wslR_4_1_argbuf_d = (wslR_4_destruct_bufchan_buf[0] ? wslR_4_destruct_bufchan_buf :
                              wslR_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslR_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((wslR_4_1_argbuf_r && wslR_4_destruct_bufchan_buf[0]))
        wslR_4_destruct_bufchan_buf <= 1'd0;
      else if (((! wslR_4_1_argbuf_r) && (! wslR_4_destruct_bufchan_buf[0])))
        wslR_4_destruct_bufchan_buf <= wslR_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (wslW_1_goMux_mux,Pointer_QTree_Bool) > (wslW_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t wslW_1_goMux_mux_bufchan_d;
  logic wslW_1_goMux_mux_bufchan_r;
  assign wslW_1_goMux_mux_r = ((! wslW_1_goMux_mux_bufchan_d[0]) || wslW_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslW_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wslW_1_goMux_mux_r)
        wslW_1_goMux_mux_bufchan_d <= wslW_1_goMux_mux_d;
  Pointer_QTree_Bool_t wslW_1_goMux_mux_bufchan_buf;
  assign wslW_1_goMux_mux_bufchan_r = (! wslW_1_goMux_mux_bufchan_buf[0]);
  assign wslW_1_1_argbuf_d = (wslW_1_goMux_mux_bufchan_buf[0] ? wslW_1_goMux_mux_bufchan_buf :
                              wslW_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wslW_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wslW_1_1_argbuf_r && wslW_1_goMux_mux_bufchan_buf[0]))
        wslW_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wslW_1_1_argbuf_r) && (! wslW_1_goMux_mux_bufchan_buf[0])))
        wslW_1_goMux_mux_bufchan_buf <= wslW_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz) : (wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1,CT$wnnz) > (lizzieLet31_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d;
  logic wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_r;
  assign wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_r = ((! wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d[0]) || wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d <= {115'd0,
                                                                                      1'd0};
    else
      if (wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_r)
        wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d <= wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_d;
  CT$wnnz_t wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf;
  assign wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_r = (! wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf[0] ? wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf :
                                   wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                        1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf[0]))
        wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf <= {115'd0,
                                                                                          1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf[0])))
        wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_buf <= wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz1) : [(wwslZ_1_destruct,Int#),
                                       (lizzieLet29_4Lcall_$wnnz2,Int#),
                                       (sc_0_8_destruct,Pointer_CT$wnnz),
                                       (q4a95_2_destruct,Pointer_QTree_Bool)] > (wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1,CT$wnnz) */
  assign wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_d = Lcall_$wnnz1_dc((& {wwslZ_1_destruct_d[0],
                                                                                                   lizzieLet29_4Lcall_$wnnz2_d[0],
                                                                                                   sc_0_8_destruct_d[0],
                                                                                                   q4a95_2_destruct_d[0]}), wwslZ_1_destruct_d, lizzieLet29_4Lcall_$wnnz2_d, sc_0_8_destruct_d, q4a95_2_destruct_d);
  assign {wwslZ_1_destruct_r,
          lizzieLet29_4Lcall_$wnnz2_r,
          sc_0_8_destruct_r,
          q4a95_2_destruct_r} = {4 {(wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_r && wwslZ_1_1lizzieLet29_4Lcall_$wnnz2_1sc_0_8_1q4a95_2_1Lcall_$wnnz1_d[0])}};
  
  /* buf (Ty CT$wnnz) : (wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0,CT$wnnz) > (lizzieLet32_1_argbuf,CT$wnnz) */
  CT$wnnz_t wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d;
  logic wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_r;
  assign wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_r = ((! wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d[0]) || wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d <= {115'd0,
                                                                                       1'd0};
    else
      if (wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_r)
        wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d <= wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_d;
  CT$wnnz_t wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf;
  assign wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_r = (! wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf[0] ? wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf :
                                   wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                         1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf[0]))
        wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf <= {115'd0,
                                                                                           1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf[0])))
        wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_buf <= wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_bufchan_d;
  
  /* dcon (Ty CT$wnnz,Dcon Lcall_$wnnz0) : [(wwslZ_2_destruct,Int#),
                                       (ww1XmJ_1_destruct,Int#),
                                       (lizzieLet29_4Lcall_$wnnz1,Int#),
                                       (sc_0_9_destruct,Pointer_CT$wnnz)] > (wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0,CT$wnnz) */
  assign wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_d = Lcall_$wnnz0_dc((& {wwslZ_2_destruct_d[0],
                                                                                                    ww1XmJ_1_destruct_d[0],
                                                                                                    lizzieLet29_4Lcall_$wnnz1_d[0],
                                                                                                    sc_0_9_destruct_d[0]}), wwslZ_2_destruct_d, ww1XmJ_1_destruct_d, lizzieLet29_4Lcall_$wnnz1_d, sc_0_9_destruct_d);
  assign {wwslZ_2_destruct_r,
          ww1XmJ_1_destruct_r,
          lizzieLet29_4Lcall_$wnnz1_r,
          sc_0_9_destruct_r} = {4 {(wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_r && wwslZ_2_1ww1XmJ_1_1lizzieLet29_4Lcall_$wnnz1_1sc_0_9_1Lcall_$wnnz0_d[0])}};
  
  /* op_add (Ty Int#) : (wwslZ_3_1ww1XmJ_2_1_Add32,Int#) (ww2XmM_1_destruct,Int#) > (es_6_1ww2XmM_1_1_Add32,Int#) */
  assign es_6_1ww2XmM_1_1_Add32_d = {(wwslZ_3_1ww1XmJ_2_1_Add32_d[32:1] + ww2XmM_1_destruct_d[32:1]),
                                     (wwslZ_3_1ww1XmJ_2_1_Add32_d[0] && ww2XmM_1_destruct_d[0])};
  assign {wwslZ_3_1ww1XmJ_2_1_Add32_r,
          ww2XmM_1_destruct_r} = {2 {(es_6_1ww2XmM_1_1_Add32_r && es_6_1ww2XmM_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwslZ_3_destruct,Int#) (ww1XmJ_2_destruct,Int#) > (wwslZ_3_1ww1XmJ_2_1_Add32,Int#) */
  assign wwslZ_3_1ww1XmJ_2_1_Add32_d = {(wwslZ_3_destruct_d[32:1] + ww1XmJ_2_destruct_d[32:1]),
                                        (wwslZ_3_destruct_d[0] && ww1XmJ_2_destruct_d[0])};
  assign {wwslZ_3_destruct_r,
          ww1XmJ_2_destruct_r} = {2 {(wwslZ_3_1ww1XmJ_2_1_Add32_r && wwslZ_3_1ww1XmJ_2_1_Add32_d[0])}};
  
  /* buf (Ty MyBool) : (xa88_1,MyBool) > (xa88_1_argbuf,MyBool) */
  MyBool_t xa88_1_bufchan_d;
  logic xa88_1_bufchan_r;
  assign xa88_1_r = ((! xa88_1_bufchan_d[0]) || xa88_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xa88_1_bufchan_d <= {1'd0, 1'd0};
    else if (xa88_1_r) xa88_1_bufchan_d <= xa88_1_d;
  MyBool_t xa88_1_bufchan_buf;
  assign xa88_1_bufchan_r = (! xa88_1_bufchan_buf[0]);
  assign xa88_1_argbuf_d = (xa88_1_bufchan_buf[0] ? xa88_1_bufchan_buf :
                            xa88_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xa88_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((xa88_1_argbuf_r && xa88_1_bufchan_buf[0]))
        xa88_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! xa88_1_argbuf_r) && (! xa88_1_bufchan_buf[0])))
        xa88_1_bufchan_buf <= xa88_1_bufchan_d;
endmodule