`timescale 1ns/1ns
import mMaskAdd_package::*;

module mMaskAdd(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Bool_src_d ,
  output logic \\QTree_Bool_src_r ,
  input QTree_Bool_t dummy_write_QTree_Bool_d,
  output logic dummy_write_QTree_Bool_r,
  input Go_t \\MaskQTree_src_d ,
  output logic \\MaskQTree_src_r ,
  input MaskQTree_t dummy_write_MaskQTree_d,
  output logic dummy_write_MaskQTree_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_MaskQTree_t m1a92_0_d,
  output logic m1a92_0_r,
  input Pointer_QTree_Bool_t m2a93_1_d,
  output logic m2a93_1_r,
  input Pointer_QTree_Bool_t m3a94_2_d,
  output logic m3a94_2_r,
  output \Word16#_t  forkHP1_QTree_Bool_snk_dout,
  input logic forkHP1_QTree_Bool_snk_rout,
  output Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_dout,
  input logic dummy_write_QTree_Bool_sink_rout,
  output \Word16#_t  forkHP1_MaskQTree_snk_dout,
  input logic forkHP1_MaskQTree_snk_rout,
  output Pointer_MaskQTree_t dummy_write_MaskQTree_sink_dout,
  input logic dummy_write_MaskQTree_sink_rout,
  output Pointer_QTree_Bool_t main_mask_Bool_resbuf_dout,
  input logic main_mask_Bool_resbuf_rout
  );
  /* --define=INPUTS=((__05CQTree_Bool_src, 0, 1, Go), (dummy_write_QTree_Bool, 66, 73786976294838206464, QTree_Bool), (__05CMaskQTree_src, 0, 1, Go), (dummy_write_MaskQTree, 66, 73786976294838206464, MaskQTree), (sourceGo, 0, 1, Go), (m1a92_0, 16, 65536, Pointer_MaskQTree), (m2a93_1, 16, 65536, Pointer_QTree_Bool), (m3a94_2, 16, 65536, Pointer_QTree_Bool)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Bool_snk, 16, 65536, Word16__023), (dummy_write_QTree_Bool_sink, 16, 65536, Pointer_QTree_Bool), (forkHP1_MaskQTree_snk, 16, 65536, Word16__023), (dummy_write_MaskQTree_sink, 16, 65536, Pointer_MaskQTree), (main_mask_Bool_resbuf, 16, 65536, Pointer_QTree_Bool)) */
  /* TYPE_START
CT__024wmAdd_Bool 16 3 (0,[0]) (1,[16p,0,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,0,16p,16p,16p,16p]) (3,[16p,16p,16p,0,16p,16p]) (4,[16p,16p,16p,16p])
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTmain_mask_Bool 16 3 (0,[0]) (1,[16p,16p,16p,16p,16p,16p,16p]) (2,[16p,16p,16p,16p,16p,16p]) (3,[16p,16p,16p,16p,16p]) (4,[16p,16p,16p,16p])
MaskQTree 16 2 (0,[0]) (1,[0]) (2,[16p,16p,16p,16p])
TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,0,16p,16p])
TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT__024wmAdd_Bool 16 0 (0,[0,0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool 16 0 (0,[0,16p,16p,16p])
TupGo___Pointer_QTree_Bool___Pointer_MaskQTree 16 0 (0,[0,16p,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go__4_d;
  logic go__4_r;
  Go_t go__5_d;
  logic go__5_r;
  Go_t go__6_d;
  logic go__6_r;
  Go_t go__7_d;
  logic go__7_r;
  \Word16#_t  initHP_CT$wmAdd_Bool_d;
  logic initHP_CT$wmAdd_Bool_r;
  \Word16#_t  incrHP_CT$wmAdd_Bool_d;
  logic incrHP_CT$wmAdd_Bool_r;
  Go_t incrHP_mergeCT$wmAdd_Bool_d;
  logic incrHP_mergeCT$wmAdd_Bool_r;
  Go_t incrHP_CT$wmAdd_Bool1_d;
  logic incrHP_CT$wmAdd_Bool1_r;
  Go_t incrHP_CT$wmAdd_Bool2_d;
  logic incrHP_CT$wmAdd_Bool2_r;
  \Word16#_t  addHP_CT$wmAdd_Bool_d;
  logic addHP_CT$wmAdd_Bool_r;
  \Word16#_t  mergeHP_CT$wmAdd_Bool_d;
  logic mergeHP_CT$wmAdd_Bool_r;
  Go_t incrHP_mergeCT$wmAdd_Bool_buf_d;
  logic incrHP_mergeCT$wmAdd_Bool_buf_r;
  \Word16#_t  mergeHP_CT$wmAdd_Bool_buf_d;
  logic mergeHP_CT$wmAdd_Bool_buf_r;
  \Word16#_t  forkHP1_CT$wmAdd_Bool_d;
  logic forkHP1_CT$wmAdd_Bool_r;
  \Word16#_t  forkHP1_CT$wmAdd_Boo2_d;
  logic forkHP1_CT$wmAdd_Boo2_r;
  \Word16#_t  forkHP1_CT$wmAdd_Boo3_d;
  logic forkHP1_CT$wmAdd_Boo3_r;
  C2_t memMergeChoice_CT$wmAdd_Bool_d;
  logic memMergeChoice_CT$wmAdd_Bool_r;
  MemIn_CT$wmAdd_Bool_t memMergeIn_CT$wmAdd_Bool_d;
  logic memMergeIn_CT$wmAdd_Bool_r;
  MemOut_CT$wmAdd_Bool_t memOut_CT$wmAdd_Bool_d;
  logic memOut_CT$wmAdd_Bool_r;
  MemOut_CT$wmAdd_Bool_t memReadOut_CT$wmAdd_Bool_d;
  logic memReadOut_CT$wmAdd_Bool_r;
  MemOut_CT$wmAdd_Bool_t memWriteOut_CT$wmAdd_Bool_d;
  logic memWriteOut_CT$wmAdd_Bool_r;
  MemIn_CT$wmAdd_Bool_t memMergeIn_CT$wmAdd_Bool_dbuf_d;
  logic memMergeIn_CT$wmAdd_Bool_dbuf_r;
  MemIn_CT$wmAdd_Bool_t memMergeIn_CT$wmAdd_Bool_rbuf_d;
  logic memMergeIn_CT$wmAdd_Bool_rbuf_r;
  MemOut_CT$wmAdd_Bool_t memOut_CT$wmAdd_Bool_dbuf_d;
  logic memOut_CT$wmAdd_Bool_dbuf_r;
  MemOut_CT$wmAdd_Bool_t memOut_CT$wmAdd_Bool_rbuf_d;
  logic memOut_CT$wmAdd_Bool_rbuf_r;
  \Word16#_t  destructReadIn_CT$wmAdd_Bool_d;
  logic destructReadIn_CT$wmAdd_Bool_r;
  MemIn_CT$wmAdd_Bool_t dconReadIn_CT$wmAdd_Bool_d;
  logic dconReadIn_CT$wmAdd_Bool_r;
  CT$wmAdd_Bool_t readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_d;
  logic readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wmAdd_Bool_d;
  logic writeMerge_choice_CT$wmAdd_Bool_r;
  CT$wmAdd_Bool_t writeMerge_data_CT$wmAdd_Bool_d;
  logic writeMerge_data_CT$wmAdd_Bool_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_d;
  logic writeCT$wmAdd_BoollizzieLet0_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_d;
  logic writeCT$wmAdd_BoollizzieLet20_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_d;
  logic writeCT$wmAdd_BoollizzieLet21_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_d;
  logic writeCT$wmAdd_BoollizzieLet22_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_d;
  logic writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_r;
  MemIn_CT$wmAdd_Bool_t dconWriteIn_CT$wmAdd_Bool_d;
  logic dconWriteIn_CT$wmAdd_Bool_r;
  Pointer_CT$wmAdd_Bool_t dconPtr_CT$wmAdd_Bool_d;
  logic dconPtr_CT$wmAdd_Bool_r;
  Pointer_CT$wmAdd_Bool_t _74_d;
  logic _74_r;
  assign _74_r = 1'd1;
  Pointer_CT$wmAdd_Bool_t demuxWriteResult_CT$wmAdd_Bool_d;
  logic demuxWriteResult_CT$wmAdd_Bool_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  Go_t go_1_dummy_write_QTree_Bool_d;
  logic go_1_dummy_write_QTree_Bool_r;
  Go_t go_2_dummy_write_QTree_Bool_d;
  logic go_2_dummy_write_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_snk_d;
  logic forkHP1_QTree_Bool_snk_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  \Word16#_t  forkHP1_QTree_Boo4_d;
  logic forkHP1_QTree_Boo4_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  C3_t readMerge_choice_QTree_Bool_d;
  logic readMerge_choice_QTree_Bool_r;
  Pointer_QTree_Bool_t readMerge_data_QTree_Bool_d;
  logic readMerge_data_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_Boolma8q_1_argbuf_d;
  logic readPointer_QTree_Boolma8q_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolw1sic_1_1_argbuf_d;
  logic readPointer_QTree_Boolw1sic_1_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolw2sid_1_1_argbuf_d;
  logic readPointer_QTree_Boolw2sid_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t destructReadOut_QTree_Bool_d;
  logic destructReadOut_QTree_Bool_r;
  C13_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_d;
  logic dummy_write_QTree_Bool_sink_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _73_d;
  logic _73_r;
  assign _73_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  initHP_CTmain_mask_Bool_d;
  logic initHP_CTmain_mask_Bool_r;
  \Word16#_t  incrHP_CTmain_mask_Bool_d;
  logic incrHP_CTmain_mask_Bool_r;
  Go_t incrHP_mergeCTmain_mask_Bool_d;
  logic incrHP_mergeCTmain_mask_Bool_r;
  Go_t incrHP_CTmain_mask_Bool1_d;
  logic incrHP_CTmain_mask_Bool1_r;
  Go_t incrHP_CTmain_mask_Bool2_d;
  logic incrHP_CTmain_mask_Bool2_r;
  \Word16#_t  addHP_CTmain_mask_Bool_d;
  logic addHP_CTmain_mask_Bool_r;
  \Word16#_t  mergeHP_CTmain_mask_Bool_d;
  logic mergeHP_CTmain_mask_Bool_r;
  Go_t incrHP_mergeCTmain_mask_Bool_buf_d;
  logic incrHP_mergeCTmain_mask_Bool_buf_r;
  \Word16#_t  mergeHP_CTmain_mask_Bool_buf_d;
  logic mergeHP_CTmain_mask_Bool_buf_r;
  \Word16#_t  forkHP1_CTmain_mask_Bool_d;
  logic forkHP1_CTmain_mask_Bool_r;
  \Word16#_t  forkHP1_CTmain_mask_Boo2_d;
  logic forkHP1_CTmain_mask_Boo2_r;
  \Word16#_t  forkHP1_CTmain_mask_Boo3_d;
  logic forkHP1_CTmain_mask_Boo3_r;
  C2_t memMergeChoice_CTmain_mask_Bool_d;
  logic memMergeChoice_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_d;
  logic memMergeIn_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_d;
  logic memOut_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memReadOut_CTmain_mask_Bool_d;
  logic memReadOut_CTmain_mask_Bool_r;
  MemOut_CTmain_mask_Bool_t memWriteOut_CTmain_mask_Bool_d;
  logic memWriteOut_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_dbuf_d;
  logic memMergeIn_CTmain_mask_Bool_dbuf_r;
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_rbuf_d;
  logic memMergeIn_CTmain_mask_Bool_rbuf_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_dbuf_d;
  logic memOut_CTmain_mask_Bool_dbuf_r;
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_rbuf_d;
  logic memOut_CTmain_mask_Bool_rbuf_r;
  \Word16#_t  destructReadIn_CTmain_mask_Bool_d;
  logic destructReadIn_CTmain_mask_Bool_r;
  MemIn_CTmain_mask_Bool_t dconReadIn_CTmain_mask_Bool_d;
  logic dconReadIn_CTmain_mask_Bool_r;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r;
  C5_t writeMerge_choice_CTmain_mask_Bool_d;
  logic writeMerge_choice_CTmain_mask_Bool_r;
  CTmain_mask_Bool_t writeMerge_data_CTmain_mask_Bool_d;
  logic writeMerge_data_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet16_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet25_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_r;
  MemIn_CTmain_mask_Bool_t dconWriteIn_CTmain_mask_Bool_d;
  logic dconWriteIn_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t dconPtr_CTmain_mask_Bool_d;
  logic dconPtr_CTmain_mask_Bool_r;
  Pointer_CTmain_mask_Bool_t _72_d;
  logic _72_r;
  assign _72_r = 1'd1;
  Pointer_CTmain_mask_Bool_t demuxWriteResult_CTmain_mask_Bool_d;
  logic demuxWriteResult_CTmain_mask_Bool_r;
  \Word16#_t  initHP_MaskQTree_d;
  logic initHP_MaskQTree_r;
  \Word16#_t  incrHP_MaskQTree_d;
  logic incrHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_d;
  logic incrHP_mergeMaskQTree_r;
  Go_t incrHP_MaskQTree1_d;
  logic incrHP_MaskQTree1_r;
  Go_t incrHP_MaskQTree2_d;
  logic incrHP_MaskQTree2_r;
  \Word16#_t  addHP_MaskQTree_d;
  logic addHP_MaskQTree_r;
  \Word16#_t  mergeHP_MaskQTree_d;
  logic mergeHP_MaskQTree_r;
  Go_t incrHP_mergeMaskQTree_buf_d;
  logic incrHP_mergeMaskQTree_buf_r;
  \Word16#_t  mergeHP_MaskQTree_buf_d;
  logic mergeHP_MaskQTree_buf_r;
  Go_t go_1_dummy_write_MaskQTree_d;
  logic go_1_dummy_write_MaskQTree_r;
  Go_t go_2_dummy_write_MaskQTree_d;
  logic go_2_dummy_write_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_d;
  logic forkHP1_MaskQTree_r;
  \Word16#_t  forkHP1_MaskQTree_snk_d;
  logic forkHP1_MaskQTree_snk_r;
  \Word16#_t  forkHP1_MaskQTre3_d;
  logic forkHP1_MaskQTre3_r;
  \Word16#_t  forkHP1_MaskQTre4_d;
  logic forkHP1_MaskQTre4_r;
  C2_t memMergeChoice_MaskQTree_d;
  logic memMergeChoice_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_d;
  logic memMergeIn_MaskQTree_r;
  MemOut_MaskQTree_t memOut_MaskQTree_d;
  logic memOut_MaskQTree_r;
  MemOut_MaskQTree_t memReadOut_MaskQTree_d;
  logic memReadOut_MaskQTree_r;
  MemOut_MaskQTree_t memWriteOut_MaskQTree_d;
  logic memWriteOut_MaskQTree_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_dbuf_d;
  logic memMergeIn_MaskQTree_dbuf_r;
  MemIn_MaskQTree_t memMergeIn_MaskQTree_rbuf_d;
  logic memMergeIn_MaskQTree_rbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_dbuf_d;
  logic memOut_MaskQTree_dbuf_r;
  MemOut_MaskQTree_t memOut_MaskQTree_rbuf_d;
  logic memOut_MaskQTree_rbuf_r;
  \Word16#_t  destructReadIn_MaskQTree_d;
  logic destructReadIn_MaskQTree_r;
  MemIn_MaskQTree_t dconReadIn_MaskQTree_d;
  logic dconReadIn_MaskQTree_r;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_r;
  MemIn_MaskQTree_t dconWriteIn_MaskQTree_d;
  logic dconWriteIn_MaskQTree_r;
  Pointer_MaskQTree_t dconPtr_MaskQTree_d;
  logic dconPtr_MaskQTree_r;
  Pointer_MaskQTree_t _71_d;
  logic _71_r;
  assign _71_r = 1'd1;
  Pointer_MaskQTree_t dummy_write_MaskQTree_sink_d;
  logic dummy_write_MaskQTree_sink_r;
  Go_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_r ;
  MyDTBool_Bool_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_r ;
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_r ;
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_r ;
  Go_t go_2_1_d;
  logic go_2_1_r;
  Go_t go_2_2_d;
  logic go_2_2_r;
  Pointer_QTree_Bool_t w1sic_1_argbuf_d;
  logic w1sic_1_argbuf_r;
  Pointer_QTree_Bool_t w2sid_1_argbuf_d;
  logic w2sid_1_argbuf_r;
  MyDTBool_Bool_Bool_t wsib_1_argbuf_d;
  logic wsib_1_argbuf_r;
  Pointer_QTree_Bool_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  Go_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r;
  MyDTBool_Bool_Bool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_r;
  MyDTBool_Bool_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTBool_Bool_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTBool_Bool_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyDTBool_Bool_Bool_t arg0_4_d;
  logic arg0_4_r;
  QTree_Bool_t es_0_1_1QVal_Bool_d;
  logic es_0_1_1QVal_Bool_r;
  MyBool_t \arg0_1Dcon_||_d ;
  logic \arg0_1Dcon_||_r ;
  MyBool_t \arg0_2Dcon_||_d ;
  logic \arg0_2Dcon_||_r ;
  MyBool_t \arg0_2Dcon_||_1_d ;
  logic \arg0_2Dcon_||_1_r ;
  MyBool_t \arg0_2Dcon_||_2_d ;
  logic \arg0_2Dcon_||_2_r ;
  MyBool_t \arg0_2Dcon_||_3_d ;
  logic \arg0_2Dcon_||_3_r ;
  MyBool_t \arg0_2Dcon_||_1MyFalse_d ;
  logic \arg0_2Dcon_||_1MyFalse_r ;
  MyBool_t _70_d;
  logic _70_r;
  assign _70_r = 1'd1;
  MyBool_t applyfnBool_Bool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_Bool_5_resbuf_r;
  Go_t _69_d;
  logic _69_r;
  assign _69_r = 1'd1;
  Go_t \arg0_2Dcon_||_2MyTrue_d ;
  logic \arg0_2Dcon_||_2MyTrue_r ;
  MyBool_t \arg0_2Dcon_||_2MyTrue_1MyTrue_d ;
  logic \arg0_2Dcon_||_2MyTrue_1MyTrue_r ;
  MyBool_t \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d ;
  logic \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_r ;
  Go_t \arg0_3Dcon_||_d ;
  logic \arg0_3Dcon_||_r ;
  MyBool_t \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_d ;
  logic \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_r ;
  Go_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_r;
  MyDTBool_Bool_Bool_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_r;
  Pointer_QTree_Bool_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_r;
  Pointer_QTree_Bool_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_r;
  Pointer_CT$wmAdd_Bool_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_r;
  Go_t call_$wmAdd_Bool_initBufi_d;
  logic call_$wmAdd_Bool_initBufi_r;
  C5_t go_4_goMux_choice_d;
  logic go_4_goMux_choice_r;
  Go_t go_4_goMux_data_d;
  logic go_4_goMux_data_r;
  Go_t call_$wmAdd_Bool_unlockFork1_d;
  logic call_$wmAdd_Bool_unlockFork1_r;
  Go_t call_$wmAdd_Bool_unlockFork2_d;
  logic call_$wmAdd_Bool_unlockFork2_r;
  Go_t call_$wmAdd_Bool_unlockFork3_d;
  logic call_$wmAdd_Bool_unlockFork3_r;
  Go_t call_$wmAdd_Bool_unlockFork4_d;
  logic call_$wmAdd_Bool_unlockFork4_r;
  Go_t call_$wmAdd_Bool_unlockFork5_d;
  logic call_$wmAdd_Bool_unlockFork5_r;
  Go_t call_$wmAdd_Bool_initBuf_d;
  logic call_$wmAdd_Bool_initBuf_r;
  Go_t call_$wmAdd_Bool_goMux1_d;
  logic call_$wmAdd_Bool_goMux1_r;
  MyDTBool_Bool_Bool_t call_$wmAdd_Bool_goMux2_d;
  logic call_$wmAdd_Bool_goMux2_r;
  Pointer_QTree_Bool_t call_$wmAdd_Bool_goMux3_d;
  logic call_$wmAdd_Bool_goMux3_r;
  Pointer_QTree_Bool_t call_$wmAdd_Bool_goMux4_d;
  logic call_$wmAdd_Bool_goMux4_r;
  Pointer_CT$wmAdd_Bool_t call_$wmAdd_Bool_goMux5_d;
  logic call_$wmAdd_Bool_goMux5_r;
  Go_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r;
  Pointer_QTree_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_r;
  Pointer_MaskQTree_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_r;
  Pointer_CTmain_mask_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r;
  Go_t call_main_mask_Bool_initBufi_d;
  logic call_main_mask_Bool_initBufi_r;
  C5_t go_5_goMux_choice_d;
  logic go_5_goMux_choice_r;
  Go_t go_5_goMux_data_d;
  logic go_5_goMux_data_r;
  Go_t call_main_mask_Bool_unlockFork1_d;
  logic call_main_mask_Bool_unlockFork1_r;
  Go_t call_main_mask_Bool_unlockFork2_d;
  logic call_main_mask_Bool_unlockFork2_r;
  Go_t call_main_mask_Bool_unlockFork3_d;
  logic call_main_mask_Bool_unlockFork3_r;
  Go_t call_main_mask_Bool_unlockFork4_d;
  logic call_main_mask_Bool_unlockFork4_r;
  Go_t call_main_mask_Bool_initBuf_d;
  logic call_main_mask_Bool_initBuf_r;
  Go_t call_main_mask_Bool_goMux1_d;
  logic call_main_mask_Bool_goMux1_r;
  Pointer_QTree_Bool_t call_main_mask_Bool_goMux2_d;
  logic call_main_mask_Bool_goMux2_r;
  Pointer_MaskQTree_t call_main_mask_Bool_goMux3_d;
  logic call_main_mask_Bool_goMux3_r;
  Pointer_CTmain_mask_Bool_t call_main_mask_Bool_goMux4_d;
  logic call_main_mask_Bool_goMux4_r;
  QTree_Bool_t lizzieLet3_1_argbuf_d;
  logic lizzieLet3_1_argbuf_r;
  MyDTBool_Bool_Bool_t \go_1Dcon_||_d ;
  logic \go_1Dcon_||_r ;
  MyDTBool_Bool_Bool_t es_2_1_argbuf_d;
  logic es_2_1_argbuf_r;
  Go_t go_2_argbuf_d;
  logic go_2_argbuf_r;
  CT$wmAdd_Bool_t go_2_1L$wmAdd_Boolsbos_d;
  logic go_2_1L$wmAdd_Boolsbos_r;
  CT$wmAdd_Bool_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_2_2_argbuf_d;
  logic go_2_2_argbuf_r;
  TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_t call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d;
  logic call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_r;
  TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ;
  Go_t go_3_argbuf_d;
  logic go_3_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r;
  C5_t go_4_goMux_choice_1_d;
  logic go_4_goMux_choice_1_r;
  C5_t go_4_goMux_choice_2_d;
  logic go_4_goMux_choice_2_r;
  C5_t go_4_goMux_choice_3_d;
  logic go_4_goMux_choice_3_r;
  C5_t go_4_goMux_choice_4_d;
  logic go_4_goMux_choice_4_r;
  MyDTBool_Bool_Bool_t wsib_1_goMux_mux_d;
  logic wsib_1_goMux_mux_r;
  Pointer_QTree_Bool_t w1sic_1_goMux_mux_d;
  logic w1sic_1_goMux_mux_r;
  Pointer_QTree_Bool_t w2sid_1_goMux_mux_d;
  logic w2sid_1_goMux_mux_r;
  Pointer_CT$wmAdd_Bool_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_5_goMux_choice_1_d;
  logic go_5_goMux_choice_1_r;
  C5_t go_5_goMux_choice_2_d;
  logic go_5_goMux_choice_2_r;
  C5_t go_5_goMux_choice_3_d;
  logic go_5_goMux_choice_3_r;
  Pointer_QTree_Bool_t ma8q_goMux_mux_d;
  logic ma8q_goMux_mux_r;
  Pointer_MaskQTree_t mska8r_goMux_mux_d;
  logic mska8r_goMux_mux_r;
  Pointer_CTmain_mask_Bool_t sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  CTmain_mask_Bool_t go_6_1Lmain_mask_Boolsbos_d;
  logic go_6_1Lmain_mask_Boolsbos_r;
  CTmain_mask_Bool_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t go_6_2_argbuf_d;
  logic go_6_2_argbuf_r;
  TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_t call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d;
  logic call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r;
  C10_t go_7_goMux_choice_1_d;
  logic go_7_goMux_choice_1_r;
  C10_t go_7_goMux_choice_2_d;
  logic go_7_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wmAdd_Bool_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C6_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C6_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  Pointer_MaskQTree_t q1a8s_destruct_d;
  logic q1a8s_destruct_r;
  Pointer_MaskQTree_t q2a8t_destruct_d;
  logic q2a8t_destruct_r;
  Pointer_MaskQTree_t q3a8u_destruct_d;
  logic q3a8u_destruct_r;
  Pointer_MaskQTree_t q4a8v_destruct_d;
  logic q4a8v_destruct_r;
  MaskQTree_t _68_d;
  logic _68_r;
  assign _68_r = 1'd1;
  MaskQTree_t _67_d;
  logic _67_r;
  assign _67_r = 1'd1;
  MaskQTree_t lizzieLet11_1_1MQNode_d;
  logic lizzieLet11_1_1MQNode_r;
  Go_t lizzieLet11_1_3MQNone_d;
  logic lizzieLet11_1_3MQNone_r;
  Go_t lizzieLet11_1_3MQVal_d;
  logic lizzieLet11_1_3MQVal_r;
  Go_t lizzieLet11_1_3MQNode_d;
  logic lizzieLet11_1_3MQNode_r;
  Go_t lizzieLet11_1_3MQNone_1_d;
  logic lizzieLet11_1_3MQNone_1_r;
  Go_t lizzieLet11_1_3MQNone_2_d;
  logic lizzieLet11_1_3MQNone_2_r;
  QTree_Bool_t lizzieLet11_1_3MQNone_1QNone_Bool_d;
  logic lizzieLet11_1_3MQNone_1QNone_Bool_r;
  QTree_Bool_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Go_t lizzieLet11_1_3MQNone_2_argbuf_d;
  logic lizzieLet11_1_3MQNone_2_argbuf_r;
  C6_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t lizzieLet11_1_3MQVal_1_argbuf_d;
  logic lizzieLet11_1_3MQVal_1_argbuf_r;
  QTree_Bool_t _66_d;
  logic _66_r;
  assign _66_r = 1'd1;
  QTree_Bool_t _65_d;
  logic _65_r;
  assign _65_r = 1'd1;
  QTree_Bool_t lizzieLet11_1_4MQNode_d;
  logic lizzieLet11_1_4MQNode_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_1_d;
  logic lizzieLet11_1_4MQNode_1_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_2_d;
  logic lizzieLet11_1_4MQNode_2_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_3_d;
  logic lizzieLet11_1_4MQNode_3_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_4_d;
  logic lizzieLet11_1_4MQNode_4_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_5_d;
  logic lizzieLet11_1_4MQNode_5_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_6_d;
  logic lizzieLet11_1_4MQNode_6_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_7_d;
  logic lizzieLet11_1_4MQNode_7_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_8_d;
  logic lizzieLet11_1_4MQNode_8_r;
  Pointer_QTree_Bool_t t1a8x_destruct_d;
  logic t1a8x_destruct_r;
  Pointer_QTree_Bool_t t2a8y_destruct_d;
  logic t2a8y_destruct_r;
  Pointer_QTree_Bool_t t3a8z_destruct_d;
  logic t3a8z_destruct_r;
  Pointer_QTree_Bool_t t4a8A_destruct_d;
  logic t4a8A_destruct_r;
  QTree_Bool_t _64_d;
  logic _64_r;
  assign _64_r = 1'd1;
  QTree_Bool_t _63_d;
  logic _63_r;
  assign _63_r = 1'd1;
  QTree_Bool_t lizzieLet11_1_4MQNode_1QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_1QNode_Bool_r;
  QTree_Bool_t _62_d;
  logic _62_r;
  assign _62_r = 1'd1;
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_r;
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_r;
  Go_t lizzieLet11_1_4MQNode_3QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_3QNode_Bool_r;
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_r;
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_1_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_1_r;
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_2_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_d;
  logic lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_1_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_1_r;
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_2_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_2_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_1_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_1_r;
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_2_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNone_Bool_d;
  logic lizzieLet11_1_4MQNode_4QNone_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QVal_Bool_d;
  logic lizzieLet11_1_4MQNode_4QVal_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_4QNode_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QError_Bool_d;
  logic lizzieLet11_1_4MQNode_4QError_Bool_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_d;
  logic lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d;
  logic lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r;
  CTmain_mask_Bool_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_d;
  logic lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_d;
  logic lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_r;
  Pointer_MaskQTree_t _61_d;
  logic _61_r;
  assign _61_r = 1'd1;
  Pointer_MaskQTree_t _60_d;
  logic _60_r;
  assign _60_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_5QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_5QNode_Bool_r;
  Pointer_MaskQTree_t _59_d;
  logic _59_r;
  assign _59_r = 1'd1;
  Pointer_MaskQTree_t _58_d;
  logic _58_r;
  assign _58_r = 1'd1;
  Pointer_MaskQTree_t _57_d;
  logic _57_r;
  assign _57_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_6QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_6QNode_Bool_r;
  Pointer_MaskQTree_t _56_d;
  logic _56_r;
  assign _56_r = 1'd1;
  Pointer_MaskQTree_t _55_d;
  logic _55_r;
  assign _55_r = 1'd1;
  Pointer_MaskQTree_t _54_d;
  logic _54_r;
  assign _54_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_7QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_7QNode_Bool_r;
  Pointer_MaskQTree_t _53_d;
  logic _53_r;
  assign _53_r = 1'd1;
  Pointer_MaskQTree_t _52_d;
  logic _52_r;
  assign _52_r = 1'd1;
  Pointer_MaskQTree_t _51_d;
  logic _51_r;
  assign _51_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_8QNode_Bool_d;
  logic lizzieLet11_1_4MQNode_8QNode_Bool_r;
  Pointer_MaskQTree_t _50_d;
  logic _50_r;
  assign _50_r = 1'd1;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_d;
  logic lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _49_d;
  logic _49_r;
  assign _49_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet11_1_5MQVal_d;
  logic lizzieLet11_1_5MQVal_r;
  Pointer_QTree_Bool_t _48_d;
  logic _48_r;
  assign _48_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet11_1_5MQVal_1_argbuf_d;
  logic lizzieLet11_1_5MQVal_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQNone_d;
  logic lizzieLet11_1_6MQNone_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQVal_d;
  logic lizzieLet11_1_6MQVal_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQNode_d;
  logic lizzieLet11_1_6MQNode_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQNone_1_argbuf_d;
  logic lizzieLet11_1_6MQNone_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQVal_1_argbuf_d;
  logic lizzieLet11_1_6MQVal_1_argbuf_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_QTree_Bool_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  Pointer_CT$wmAdd_Bool_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Bool_t es_3_destruct_d;
  logic es_3_destruct_r;
  Pointer_QTree_Bool_t es_4_1_destruct_d;
  logic es_4_1_destruct_r;
  Pointer_CT$wmAdd_Bool_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  MyDTBool_Bool_Bool_t wsib_4_destruct_d;
  logic wsib_4_destruct_r;
  Pointer_QTree_Bool_t q1a8h_3_destruct_d;
  logic q1a8h_3_destruct_r;
  Pointer_QTree_Bool_t t1a8m_3_destruct_d;
  logic t1a8m_3_destruct_r;
  Pointer_QTree_Bool_t es_4_destruct_d;
  logic es_4_destruct_r;
  Pointer_CT$wmAdd_Bool_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  MyDTBool_Bool_Bool_t wsib_3_destruct_d;
  logic wsib_3_destruct_r;
  Pointer_QTree_Bool_t q1a8h_2_destruct_d;
  logic q1a8h_2_destruct_r;
  Pointer_QTree_Bool_t t1a8m_2_destruct_d;
  logic t1a8m_2_destruct_r;
  Pointer_QTree_Bool_t q2a8i_2_destruct_d;
  logic q2a8i_2_destruct_r;
  Pointer_QTree_Bool_t t2a8n_2_destruct_d;
  logic t2a8n_2_destruct_r;
  Pointer_CT$wmAdd_Bool_t sc_0_2_destruct_d;
  logic sc_0_2_destruct_r;
  MyDTBool_Bool_Bool_t wsib_2_destruct_d;
  logic wsib_2_destruct_r;
  Pointer_QTree_Bool_t q1a8h_1_destruct_d;
  logic q1a8h_1_destruct_r;
  Pointer_QTree_Bool_t t1a8m_1_destruct_d;
  logic t1a8m_1_destruct_r;
  Pointer_QTree_Bool_t q2a8i_1_destruct_d;
  logic q2a8i_1_destruct_r;
  Pointer_QTree_Bool_t t2a8n_1_destruct_d;
  logic t2a8n_1_destruct_r;
  Pointer_QTree_Bool_t q3a8j_1_destruct_d;
  logic q3a8j_1_destruct_r;
  Pointer_QTree_Bool_t t3a8o_1_destruct_d;
  logic t3a8o_1_destruct_r;
  CT$wmAdd_Bool_t _47_d;
  logic _47_r;
  assign _47_r = 1'd1;
  CT$wmAdd_Bool_t lizzieLet19_1Lcall_$wmAdd_Bool3_d;
  logic lizzieLet19_1Lcall_$wmAdd_Bool3_r;
  CT$wmAdd_Bool_t lizzieLet19_1Lcall_$wmAdd_Bool2_d;
  logic lizzieLet19_1Lcall_$wmAdd_Bool2_r;
  CT$wmAdd_Bool_t lizzieLet19_1Lcall_$wmAdd_Bool1_d;
  logic lizzieLet19_1Lcall_$wmAdd_Bool1_r;
  CT$wmAdd_Bool_t lizzieLet19_1Lcall_$wmAdd_Bool0_d;
  logic lizzieLet19_1Lcall_$wmAdd_Bool0_r;
  Go_t _46_d;
  logic _46_r;
  assign _46_r = 1'd1;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool3_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool3_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool2_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool2_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool1_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool1_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool0_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool0_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet19_4L$wmAdd_Boolsbos_d;
  logic lizzieLet19_4L$wmAdd_Boolsbos_r;
  Pointer_QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool3_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool3_r;
  Pointer_QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool2_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool2_r;
  Pointer_QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool1_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool1_r;
  Pointer_QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool0_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool0_r;
  Pointer_QTree_Bool_t lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_d;
  logic lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_d;
  logic lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_r;
  Go_t call_$wmAdd_Bool_goConst_d;
  logic call_$wmAdd_Bool_goConst_r;
  Pointer_QTree_Bool_t \$wmAdd_Bool_resbuf_d ;
  logic \$wmAdd_Bool_resbuf_r ;
  QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_r;
  QTree_Bool_t lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_r;
  CT$wmAdd_Bool_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_r;
  CT$wmAdd_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_r;
  CT$wmAdd_Bool_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Pointer_QTree_Bool_t q1a8h_destruct_d;
  logic q1a8h_destruct_r;
  Pointer_QTree_Bool_t q2a8i_destruct_d;
  logic q2a8i_destruct_r;
  Pointer_QTree_Bool_t q3a8j_destruct_d;
  logic q3a8j_destruct_r;
  Pointer_QTree_Bool_t q4a8k_destruct_d;
  logic q4a8k_destruct_r;
  MyBool_t v1a8b_destruct_d;
  logic v1a8b_destruct_r;
  QTree_Bool_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  QTree_Bool_t lizzieLet1_1QVal_Bool_d;
  logic lizzieLet1_1QVal_Bool_r;
  QTree_Bool_t lizzieLet1_1QNode_Bool_d;
  logic lizzieLet1_1QNode_Bool_r;
  QTree_Bool_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Go_t lizzieLet1_3QNone_Bool_d;
  logic lizzieLet1_3QNone_Bool_r;
  Go_t lizzieLet1_3QVal_Bool_d;
  logic lizzieLet1_3QVal_Bool_r;
  Go_t lizzieLet1_3QNode_Bool_d;
  logic lizzieLet1_3QNode_Bool_r;
  Go_t lizzieLet1_3QError_Bool_d;
  logic lizzieLet1_3QError_Bool_r;
  Go_t lizzieLet1_3QError_Bool_1_d;
  logic lizzieLet1_3QError_Bool_1_r;
  Go_t lizzieLet1_3QError_Bool_2_d;
  logic lizzieLet1_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet1_3QError_Bool_1QError_Bool_d;
  logic lizzieLet1_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Go_t lizzieLet1_3QError_Bool_2_argbuf_d;
  logic lizzieLet1_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet1_3QNone_Bool_1_argbuf_d;
  logic lizzieLet1_3QNone_Bool_1_argbuf_r;
  C10_t go_7_goMux_choice_d;
  logic go_7_goMux_choice_r;
  Go_t go_7_goMux_data_d;
  logic go_7_goMux_data_r;
  QTree_Bool_t _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  QTree_Bool_t lizzieLet1_4QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_r;
  QTree_Bool_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  QTree_Bool_t lizzieLet1_4QNode_Bool_1_d;
  logic lizzieLet1_4QNode_Bool_1_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_2_d;
  logic lizzieLet1_4QNode_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_3_d;
  logic lizzieLet1_4QNode_Bool_3_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_4_d;
  logic lizzieLet1_4QNode_Bool_4_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_5_d;
  logic lizzieLet1_4QNode_Bool_5_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_6_d;
  logic lizzieLet1_4QNode_Bool_6_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_7_d;
  logic lizzieLet1_4QNode_Bool_7_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_8_d;
  logic lizzieLet1_4QNode_Bool_8_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_9_d;
  logic lizzieLet1_4QNode_Bool_9_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_10_d;
  logic lizzieLet1_4QNode_Bool_10_r;
  Pointer_QTree_Bool_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  Pointer_QTree_Bool_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_10QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_10QNode_Bool_r;
  Pointer_QTree_Bool_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8m_destruct_d;
  logic t1a8m_destruct_r;
  Pointer_QTree_Bool_t t2a8n_destruct_d;
  logic t2a8n_destruct_r;
  Pointer_QTree_Bool_t t3a8o_destruct_d;
  logic t3a8o_destruct_r;
  Pointer_QTree_Bool_t t4a8p_destruct_d;
  logic t4a8p_destruct_r;
  QTree_Bool_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  QTree_Bool_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  QTree_Bool_t lizzieLet1_4QNode_Bool_1QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_1QNode_Bool_r;
  QTree_Bool_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  Go_t lizzieLet1_4QNode_Bool_3QNone_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QNone_Bool_r;
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_r;
  Go_t lizzieLet1_4QNode_Bool_3QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QNode_Bool_r;
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_r;
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_1_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_1_r;
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_2_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_r;
  Go_t lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_1_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_2_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNone_Bool_d;
  logic lizzieLet1_4QNode_Bool_4QNone_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QVal_Bool_d;
  logic lizzieLet1_4QNode_Bool_4QVal_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_4QNode_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QError_Bool_d;
  logic lizzieLet1_4QNode_Bool_4QError_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_r;
  CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_d;
  logic lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_r;
  CT$wmAdd_Bool_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_5QNone_Bool_d;
  logic lizzieLet1_4QNode_Bool_5QNone_Bool_r;
  Pointer_QTree_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_QTree_Bool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Pointer_QTree_Bool_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_r;
  MyDTBool_Bool_Bool_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  MyDTBool_Bool_Bool_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_6QNode_Bool_r;
  MyDTBool_Bool_Bool_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_1_d;
  logic lizzieLet1_4QNode_Bool_6QNode_Bool_1_r;
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_2_d;
  logic lizzieLet1_4QNode_Bool_6QNode_Bool_2_r;
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_d;
  logic lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  Pointer_QTree_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_7QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_7QNode_Bool_r;
  Pointer_QTree_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  Pointer_QTree_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  Pointer_QTree_Bool_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_8QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_8QNode_Bool_r;
  Pointer_QTree_Bool_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Bool_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Bool_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_9QNode_Bool_d;
  logic lizzieLet1_4QNode_Bool_9QNode_Bool_r;
  Pointer_QTree_Bool_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  QTree_Bool_t lizzieLet1_4QVal_Bool_1_d;
  logic lizzieLet1_4QVal_Bool_1_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_2_d;
  logic lizzieLet1_4QVal_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_3_d;
  logic lizzieLet1_4QVal_Bool_3_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_4_d;
  logic lizzieLet1_4QVal_Bool_4_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_5_d;
  logic lizzieLet1_4QVal_Bool_5_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_6_d;
  logic lizzieLet1_4QVal_Bool_6_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_7_d;
  logic lizzieLet1_4QVal_Bool_7_r;
  MyBool_t va8c_destruct_d;
  logic va8c_destruct_r;
  QTree_Bool_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  QTree_Bool_t lizzieLet1_4QVal_Bool_1QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_1QVal_Bool_r;
  QTree_Bool_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  QTree_Bool_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Go_t lizzieLet1_4QVal_Bool_3QNone_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QNone_Bool_r;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_r;
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_r;
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_r;
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_1_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_1_r;
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_2_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_r;
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_1_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_1_r;
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_2_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_2_r;
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_r;
  Go_t lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_r;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_1_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_1_r;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_2_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_2_r;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNone_Bool_d;
  logic lizzieLet1_4QVal_Bool_4QNone_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_4QVal_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNode_Bool_d;
  logic lizzieLet1_4QVal_Bool_4QNode_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QError_Bool_d;
  logic lizzieLet1_4QVal_Bool_4QError_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet1_4QVal_Bool_5QNone_Bool_d;
  logic lizzieLet1_4QVal_Bool_5QNone_Bool_r;
  Pointer_QTree_Bool_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Pointer_QTree_Bool_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Pointer_QTree_Bool_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_r;
  MyDTBool_Bool_Bool_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet1_4QVal_Bool_6QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_6QVal_Bool_r;
  MyDTBool_Bool_Bool_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  MyDTBool_Bool_Bool_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_r;
  MyBool_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  MyBool_t lizzieLet1_4QVal_Bool_7QVal_Bool_d;
  logic lizzieLet1_4QVal_Bool_7QVal_Bool_r;
  MyBool_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  MyBool_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  MyBool_t lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_d;
  logic lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QNone_Bool_d;
  logic lizzieLet1_5QNone_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QVal_Bool_d;
  logic lizzieLet1_5QVal_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QNode_Bool_d;
  logic lizzieLet1_5QNode_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QError_Bool_d;
  logic lizzieLet1_5QError_Bool_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QError_Bool_1_argbuf_d;
  logic lizzieLet1_5QError_Bool_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QNone_Bool_1_argbuf_d;
  logic lizzieLet1_5QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_6QVal_Bool_d;
  logic lizzieLet1_6QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet1_6QNode_Bool_d;
  logic lizzieLet1_6QNode_Bool_r;
  Pointer_QTree_Bool_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_7QNone_Bool_d;
  logic lizzieLet1_7QNone_Bool_r;
  Pointer_QTree_Bool_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Pointer_QTree_Bool_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  Pointer_QTree_Bool_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet1_7QNone_Bool_1_argbuf_d;
  logic lizzieLet1_7QNone_Bool_1_argbuf_r;
  MyDTBool_Bool_Bool_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet1_8QVal_Bool_d;
  logic lizzieLet1_8QVal_Bool_r;
  MyDTBool_Bool_Bool_t lizzieLet1_8QNode_Bool_d;
  logic lizzieLet1_8QNode_Bool_r;
  MyDTBool_Bool_Bool_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  Pointer_QTree_Bool_t es_1_destruct_d;
  logic es_1_destruct_r;
  Pointer_QTree_Bool_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Bool_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Bool_t t1a8x_3_destruct_d;
  logic t1a8x_3_destruct_r;
  Pointer_MaskQTree_t q1a8s_3_destruct_d;
  logic q1a8s_3_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Bool_t t1a8x_2_destruct_d;
  logic t1a8x_2_destruct_r;
  Pointer_MaskQTree_t q1a8s_2_destruct_d;
  logic q1a8s_2_destruct_r;
  Pointer_QTree_Bool_t t2a8y_2_destruct_d;
  logic t2a8y_2_destruct_r;
  Pointer_MaskQTree_t q2a8t_2_destruct_d;
  logic q2a8t_2_destruct_r;
  Pointer_CTmain_mask_Bool_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Bool_t t1a8x_1_destruct_d;
  logic t1a8x_1_destruct_r;
  Pointer_MaskQTree_t q1a8s_1_destruct_d;
  logic q1a8s_1_destruct_r;
  Pointer_QTree_Bool_t t2a8y_1_destruct_d;
  logic t2a8y_1_destruct_r;
  Pointer_MaskQTree_t q2a8t_1_destruct_d;
  logic q2a8t_1_destruct_r;
  Pointer_QTree_Bool_t t3a8z_1_destruct_d;
  logic t3a8z_1_destruct_r;
  Pointer_MaskQTree_t q3a8u_1_destruct_d;
  logic q3a8u_1_destruct_r;
  CTmain_mask_Bool_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  CTmain_mask_Bool_t lizzieLet24_1Lcall_main_mask_Bool3_d;
  logic lizzieLet24_1Lcall_main_mask_Bool3_r;
  CTmain_mask_Bool_t lizzieLet24_1Lcall_main_mask_Bool2_d;
  logic lizzieLet24_1Lcall_main_mask_Bool2_r;
  CTmain_mask_Bool_t lizzieLet24_1Lcall_main_mask_Bool1_d;
  logic lizzieLet24_1Lcall_main_mask_Bool1_r;
  CTmain_mask_Bool_t lizzieLet24_1Lcall_main_mask_Bool0_d;
  logic lizzieLet24_1Lcall_main_mask_Bool0_r;
  Go_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Go_t lizzieLet24_3Lcall_main_mask_Bool3_d;
  logic lizzieLet24_3Lcall_main_mask_Bool3_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool2_d;
  logic lizzieLet24_3Lcall_main_mask_Bool2_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool1_d;
  logic lizzieLet24_3Lcall_main_mask_Bool1_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool0_d;
  logic lizzieLet24_3Lcall_main_mask_Bool0_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_d;
  logic lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_d;
  logic lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_d;
  logic lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_d;
  logic lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lmain_mask_Boolsbos_d;
  logic lizzieLet24_4Lmain_mask_Boolsbos_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool3_d;
  logic lizzieLet24_4Lcall_main_mask_Bool3_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool2_d;
  logic lizzieLet24_4Lcall_main_mask_Bool2_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool1_d;
  logic lizzieLet24_4Lcall_main_mask_Bool1_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool0_d;
  logic lizzieLet24_4Lcall_main_mask_Bool0_r;
  QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_d;
  logic lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_r;
  QTree_Bool_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_d;
  logic lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_r;
  CTmain_mask_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_d;
  logic lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_r;
  CTmain_mask_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_d;
  logic lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_r;
  CTmain_mask_Bool_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d;
  logic lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d;
  logic lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r;
  Go_t call_main_mask_Bool_goConst_d;
  logic call_main_mask_Bool_goConst_r;
  Pointer_QTree_Bool_t main_mask_Bool_resbuf_d;
  logic main_mask_Bool_resbuf_r;
  Pointer_QTree_Bool_t ma8q_1_argbuf_d;
  logic ma8q_1_argbuf_r;
  Pointer_QTree_Bool_t ma8q_1_d;
  logic ma8q_1_r;
  Pointer_QTree_Bool_t ma8q_2_d;
  logic ma8q_2_r;
  Go_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_r;
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_r;
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_r;
  Go_t go_6_1_d;
  logic go_6_1_r;
  Go_t go_6_2_d;
  logic go_6_2_r;
  Pointer_QTree_Bool_t ma8q_1_1_argbuf_d;
  logic ma8q_1_1_argbuf_r;
  Pointer_MaskQTree_t mska8r_1_1_argbuf_d;
  logic mska8r_1_1_argbuf_r;
  Pointer_MaskQTree_t mska8r_1_argbuf_d;
  logic mska8r_1_argbuf_r;
  Pointer_QTree_Bool_t q1a8h_3_1_argbuf_d;
  logic q1a8h_3_1_argbuf_r;
  Pointer_MaskQTree_t q1a8s_3_1_argbuf_d;
  logic q1a8s_3_1_argbuf_r;
  Pointer_QTree_Bool_t q2a8i_2_1_argbuf_d;
  logic q2a8i_2_1_argbuf_r;
  Pointer_MaskQTree_t q2a8t_2_1_argbuf_d;
  logic q2a8t_2_1_argbuf_r;
  Pointer_QTree_Bool_t q3a8j_1_1_argbuf_d;
  logic q3a8j_1_1_argbuf_r;
  Pointer_MaskQTree_t q3a8u_1_1_argbuf_d;
  logic q3a8u_1_1_argbuf_r;
  CT$wmAdd_Bool_t readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_r;
  CT$wmAdd_Bool_t lizzieLet19_1_d;
  logic lizzieLet19_1_r;
  CT$wmAdd_Bool_t lizzieLet19_2_d;
  logic lizzieLet19_2_r;
  CT$wmAdd_Bool_t lizzieLet19_3_d;
  logic lizzieLet19_3_r;
  CT$wmAdd_Bool_t lizzieLet19_4_d;
  logic lizzieLet19_4_r;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r;
  CTmain_mask_Bool_t lizzieLet24_1_d;
  logic lizzieLet24_1_r;
  CTmain_mask_Bool_t lizzieLet24_2_d;
  logic lizzieLet24_2_r;
  CTmain_mask_Bool_t lizzieLet24_3_d;
  logic lizzieLet24_3_r;
  CTmain_mask_Bool_t lizzieLet24_4_d;
  logic lizzieLet24_4_r;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_rwb_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_rwb_r;
  MaskQTree_t lizzieLet11_1_1_d;
  logic lizzieLet11_1_1_r;
  MaskQTree_t lizzieLet11_1_2_d;
  logic lizzieLet11_1_2_r;
  MaskQTree_t lizzieLet11_1_3_d;
  logic lizzieLet11_1_3_r;
  MaskQTree_t lizzieLet11_1_4_d;
  logic lizzieLet11_1_4_r;
  MaskQTree_t lizzieLet11_1_5_d;
  logic lizzieLet11_1_5_r;
  MaskQTree_t lizzieLet11_1_6_d;
  logic lizzieLet11_1_6_r;
  QTree_Bool_t readPointer_QTree_Boolma8q_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolma8q_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet1_1_d;
  logic lizzieLet1_1_r;
  QTree_Bool_t lizzieLet1_2_d;
  logic lizzieLet1_2_r;
  QTree_Bool_t lizzieLet1_3_d;
  logic lizzieLet1_3_r;
  QTree_Bool_t lizzieLet1_4_d;
  logic lizzieLet1_4_r;
  QTree_Bool_t lizzieLet1_5_d;
  logic lizzieLet1_5_r;
  QTree_Bool_t lizzieLet1_6_d;
  logic lizzieLet1_6_r;
  QTree_Bool_t lizzieLet1_7_d;
  logic lizzieLet1_7_r;
  QTree_Bool_t lizzieLet1_8_d;
  logic lizzieLet1_8_r;
  QTree_Bool_t readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t sc_0_5_1_argbuf_d;
  logic sc_0_5_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t sc_0_9_1_argbuf_d;
  logic sc_0_9_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8m_3_1_argbuf_d;
  logic t1a8m_3_1_argbuf_r;
  Pointer_QTree_Bool_t t1a8x_3_1_argbuf_d;
  logic t1a8x_3_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8n_2_1_argbuf_d;
  logic t2a8n_2_1_argbuf_r;
  Pointer_QTree_Bool_t t2a8y_2_1_argbuf_d;
  logic t2a8y_2_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8o_1_1_argbuf_d;
  logic t3a8o_1_1_argbuf_r;
  Pointer_QTree_Bool_t t3a8z_1_1_argbuf_d;
  logic t3a8z_1_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8A_1_argbuf_d;
  logic t4a8A_1_argbuf_r;
  Pointer_QTree_Bool_t t4a8p_1_argbuf_d;
  logic t4a8p_1_argbuf_r;
  MyBool_t va8c_1_argbuf_d;
  logic va8c_1_argbuf_r;
  Pointer_QTree_Bool_t w1sic_1_1_argbuf_d;
  logic w1sic_1_1_argbuf_r;
  Pointer_QTree_Bool_t w1sic_1_1_d;
  logic w1sic_1_1_r;
  Pointer_QTree_Bool_t w1sic_1_2_d;
  logic w1sic_1_2_r;
  Pointer_QTree_Bool_t w2sid_1_1_argbuf_d;
  logic w2sid_1_1_argbuf_r;
  Pointer_QTree_Bool_t w2sid_1_1_d;
  logic w2sid_1_1_r;
  Pointer_QTree_Bool_t w2sid_1_2_d;
  logic w2sid_1_2_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_d;
  logic writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_d;
  logic writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_d;
  logic writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_d;
  logic writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_r;
  Pointer_CT$wmAdd_Bool_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r;
  Pointer_CTmain_mask_Bool_t sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet0_1_1_argbuf_d;
  logic lizzieLet0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_argbuf_d;
  logic lizzieLet6_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet5_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet7_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  MyDTBool_Bool_Bool_t wsib_2_2_argbuf_d;
  logic wsib_2_2_argbuf_r;
  MyDTBool_Bool_Bool_t wsib_2_1_d;
  logic wsib_2_1_r;
  MyDTBool_Bool_Bool_t wsib_2_2_d;
  logic wsib_2_2_r;
  MyDTBool_Bool_Bool_t wsib_3_2_argbuf_d;
  logic wsib_3_2_argbuf_r;
  MyDTBool_Bool_Bool_t wsib_3_1_d;
  logic wsib_3_1_r;
  MyDTBool_Bool_Bool_t wsib_3_2_d;
  logic wsib_3_2_r;
  MyDTBool_Bool_Bool_t wsib_4_1_argbuf_d;
  logic wsib_4_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go__4,Go),
                                (go__5,Go),
                                (go__6,Go),
                                (go__7,Go)] */
  logic [6:0] sourceGo_emitted;
  logic [6:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go__4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go__5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go__6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign sourceGo_done = (sourceGo_emitted | ({go__7_d[0],
                                               go__6_d[0],
                                               go__5_d[0],
                                               go__4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__7_r,
                                                             go__6_r,
                                                             go__5_r,
                                                             go__4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 7'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 7'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go__4,Go) > (initHP_CT$wmAdd_Bool,Word16#) */
  assign initHP_CT$wmAdd_Bool_d = {16'd0, go__4_d[0]};
  assign go__4_r = initHP_CT$wmAdd_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wmAdd_Bool1,Go) > (incrHP_CT$wmAdd_Bool,Word16#) */
  assign incrHP_CT$wmAdd_Bool_d = {16'd1,
                                   incrHP_CT$wmAdd_Bool1_d[0]};
  assign incrHP_CT$wmAdd_Bool1_r = incrHP_CT$wmAdd_Bool_r;
  
  /* merge (Ty Go) : [(go__5,Go),
                 (incrHP_CT$wmAdd_Bool2,Go)] > (incrHP_mergeCT$wmAdd_Bool,Go) */
  logic [1:0] incrHP_mergeCT$wmAdd_Bool_selected;
  logic [1:0] incrHP_mergeCT$wmAdd_Bool_select;
  always_comb
    begin
      incrHP_mergeCT$wmAdd_Bool_selected = 2'd0;
      if ((| incrHP_mergeCT$wmAdd_Bool_select))
        incrHP_mergeCT$wmAdd_Bool_selected = incrHP_mergeCT$wmAdd_Bool_select;
      else
        if (go__5_d[0]) incrHP_mergeCT$wmAdd_Bool_selected[0] = 1'd1;
        else if (incrHP_CT$wmAdd_Bool2_d[0])
          incrHP_mergeCT$wmAdd_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Bool_select <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Bool_select <= (incrHP_mergeCT$wmAdd_Bool_r ? 2'd0 :
                                           incrHP_mergeCT$wmAdd_Bool_selected);
  always_comb
    if (incrHP_mergeCT$wmAdd_Bool_selected[0])
      incrHP_mergeCT$wmAdd_Bool_d = go__5_d;
    else if (incrHP_mergeCT$wmAdd_Bool_selected[1])
      incrHP_mergeCT$wmAdd_Bool_d = incrHP_CT$wmAdd_Bool2_d;
    else incrHP_mergeCT$wmAdd_Bool_d = 1'd0;
  assign {incrHP_CT$wmAdd_Bool2_r,
          go__5_r} = (incrHP_mergeCT$wmAdd_Bool_r ? incrHP_mergeCT$wmAdd_Bool_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wmAdd_Bool_buf,Go) > [(incrHP_CT$wmAdd_Bool1,Go),
                                                     (incrHP_CT$wmAdd_Bool2,Go)] */
  logic [1:0] incrHP_mergeCT$wmAdd_Bool_buf_emitted;
  logic [1:0] incrHP_mergeCT$wmAdd_Bool_buf_done;
  assign incrHP_CT$wmAdd_Bool1_d = (incrHP_mergeCT$wmAdd_Bool_buf_d[0] && (! incrHP_mergeCT$wmAdd_Bool_buf_emitted[0]));
  assign incrHP_CT$wmAdd_Bool2_d = (incrHP_mergeCT$wmAdd_Bool_buf_d[0] && (! incrHP_mergeCT$wmAdd_Bool_buf_emitted[1]));
  assign incrHP_mergeCT$wmAdd_Bool_buf_done = (incrHP_mergeCT$wmAdd_Bool_buf_emitted | ({incrHP_CT$wmAdd_Bool2_d[0],
                                                                                         incrHP_CT$wmAdd_Bool1_d[0]} & {incrHP_CT$wmAdd_Bool2_r,
                                                                                                                        incrHP_CT$wmAdd_Bool1_r}));
  assign incrHP_mergeCT$wmAdd_Bool_buf_r = (& incrHP_mergeCT$wmAdd_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wmAdd_Bool_buf_emitted <= (incrHP_mergeCT$wmAdd_Bool_buf_r ? 2'd0 :
                                                incrHP_mergeCT$wmAdd_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wmAdd_Bool,Word16#) (forkHP1_CT$wmAdd_Bool,Word16#) > (addHP_CT$wmAdd_Bool,Word16#) */
  assign addHP_CT$wmAdd_Bool_d = {(incrHP_CT$wmAdd_Bool_d[16:1] + forkHP1_CT$wmAdd_Bool_d[16:1]),
                                  (incrHP_CT$wmAdd_Bool_d[0] && forkHP1_CT$wmAdd_Bool_d[0])};
  assign {incrHP_CT$wmAdd_Bool_r,
          forkHP1_CT$wmAdd_Bool_r} = {2 {(addHP_CT$wmAdd_Bool_r && addHP_CT$wmAdd_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wmAdd_Bool,Word16#),
                      (addHP_CT$wmAdd_Bool,Word16#)] > (mergeHP_CT$wmAdd_Bool,Word16#) */
  logic [1:0] mergeHP_CT$wmAdd_Bool_selected;
  logic [1:0] mergeHP_CT$wmAdd_Bool_select;
  always_comb
    begin
      mergeHP_CT$wmAdd_Bool_selected = 2'd0;
      if ((| mergeHP_CT$wmAdd_Bool_select))
        mergeHP_CT$wmAdd_Bool_selected = mergeHP_CT$wmAdd_Bool_select;
      else
        if (initHP_CT$wmAdd_Bool_d[0])
          mergeHP_CT$wmAdd_Bool_selected[0] = 1'd1;
        else if (addHP_CT$wmAdd_Bool_d[0])
          mergeHP_CT$wmAdd_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Bool_select <= 2'd0;
    else
      mergeHP_CT$wmAdd_Bool_select <= (mergeHP_CT$wmAdd_Bool_r ? 2'd0 :
                                       mergeHP_CT$wmAdd_Bool_selected);
  always_comb
    if (mergeHP_CT$wmAdd_Bool_selected[0])
      mergeHP_CT$wmAdd_Bool_d = initHP_CT$wmAdd_Bool_d;
    else if (mergeHP_CT$wmAdd_Bool_selected[1])
      mergeHP_CT$wmAdd_Bool_d = addHP_CT$wmAdd_Bool_d;
    else mergeHP_CT$wmAdd_Bool_d = {16'd0, 1'd0};
  assign {addHP_CT$wmAdd_Bool_r,
          initHP_CT$wmAdd_Bool_r} = (mergeHP_CT$wmAdd_Bool_r ? mergeHP_CT$wmAdd_Bool_selected :
                                     2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wmAdd_Bool,Go) > (incrHP_mergeCT$wmAdd_Bool_buf,Go) */
  Go_t incrHP_mergeCT$wmAdd_Bool_bufchan_d;
  logic incrHP_mergeCT$wmAdd_Bool_bufchan_r;
  assign incrHP_mergeCT$wmAdd_Bool_r = ((! incrHP_mergeCT$wmAdd_Bool_bufchan_d[0]) || incrHP_mergeCT$wmAdd_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wmAdd_Bool_r)
        incrHP_mergeCT$wmAdd_Bool_bufchan_d <= incrHP_mergeCT$wmAdd_Bool_d;
  Go_t incrHP_mergeCT$wmAdd_Bool_bufchan_buf;
  assign incrHP_mergeCT$wmAdd_Bool_bufchan_r = (! incrHP_mergeCT$wmAdd_Bool_bufchan_buf[0]);
  assign incrHP_mergeCT$wmAdd_Bool_buf_d = (incrHP_mergeCT$wmAdd_Bool_bufchan_buf[0] ? incrHP_mergeCT$wmAdd_Bool_bufchan_buf :
                                            incrHP_mergeCT$wmAdd_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wmAdd_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wmAdd_Bool_buf_r && incrHP_mergeCT$wmAdd_Bool_bufchan_buf[0]))
        incrHP_mergeCT$wmAdd_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wmAdd_Bool_buf_r) && (! incrHP_mergeCT$wmAdd_Bool_bufchan_buf[0])))
        incrHP_mergeCT$wmAdd_Bool_bufchan_buf <= incrHP_mergeCT$wmAdd_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wmAdd_Bool,Word16#) > (mergeHP_CT$wmAdd_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wmAdd_Bool_bufchan_d;
  logic mergeHP_CT$wmAdd_Bool_bufchan_r;
  assign mergeHP_CT$wmAdd_Bool_r = ((! mergeHP_CT$wmAdd_Bool_bufchan_d[0]) || mergeHP_CT$wmAdd_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wmAdd_Bool_r)
        mergeHP_CT$wmAdd_Bool_bufchan_d <= mergeHP_CT$wmAdd_Bool_d;
  \Word16#_t  mergeHP_CT$wmAdd_Bool_bufchan_buf;
  assign mergeHP_CT$wmAdd_Bool_bufchan_r = (! mergeHP_CT$wmAdd_Bool_bufchan_buf[0]);
  assign mergeHP_CT$wmAdd_Bool_buf_d = (mergeHP_CT$wmAdd_Bool_bufchan_buf[0] ? mergeHP_CT$wmAdd_Bool_bufchan_buf :
                                        mergeHP_CT$wmAdd_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wmAdd_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wmAdd_Bool_buf_r && mergeHP_CT$wmAdd_Bool_bufchan_buf[0]))
        mergeHP_CT$wmAdd_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wmAdd_Bool_buf_r) && (! mergeHP_CT$wmAdd_Bool_bufchan_buf[0])))
        mergeHP_CT$wmAdd_Bool_bufchan_buf <= mergeHP_CT$wmAdd_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wmAdd_Bool_buf,Word16#) > [(forkHP1_CT$wmAdd_Bool,Word16#),
                                                           (forkHP1_CT$wmAdd_Boo2,Word16#),
                                                           (forkHP1_CT$wmAdd_Boo3,Word16#)] */
  logic [2:0] mergeHP_CT$wmAdd_Bool_buf_emitted;
  logic [2:0] mergeHP_CT$wmAdd_Bool_buf_done;
  assign forkHP1_CT$wmAdd_Bool_d = {mergeHP_CT$wmAdd_Bool_buf_d[16:1],
                                    (mergeHP_CT$wmAdd_Bool_buf_d[0] && (! mergeHP_CT$wmAdd_Bool_buf_emitted[0]))};
  assign forkHP1_CT$wmAdd_Boo2_d = {mergeHP_CT$wmAdd_Bool_buf_d[16:1],
                                    (mergeHP_CT$wmAdd_Bool_buf_d[0] && (! mergeHP_CT$wmAdd_Bool_buf_emitted[1]))};
  assign forkHP1_CT$wmAdd_Boo3_d = {mergeHP_CT$wmAdd_Bool_buf_d[16:1],
                                    (mergeHP_CT$wmAdd_Bool_buf_d[0] && (! mergeHP_CT$wmAdd_Bool_buf_emitted[2]))};
  assign mergeHP_CT$wmAdd_Bool_buf_done = (mergeHP_CT$wmAdd_Bool_buf_emitted | ({forkHP1_CT$wmAdd_Boo3_d[0],
                                                                                 forkHP1_CT$wmAdd_Boo2_d[0],
                                                                                 forkHP1_CT$wmAdd_Bool_d[0]} & {forkHP1_CT$wmAdd_Boo3_r,
                                                                                                                forkHP1_CT$wmAdd_Boo2_r,
                                                                                                                forkHP1_CT$wmAdd_Bool_r}));
  assign mergeHP_CT$wmAdd_Bool_buf_r = (& mergeHP_CT$wmAdd_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wmAdd_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wmAdd_Bool_buf_emitted <= (mergeHP_CT$wmAdd_Bool_buf_r ? 3'd0 :
                                            mergeHP_CT$wmAdd_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wmAdd_Bool) : [(dconReadIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool),
                                      (dconWriteIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool)] > (memMergeChoice_CT$wmAdd_Bool,C2) (memMergeIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool) */
  logic [1:0] dconReadIn_CT$wmAdd_Bool_select_d;
  assign dconReadIn_CT$wmAdd_Bool_select_d = ((| dconReadIn_CT$wmAdd_Bool_select_q) ? dconReadIn_CT$wmAdd_Bool_select_q :
                                              (dconReadIn_CT$wmAdd_Bool_d[0] ? 2'd1 :
                                               (dconWriteIn_CT$wmAdd_Bool_d[0] ? 2'd2 :
                                                2'd0)));
  logic [1:0] dconReadIn_CT$wmAdd_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Bool_select_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Bool_select_q <= (dconReadIn_CT$wmAdd_Bool_done ? 2'd0 :
                                            dconReadIn_CT$wmAdd_Bool_select_d);
  logic [1:0] dconReadIn_CT$wmAdd_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wmAdd_Bool_emit_q <= 2'd0;
    else
      dconReadIn_CT$wmAdd_Bool_emit_q <= (dconReadIn_CT$wmAdd_Bool_done ? 2'd0 :
                                          dconReadIn_CT$wmAdd_Bool_emit_d);
  logic [1:0] dconReadIn_CT$wmAdd_Bool_emit_d;
  assign dconReadIn_CT$wmAdd_Bool_emit_d = (dconReadIn_CT$wmAdd_Bool_emit_q | ({memMergeChoice_CT$wmAdd_Bool_d[0],
                                                                                memMergeIn_CT$wmAdd_Bool_d[0]} & {memMergeChoice_CT$wmAdd_Bool_r,
                                                                                                                  memMergeIn_CT$wmAdd_Bool_r}));
  logic dconReadIn_CT$wmAdd_Bool_done;
  assign dconReadIn_CT$wmAdd_Bool_done = (& dconReadIn_CT$wmAdd_Bool_emit_d);
  assign {dconWriteIn_CT$wmAdd_Bool_r,
          dconReadIn_CT$wmAdd_Bool_r} = (dconReadIn_CT$wmAdd_Bool_done ? dconReadIn_CT$wmAdd_Bool_select_d :
                                         2'd0);
  assign memMergeIn_CT$wmAdd_Bool_d = ((dconReadIn_CT$wmAdd_Bool_select_d[0] && (! dconReadIn_CT$wmAdd_Bool_emit_q[0])) ? dconReadIn_CT$wmAdd_Bool_d :
                                       ((dconReadIn_CT$wmAdd_Bool_select_d[1] && (! dconReadIn_CT$wmAdd_Bool_emit_q[0])) ? dconWriteIn_CT$wmAdd_Bool_d :
                                        {132'd0, 1'd0}));
  assign memMergeChoice_CT$wmAdd_Bool_d = ((dconReadIn_CT$wmAdd_Bool_select_d[0] && (! dconReadIn_CT$wmAdd_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                           ((dconReadIn_CT$wmAdd_Bool_select_d[1] && (! dconReadIn_CT$wmAdd_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                            {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wmAdd_Bool,
      Ty MemOut_CT$wmAdd_Bool) : (memMergeIn_CT$wmAdd_Bool_dbuf,MemIn_CT$wmAdd_Bool) > (memOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool) */
  logic [114:0] memMergeIn_CT$wmAdd_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wmAdd_Bool_dbuf_address;
  logic [114:0] memMergeIn_CT$wmAdd_Bool_dbuf_din;
  logic [114:0] memOut_CT$wmAdd_Bool_q;
  logic memOut_CT$wmAdd_Bool_valid;
  logic memMergeIn_CT$wmAdd_Bool_dbuf_we;
  logic memOut_CT$wmAdd_Bool_we;
  assign memMergeIn_CT$wmAdd_Bool_dbuf_din = memMergeIn_CT$wmAdd_Bool_dbuf_d[132:18];
  assign memMergeIn_CT$wmAdd_Bool_dbuf_address = memMergeIn_CT$wmAdd_Bool_dbuf_d[17:2];
  assign memMergeIn_CT$wmAdd_Bool_dbuf_we = (memMergeIn_CT$wmAdd_Bool_dbuf_d[1:1] && memMergeIn_CT$wmAdd_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wmAdd_Bool_we <= 1'd0;
        memOut_CT$wmAdd_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wmAdd_Bool_we <= memMergeIn_CT$wmAdd_Bool_dbuf_we;
        memOut_CT$wmAdd_Bool_valid <= memMergeIn_CT$wmAdd_Bool_dbuf_d[0];
        if (memMergeIn_CT$wmAdd_Bool_dbuf_we)
          begin
            memMergeIn_CT$wmAdd_Bool_dbuf_mem[memMergeIn_CT$wmAdd_Bool_dbuf_address] <= memMergeIn_CT$wmAdd_Bool_dbuf_din;
            memOut_CT$wmAdd_Bool_q <= memMergeIn_CT$wmAdd_Bool_dbuf_din;
          end
        else
          memOut_CT$wmAdd_Bool_q <= memMergeIn_CT$wmAdd_Bool_dbuf_mem[memMergeIn_CT$wmAdd_Bool_dbuf_address];
      end
  assign memOut_CT$wmAdd_Bool_d = {memOut_CT$wmAdd_Bool_q,
                                   memOut_CT$wmAdd_Bool_we,
                                   memOut_CT$wmAdd_Bool_valid};
  assign memMergeIn_CT$wmAdd_Bool_dbuf_r = ((! memOut_CT$wmAdd_Bool_valid) || memOut_CT$wmAdd_Bool_r);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wmAdd_Bool) : (memMergeChoice_CT$wmAdd_Bool,C2) (memOut_CT$wmAdd_Bool_dbuf,MemOut_CT$wmAdd_Bool) > [(memReadOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool),
                                                                                                                        (memWriteOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool)] */
  logic [1:0] memOut_CT$wmAdd_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wmAdd_Bool_d[0] && memOut_CT$wmAdd_Bool_dbuf_d[0]))
      unique case (memMergeChoice_CT$wmAdd_Bool_d[1:1])
        1'd0: memOut_CT$wmAdd_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wmAdd_Bool_dbuf_onehotd = 2'd2;
        default: memOut_CT$wmAdd_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wmAdd_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wmAdd_Bool_d = {memOut_CT$wmAdd_Bool_dbuf_d[116:1],
                                       memOut_CT$wmAdd_Bool_dbuf_onehotd[0]};
  assign memWriteOut_CT$wmAdd_Bool_d = {memOut_CT$wmAdd_Bool_dbuf_d[116:1],
                                        memOut_CT$wmAdd_Bool_dbuf_onehotd[1]};
  assign memOut_CT$wmAdd_Bool_dbuf_r = (| (memOut_CT$wmAdd_Bool_dbuf_onehotd & {memWriteOut_CT$wmAdd_Bool_r,
                                                                                memReadOut_CT$wmAdd_Bool_r}));
  assign memMergeChoice_CT$wmAdd_Bool_r = memOut_CT$wmAdd_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wmAdd_Bool) : (memMergeIn_CT$wmAdd_Bool_rbuf,MemIn_CT$wmAdd_Bool) > (memMergeIn_CT$wmAdd_Bool_dbuf,MemIn_CT$wmAdd_Bool) */
  assign memMergeIn_CT$wmAdd_Bool_rbuf_r = ((! memMergeIn_CT$wmAdd_Bool_dbuf_d[0]) || memMergeIn_CT$wmAdd_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wmAdd_Bool_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wmAdd_Bool_rbuf_r)
        memMergeIn_CT$wmAdd_Bool_dbuf_d <= memMergeIn_CT$wmAdd_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wmAdd_Bool) : (memMergeIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool) > (memMergeIn_CT$wmAdd_Bool_rbuf,MemIn_CT$wmAdd_Bool) */
  MemIn_CT$wmAdd_Bool_t memMergeIn_CT$wmAdd_Bool_buf;
  assign memMergeIn_CT$wmAdd_Bool_r = (! memMergeIn_CT$wmAdd_Bool_buf[0]);
  assign memMergeIn_CT$wmAdd_Bool_rbuf_d = (memMergeIn_CT$wmAdd_Bool_buf[0] ? memMergeIn_CT$wmAdd_Bool_buf :
                                            memMergeIn_CT$wmAdd_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wmAdd_Bool_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wmAdd_Bool_rbuf_r && memMergeIn_CT$wmAdd_Bool_buf[0]))
        memMergeIn_CT$wmAdd_Bool_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wmAdd_Bool_rbuf_r) && (! memMergeIn_CT$wmAdd_Bool_buf[0])))
        memMergeIn_CT$wmAdd_Bool_buf <= memMergeIn_CT$wmAdd_Bool_d;
  
  /* dbuf (Ty MemOut_CT$wmAdd_Bool) : (memOut_CT$wmAdd_Bool_rbuf,MemOut_CT$wmAdd_Bool) > (memOut_CT$wmAdd_Bool_dbuf,MemOut_CT$wmAdd_Bool) */
  assign memOut_CT$wmAdd_Bool_rbuf_r = ((! memOut_CT$wmAdd_Bool_dbuf_d[0]) || memOut_CT$wmAdd_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Bool_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wmAdd_Bool_rbuf_r)
        memOut_CT$wmAdd_Bool_dbuf_d <= memOut_CT$wmAdd_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wmAdd_Bool) : (memOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool) > (memOut_CT$wmAdd_Bool_rbuf,MemOut_CT$wmAdd_Bool) */
  MemOut_CT$wmAdd_Bool_t memOut_CT$wmAdd_Bool_buf;
  assign memOut_CT$wmAdd_Bool_r = (! memOut_CT$wmAdd_Bool_buf[0]);
  assign memOut_CT$wmAdd_Bool_rbuf_d = (memOut_CT$wmAdd_Bool_buf[0] ? memOut_CT$wmAdd_Bool_buf :
                                        memOut_CT$wmAdd_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wmAdd_Bool_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wmAdd_Bool_rbuf_r && memOut_CT$wmAdd_Bool_buf[0]))
        memOut_CT$wmAdd_Bool_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wmAdd_Bool_rbuf_r) && (! memOut_CT$wmAdd_Bool_buf[0])))
        memOut_CT$wmAdd_Bool_buf <= memOut_CT$wmAdd_Bool_d;
  
  /* destruct (Ty Pointer_CT$wmAdd_Bool,
          Dcon Pointer_CT$wmAdd_Bool) : (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Bool) > [(destructReadIn_CT$wmAdd_Bool,Word16#)] */
  assign destructReadIn_CT$wmAdd_Bool_d = {scfarg_0_1_argbuf_d[16:1],
                                           scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wmAdd_Bool_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Bool,
      Dcon ReadIn_CT$wmAdd_Bool) : [(destructReadIn_CT$wmAdd_Bool,Word16#)] > (dconReadIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool) */
  assign dconReadIn_CT$wmAdd_Bool_d = ReadIn_CT$wmAdd_Bool_dc((& {destructReadIn_CT$wmAdd_Bool_d[0]}), destructReadIn_CT$wmAdd_Bool_d);
  assign {destructReadIn_CT$wmAdd_Bool_r} = {1 {(dconReadIn_CT$wmAdd_Bool_r && dconReadIn_CT$wmAdd_Bool_d[0])}};
  
  /* destruct (Ty MemOut_CT$wmAdd_Bool,
          Dcon ReadOut_CT$wmAdd_Bool) : (memReadOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool) > [(readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf,CT$wmAdd_Bool)] */
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_d = {memReadOut_CT$wmAdd_Bool_d[116:2],
                                                         memReadOut_CT$wmAdd_Bool_d[0]};
  assign memReadOut_CT$wmAdd_Bool_r = readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wmAdd_Bool) : [(lizzieLet0_1_argbuf,CT$wmAdd_Bool),
                                (lizzieLet20_1_argbuf,CT$wmAdd_Bool),
                                (lizzieLet21_1_argbuf,CT$wmAdd_Bool),
                                (lizzieLet22_1_argbuf,CT$wmAdd_Bool),
                                (lizzieLet8_1_1_argbuf,CT$wmAdd_Bool)] > (writeMerge_choice_CT$wmAdd_Bool,C5) (writeMerge_data_CT$wmAdd_Bool,CT$wmAdd_Bool) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet20_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet21_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet22_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet8_1_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wmAdd_Bool_d[0],
                                                                      writeMerge_data_CT$wmAdd_Bool_d[0]} & {writeMerge_choice_CT$wmAdd_Bool_r,
                                                                                                             writeMerge_data_CT$wmAdd_Bool_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet8_1_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wmAdd_Bool_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                              ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                               ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet8_1_1_argbuf_d :
                                                {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wmAdd_Bool_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                 ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                  {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wmAdd_Bool) : (writeMerge_choice_CT$wmAdd_Bool,C5) (demuxWriteResult_CT$wmAdd_Bool,Pointer_CT$wmAdd_Bool) > [(writeCT$wmAdd_BoollizzieLet0_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                                                                                                  (writeCT$wmAdd_BoollizzieLet20_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                                                                                                  (writeCT$wmAdd_BoollizzieLet21_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                                                                                                  (writeCT$wmAdd_BoollizzieLet22_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                                                                                                  (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf,Pointer_CT$wmAdd_Bool)] */
  logic [4:0] demuxWriteResult_CT$wmAdd_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wmAdd_Bool_d[0] && demuxWriteResult_CT$wmAdd_Bool_d[0]))
      unique case (writeMerge_choice_CT$wmAdd_Bool_d[3:1])
        3'd0: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd16;
        default: demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wmAdd_Bool_onehotd = 5'd0;
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Bool_d[16:1],
                                                    demuxWriteResult_CT$wmAdd_Bool_onehotd[0]};
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Bool_d[16:1],
                                                     demuxWriteResult_CT$wmAdd_Bool_onehotd[1]};
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Bool_d[16:1],
                                                     demuxWriteResult_CT$wmAdd_Bool_onehotd[2]};
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Bool_d[16:1],
                                                     demuxWriteResult_CT$wmAdd_Bool_onehotd[3]};
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_d = {demuxWriteResult_CT$wmAdd_Bool_d[16:1],
                                                      demuxWriteResult_CT$wmAdd_Bool_onehotd[4]};
  assign demuxWriteResult_CT$wmAdd_Bool_r = (| (demuxWriteResult_CT$wmAdd_Bool_onehotd & {writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_r,
                                                                                          writeCT$wmAdd_BoollizzieLet22_1_argbuf_r,
                                                                                          writeCT$wmAdd_BoollizzieLet21_1_argbuf_r,
                                                                                          writeCT$wmAdd_BoollizzieLet20_1_argbuf_r,
                                                                                          writeCT$wmAdd_BoollizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wmAdd_Bool_r = demuxWriteResult_CT$wmAdd_Bool_r;
  
  /* dcon (Ty MemIn_CT$wmAdd_Bool,
      Dcon WriteIn_CT$wmAdd_Bool) : [(forkHP1_CT$wmAdd_Boo2,Word16#),
                                     (writeMerge_data_CT$wmAdd_Bool,CT$wmAdd_Bool)] > (dconWriteIn_CT$wmAdd_Bool,MemIn_CT$wmAdd_Bool) */
  assign dconWriteIn_CT$wmAdd_Bool_d = WriteIn_CT$wmAdd_Bool_dc((& {forkHP1_CT$wmAdd_Boo2_d[0],
                                                                    writeMerge_data_CT$wmAdd_Bool_d[0]}), forkHP1_CT$wmAdd_Boo2_d, writeMerge_data_CT$wmAdd_Bool_d);
  assign {forkHP1_CT$wmAdd_Boo2_r,
          writeMerge_data_CT$wmAdd_Bool_r} = {2 {(dconWriteIn_CT$wmAdd_Bool_r && dconWriteIn_CT$wmAdd_Bool_d[0])}};
  
  /* dcon (Ty Pointer_CT$wmAdd_Bool,
      Dcon Pointer_CT$wmAdd_Bool) : [(forkHP1_CT$wmAdd_Boo3,Word16#)] > (dconPtr_CT$wmAdd_Bool,Pointer_CT$wmAdd_Bool) */
  assign dconPtr_CT$wmAdd_Bool_d = Pointer_CT$wmAdd_Bool_dc((& {forkHP1_CT$wmAdd_Boo3_d[0]}), forkHP1_CT$wmAdd_Boo3_d);
  assign {forkHP1_CT$wmAdd_Boo3_r} = {1 {(dconPtr_CT$wmAdd_Bool_r && dconPtr_CT$wmAdd_Bool_d[0])}};
  
  /* demux (Ty MemOut_CT$wmAdd_Bool,
       Ty Pointer_CT$wmAdd_Bool) : (memWriteOut_CT$wmAdd_Bool,MemOut_CT$wmAdd_Bool) (dconPtr_CT$wmAdd_Bool,Pointer_CT$wmAdd_Bool) > [(_74,Pointer_CT$wmAdd_Bool),
                                                                                                                                     (demuxWriteResult_CT$wmAdd_Bool,Pointer_CT$wmAdd_Bool)] */
  logic [1:0] dconPtr_CT$wmAdd_Bool_onehotd;
  always_comb
    if ((memWriteOut_CT$wmAdd_Bool_d[0] && dconPtr_CT$wmAdd_Bool_d[0]))
      unique case (memWriteOut_CT$wmAdd_Bool_d[1:1])
        1'd0: dconPtr_CT$wmAdd_Bool_onehotd = 2'd1;
        1'd1: dconPtr_CT$wmAdd_Bool_onehotd = 2'd2;
        default: dconPtr_CT$wmAdd_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wmAdd_Bool_onehotd = 2'd0;
  assign _74_d = {dconPtr_CT$wmAdd_Bool_d[16:1],
                  dconPtr_CT$wmAdd_Bool_onehotd[0]};
  assign demuxWriteResult_CT$wmAdd_Bool_d = {dconPtr_CT$wmAdd_Bool_d[16:1],
                                             dconPtr_CT$wmAdd_Bool_onehotd[1]};
  assign dconPtr_CT$wmAdd_Bool_r = (| (dconPtr_CT$wmAdd_Bool_onehotd & {demuxWriteResult_CT$wmAdd_Bool_r,
                                                                        _74_r}));
  assign memWriteOut_CT$wmAdd_Bool_r = dconPtr_CT$wmAdd_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Bool,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0,
                                go_1_dummy_write_QTree_Bool_d[0]};
  assign go_1_dummy_write_QTree_Bool_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Bool,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go_2_dummy_write_QTree_Bool_d[0])
          incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go_2_dummy_write_QTree_Bool_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go_2_dummy_write_QTree_Bool_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                                            2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Bool_snk,Word16#) > */
  assign {forkHP1_QTree_Bool_snk_r,
          forkHP1_QTree_Bool_snk_dout} = {forkHP1_QTree_Bool_snk_rout,
                                          forkHP1_QTree_Bool_snk_d};
  
  /* source (Ty Go) : > (\QTree_Bool_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Bool_src,Go) > [(go_1_dummy_write_QTree_Bool,Go),
                                       (go_2_dummy_write_QTree_Bool,Go)] */
  logic [1:0] \\QTree_Bool_src_emitted ;
  logic [1:0] \\QTree_Bool_src_done ;
  assign go_1_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [0]));
  assign go_2_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [1]));
  assign \\QTree_Bool_src_done  = (\\QTree_Bool_src_emitted  | ({go_2_dummy_write_QTree_Bool_d[0],
                                                                 go_1_dummy_write_QTree_Bool_d[0]} & {go_2_dummy_write_QTree_Bool_r,
                                                                                                      go_1_dummy_write_QTree_Bool_r}));
  assign \\QTree_Bool_src_r  = (& \\QTree_Bool_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Bool_src_emitted  <= 2'd0;
    else
      \\QTree_Bool_src_emitted  <= (\\QTree_Bool_src_r  ? 2'd0 :
                                    \\QTree_Bool_src_done );
  
  /* source (Ty QTree_Bool) : > (dummy_write_QTree_Bool,QTree_Bool) */
  
  /* sink (Ty Pointer_QTree_Bool) : (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool) > */
  assign {dummy_write_QTree_Bool_sink_r,
          dummy_write_QTree_Bool_sink_dout} = {dummy_write_QTree_Bool_sink_rout,
                                               dummy_write_QTree_Bool_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Bool_snk,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#),
                                                        (forkHP1_QTree_Boo4,Word16#)] */
  logic [3:0] mergeHP_QTree_Bool_buf_emitted;
  logic [3:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Bool_snk_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                     (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign forkHP1_QTree_Boo4_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[3]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo4_d[0],
                                                                           forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Bool_snk_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo4_r,
                                                                                                       forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Bool_snk_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 4'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Bool) : [(ma8q_1_argbuf,Pointer_QTree_Bool),
                                     (w1sic_1_1_argbuf,Pointer_QTree_Bool),
                                     (w2sid_1_1_argbuf,Pointer_QTree_Bool)] > (readMerge_choice_QTree_Bool,C3) (readMerge_data_QTree_Bool,Pointer_QTree_Bool) */
  logic [2:0] ma8q_1_argbuf_select_d;
  assign ma8q_1_argbuf_select_d = ((| ma8q_1_argbuf_select_q) ? ma8q_1_argbuf_select_q :
                                   (ma8q_1_argbuf_d[0] ? 3'd1 :
                                    (w1sic_1_1_argbuf_d[0] ? 3'd2 :
                                     (w2sid_1_1_argbuf_d[0] ? 3'd4 :
                                      3'd0))));
  logic [2:0] ma8q_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_argbuf_select_q <= 3'd0;
    else
      ma8q_1_argbuf_select_q <= (ma8q_1_argbuf_done ? 3'd0 :
                                 ma8q_1_argbuf_select_d);
  logic [1:0] ma8q_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_argbuf_emit_q <= 2'd0;
    else
      ma8q_1_argbuf_emit_q <= (ma8q_1_argbuf_done ? 2'd0 :
                               ma8q_1_argbuf_emit_d);
  logic [1:0] ma8q_1_argbuf_emit_d;
  assign ma8q_1_argbuf_emit_d = (ma8q_1_argbuf_emit_q | ({readMerge_choice_QTree_Bool_d[0],
                                                          readMerge_data_QTree_Bool_d[0]} & {readMerge_choice_QTree_Bool_r,
                                                                                             readMerge_data_QTree_Bool_r}));
  logic ma8q_1_argbuf_done;
  assign ma8q_1_argbuf_done = (& ma8q_1_argbuf_emit_d);
  assign {w2sid_1_1_argbuf_r,
          w1sic_1_1_argbuf_r,
          ma8q_1_argbuf_r} = (ma8q_1_argbuf_done ? ma8q_1_argbuf_select_d :
                              3'd0);
  assign readMerge_data_QTree_Bool_d = ((ma8q_1_argbuf_select_d[0] && (! ma8q_1_argbuf_emit_q[0])) ? ma8q_1_argbuf_d :
                                        ((ma8q_1_argbuf_select_d[1] && (! ma8q_1_argbuf_emit_q[0])) ? w1sic_1_1_argbuf_d :
                                         ((ma8q_1_argbuf_select_d[2] && (! ma8q_1_argbuf_emit_q[0])) ? w2sid_1_1_argbuf_d :
                                          {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Bool_d = ((ma8q_1_argbuf_select_d[0] && (! ma8q_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((ma8q_1_argbuf_select_d[1] && (! ma8q_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((ma8q_1_argbuf_select_d[2] && (! ma8q_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Bool) : (readMerge_choice_QTree_Bool,C3) (destructReadOut_QTree_Bool,QTree_Bool) > [(readPointer_QTree_Boolma8q_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolw1sic_1_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolw2sid_1_1_argbuf,QTree_Bool)] */
  logic [2:0] destructReadOut_QTree_Bool_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Bool_d[0] && destructReadOut_QTree_Bool_d[0]))
      unique case (readMerge_choice_QTree_Bool_d[2:1])
        2'd0: destructReadOut_QTree_Bool_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Bool_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Bool_onehotd = 3'd4;
        default: destructReadOut_QTree_Bool_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Bool_onehotd = 3'd0;
  assign readPointer_QTree_Boolma8q_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                  destructReadOut_QTree_Bool_onehotd[0]};
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                     destructReadOut_QTree_Bool_onehotd[1]};
  assign readPointer_QTree_Boolw2sid_1_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                     destructReadOut_QTree_Bool_onehotd[2]};
  assign destructReadOut_QTree_Bool_r = (| (destructReadOut_QTree_Bool_onehotd & {readPointer_QTree_Boolw2sid_1_1_argbuf_r,
                                                                                  readPointer_QTree_Boolw1sic_1_1_argbuf_r,
                                                                                  readPointer_QTree_Boolma8q_1_argbuf_r}));
  assign readMerge_choice_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (readMerge_data_QTree_Bool,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {readMerge_data_QTree_Bool_d[16:1],
                                        readMerge_data_QTree_Bool_d[0]};
  assign readMerge_data_QTree_Bool_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(destructReadOut_QTree_Bool,QTree_Bool)] */
  assign destructReadOut_QTree_Bool_d = {memReadOut_QTree_Bool_d[67:2],
                                         memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* mergectrl (Ty C13,
           Ty QTree_Bool) : [(lizzieLet10_1_1_argbuf,QTree_Bool),
                             (lizzieLet12_1_argbuf,QTree_Bool),
                             (lizzieLet14_1_argbuf,QTree_Bool),
                             (lizzieLet15_1_argbuf,QTree_Bool),
                             (lizzieLet17_1_argbuf,QTree_Bool),
                             (lizzieLet23_1_argbuf,QTree_Bool),
                             (lizzieLet28_1_argbuf,QTree_Bool),
                             (lizzieLet3_1_argbuf,QTree_Bool),
                             (lizzieLet4_1_argbuf,QTree_Bool),
                             (lizzieLet5_1_1_argbuf,QTree_Bool),
                             (lizzieLet7_1_1_argbuf,QTree_Bool),
                             (lizzieLet9_1_1_argbuf,QTree_Bool),
                             (dummy_write_QTree_Bool,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C13) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [12:0] lizzieLet10_1_1_argbuf_select_d;
  assign lizzieLet10_1_1_argbuf_select_d = ((| lizzieLet10_1_1_argbuf_select_q) ? lizzieLet10_1_1_argbuf_select_q :
                                            (lizzieLet10_1_1_argbuf_d[0] ? 13'd1 :
                                             (lizzieLet12_1_argbuf_d[0] ? 13'd2 :
                                              (lizzieLet14_1_argbuf_d[0] ? 13'd4 :
                                               (lizzieLet15_1_argbuf_d[0] ? 13'd8 :
                                                (lizzieLet17_1_argbuf_d[0] ? 13'd16 :
                                                 (lizzieLet23_1_argbuf_d[0] ? 13'd32 :
                                                  (lizzieLet28_1_argbuf_d[0] ? 13'd64 :
                                                   (lizzieLet3_1_argbuf_d[0] ? 13'd128 :
                                                    (lizzieLet4_1_argbuf_d[0] ? 13'd256 :
                                                     (lizzieLet5_1_1_argbuf_d[0] ? 13'd512 :
                                                      (lizzieLet7_1_1_argbuf_d[0] ? 13'd1024 :
                                                       (lizzieLet9_1_1_argbuf_d[0] ? 13'd2048 :
                                                        (dummy_write_QTree_Bool_d[0] ? 13'd4096 :
                                                         13'd0))))))))))))));
  logic [12:0] lizzieLet10_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_select_q <= 13'd0;
    else
      lizzieLet10_1_1_argbuf_select_q <= (lizzieLet10_1_1_argbuf_done ? 13'd0 :
                                          lizzieLet10_1_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_1_argbuf_emit_q <= (lizzieLet10_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet10_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_1_argbuf_emit_d;
  assign lizzieLet10_1_1_argbuf_emit_d = (lizzieLet10_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                            writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                                writeMerge_data_QTree_Bool_r}));
  logic lizzieLet10_1_1_argbuf_done;
  assign lizzieLet10_1_1_argbuf_done = (& lizzieLet10_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Bool_r,
          lizzieLet9_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r,
          lizzieLet4_1_argbuf_r,
          lizzieLet3_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = (lizzieLet10_1_1_argbuf_done ? lizzieLet10_1_1_argbuf_select_d :
                                       13'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet10_1_1_argbuf_d :
                                         ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet12_1_argbuf_d :
                                          ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                           ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                            ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                             ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                              ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                               ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet3_1_argbuf_d :
                                                ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet4_1_argbuf_d :
                                                 ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet5_1_1_argbuf_d :
                                                  ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_1_argbuf_d :
                                                   ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_1_argbuf_d :
                                                    ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Bool_d :
                                                     {66'd0, 1'd0})))))))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet10_1_1_argbuf_select_d[0] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C1_13_dc(1'd1) :
                                           ((lizzieLet10_1_1_argbuf_select_d[1] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C2_13_dc(1'd1) :
                                            ((lizzieLet10_1_1_argbuf_select_d[2] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C3_13_dc(1'd1) :
                                             ((lizzieLet10_1_1_argbuf_select_d[3] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C4_13_dc(1'd1) :
                                              ((lizzieLet10_1_1_argbuf_select_d[4] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C5_13_dc(1'd1) :
                                               ((lizzieLet10_1_1_argbuf_select_d[5] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C6_13_dc(1'd1) :
                                                ((lizzieLet10_1_1_argbuf_select_d[6] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C7_13_dc(1'd1) :
                                                 ((lizzieLet10_1_1_argbuf_select_d[7] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C8_13_dc(1'd1) :
                                                  ((lizzieLet10_1_1_argbuf_select_d[8] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C9_13_dc(1'd1) :
                                                   ((lizzieLet10_1_1_argbuf_select_d[9] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C10_13_dc(1'd1) :
                                                    ((lizzieLet10_1_1_argbuf_select_d[10] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C11_13_dc(1'd1) :
                                                     ((lizzieLet10_1_1_argbuf_select_d[11] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C12_13_dc(1'd1) :
                                                      ((lizzieLet10_1_1_argbuf_select_d[12] && (! lizzieLet10_1_1_argbuf_emit_q[1])) ? C13_13_dc(1'd1) :
                                                       {4'd0, 1'd0})))))))))))));
  
  /* demux (Ty C13,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C13) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet12_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet15_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet17_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet23_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet5_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet7_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                       (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool)] */
  logic [12:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[4:1])
        4'd0: demuxWriteResult_QTree_Bool_onehotd = 13'd1;
        4'd1: demuxWriteResult_QTree_Bool_onehotd = 13'd2;
        4'd2: demuxWriteResult_QTree_Bool_onehotd = 13'd4;
        4'd3: demuxWriteResult_QTree_Bool_onehotd = 13'd8;
        4'd4: demuxWriteResult_QTree_Bool_onehotd = 13'd16;
        4'd5: demuxWriteResult_QTree_Bool_onehotd = 13'd32;
        4'd6: demuxWriteResult_QTree_Bool_onehotd = 13'd64;
        4'd7: demuxWriteResult_QTree_Bool_onehotd = 13'd128;
        4'd8: demuxWriteResult_QTree_Bool_onehotd = 13'd256;
        4'd9: demuxWriteResult_QTree_Bool_onehotd = 13'd512;
        4'd10: demuxWriteResult_QTree_Bool_onehotd = 13'd1024;
        4'd11: demuxWriteResult_QTree_Bool_onehotd = 13'd2048;
        4'd12: demuxWriteResult_QTree_Bool_onehotd = 13'd4096;
        default: demuxWriteResult_QTree_Bool_onehotd = 13'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 13'd0;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet12_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet17_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet23_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet3_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[7]};
  assign writeQTree_BoollizzieLet4_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[8]};
  assign writeQTree_BoollizzieLet5_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                   demuxWriteResult_QTree_Bool_onehotd[9]};
  assign writeQTree_BoollizzieLet7_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                   demuxWriteResult_QTree_Bool_onehotd[10]};
  assign writeQTree_BoollizzieLet9_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                   demuxWriteResult_QTree_Bool_onehotd[11]};
  assign dummy_write_QTree_Bool_sink_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                          demuxWriteResult_QTree_Bool_onehotd[12]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {dummy_write_QTree_Bool_sink_r,
                                                                                    writeQTree_BoollizzieLet9_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet7_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet5_1_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet4_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet3_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet28_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet23_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet17_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet15_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet14_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet12_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet10_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo3_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo3_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo4,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo4_d[0]}), forkHP1_QTree_Boo4_d);
  assign {forkHP1_QTree_Boo4_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_73,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _73_d = {dconPtr_QTree_Bool_d[16:1],
                  dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _73_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__6,Go) > (initHP_CTmain_mask_Bool,Word16#) */
  assign initHP_CTmain_mask_Bool_d = {16'd0, go__6_d[0]};
  assign go__6_r = initHP_CTmain_mask_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_mask_Bool1,Go) > (incrHP_CTmain_mask_Bool,Word16#) */
  assign incrHP_CTmain_mask_Bool_d = {16'd1,
                                      incrHP_CTmain_mask_Bool1_d[0]};
  assign incrHP_CTmain_mask_Bool1_r = incrHP_CTmain_mask_Bool_r;
  
  /* merge (Ty Go) : [(go__7,Go),
                 (incrHP_CTmain_mask_Bool2,Go)] > (incrHP_mergeCTmain_mask_Bool,Go) */
  logic [1:0] incrHP_mergeCTmain_mask_Bool_selected;
  logic [1:0] incrHP_mergeCTmain_mask_Bool_select;
  always_comb
    begin
      incrHP_mergeCTmain_mask_Bool_selected = 2'd0;
      if ((| incrHP_mergeCTmain_mask_Bool_select))
        incrHP_mergeCTmain_mask_Bool_selected = incrHP_mergeCTmain_mask_Bool_select;
      else
        if (go__7_d[0]) incrHP_mergeCTmain_mask_Bool_selected[0] = 1'd1;
        else if (incrHP_CTmain_mask_Bool2_d[0])
          incrHP_mergeCTmain_mask_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCTmain_mask_Bool_select <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Bool_select <= (incrHP_mergeCTmain_mask_Bool_r ? 2'd0 :
                                              incrHP_mergeCTmain_mask_Bool_selected);
  always_comb
    if (incrHP_mergeCTmain_mask_Bool_selected[0])
      incrHP_mergeCTmain_mask_Bool_d = go__7_d;
    else if (incrHP_mergeCTmain_mask_Bool_selected[1])
      incrHP_mergeCTmain_mask_Bool_d = incrHP_CTmain_mask_Bool2_d;
    else incrHP_mergeCTmain_mask_Bool_d = 1'd0;
  assign {incrHP_CTmain_mask_Bool2_r,
          go__7_r} = (incrHP_mergeCTmain_mask_Bool_r ? incrHP_mergeCTmain_mask_Bool_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_mask_Bool_buf,Go) > [(incrHP_CTmain_mask_Bool1,Go),
                                                        (incrHP_CTmain_mask_Bool2,Go)] */
  logic [1:0] incrHP_mergeCTmain_mask_Bool_buf_emitted;
  logic [1:0] incrHP_mergeCTmain_mask_Bool_buf_done;
  assign incrHP_CTmain_mask_Bool1_d = (incrHP_mergeCTmain_mask_Bool_buf_d[0] && (! incrHP_mergeCTmain_mask_Bool_buf_emitted[0]));
  assign incrHP_CTmain_mask_Bool2_d = (incrHP_mergeCTmain_mask_Bool_buf_d[0] && (! incrHP_mergeCTmain_mask_Bool_buf_emitted[1]));
  assign incrHP_mergeCTmain_mask_Bool_buf_done = (incrHP_mergeCTmain_mask_Bool_buf_emitted | ({incrHP_CTmain_mask_Bool2_d[0],
                                                                                               incrHP_CTmain_mask_Bool1_d[0]} & {incrHP_CTmain_mask_Bool2_r,
                                                                                                                                 incrHP_CTmain_mask_Bool1_r}));
  assign incrHP_mergeCTmain_mask_Bool_buf_r = (& incrHP_mergeCTmain_mask_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTmain_mask_Bool_buf_emitted <= (incrHP_mergeCTmain_mask_Bool_buf_r ? 2'd0 :
                                                   incrHP_mergeCTmain_mask_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_mask_Bool,Word16#) (forkHP1_CTmain_mask_Bool,Word16#) > (addHP_CTmain_mask_Bool,Word16#) */
  assign addHP_CTmain_mask_Bool_d = {(incrHP_CTmain_mask_Bool_d[16:1] + forkHP1_CTmain_mask_Bool_d[16:1]),
                                     (incrHP_CTmain_mask_Bool_d[0] && forkHP1_CTmain_mask_Bool_d[0])};
  assign {incrHP_CTmain_mask_Bool_r,
          forkHP1_CTmain_mask_Bool_r} = {2 {(addHP_CTmain_mask_Bool_r && addHP_CTmain_mask_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_mask_Bool,Word16#),
                      (addHP_CTmain_mask_Bool,Word16#)] > (mergeHP_CTmain_mask_Bool,Word16#) */
  logic [1:0] mergeHP_CTmain_mask_Bool_selected;
  logic [1:0] mergeHP_CTmain_mask_Bool_select;
  always_comb
    begin
      mergeHP_CTmain_mask_Bool_selected = 2'd0;
      if ((| mergeHP_CTmain_mask_Bool_select))
        mergeHP_CTmain_mask_Bool_selected = mergeHP_CTmain_mask_Bool_select;
      else
        if (initHP_CTmain_mask_Bool_d[0])
          mergeHP_CTmain_mask_Bool_selected[0] = 1'd1;
        else if (addHP_CTmain_mask_Bool_d[0])
          mergeHP_CTmain_mask_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Bool_select <= 2'd0;
    else
      mergeHP_CTmain_mask_Bool_select <= (mergeHP_CTmain_mask_Bool_r ? 2'd0 :
                                          mergeHP_CTmain_mask_Bool_selected);
  always_comb
    if (mergeHP_CTmain_mask_Bool_selected[0])
      mergeHP_CTmain_mask_Bool_d = initHP_CTmain_mask_Bool_d;
    else if (mergeHP_CTmain_mask_Bool_selected[1])
      mergeHP_CTmain_mask_Bool_d = addHP_CTmain_mask_Bool_d;
    else mergeHP_CTmain_mask_Bool_d = {16'd0, 1'd0};
  assign {addHP_CTmain_mask_Bool_r,
          initHP_CTmain_mask_Bool_r} = (mergeHP_CTmain_mask_Bool_r ? mergeHP_CTmain_mask_Bool_selected :
                                        2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_mask_Bool,Go) > (incrHP_mergeCTmain_mask_Bool_buf,Go) */
  Go_t incrHP_mergeCTmain_mask_Bool_bufchan_d;
  logic incrHP_mergeCTmain_mask_Bool_bufchan_r;
  assign incrHP_mergeCTmain_mask_Bool_r = ((! incrHP_mergeCTmain_mask_Bool_bufchan_d[0]) || incrHP_mergeCTmain_mask_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTmain_mask_Bool_r)
        incrHP_mergeCTmain_mask_Bool_bufchan_d <= incrHP_mergeCTmain_mask_Bool_d;
  Go_t incrHP_mergeCTmain_mask_Bool_bufchan_buf;
  assign incrHP_mergeCTmain_mask_Bool_bufchan_r = (! incrHP_mergeCTmain_mask_Bool_bufchan_buf[0]);
  assign incrHP_mergeCTmain_mask_Bool_buf_d = (incrHP_mergeCTmain_mask_Bool_bufchan_buf[0] ? incrHP_mergeCTmain_mask_Bool_bufchan_buf :
                                               incrHP_mergeCTmain_mask_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTmain_mask_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTmain_mask_Bool_buf_r && incrHP_mergeCTmain_mask_Bool_bufchan_buf[0]))
        incrHP_mergeCTmain_mask_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTmain_mask_Bool_buf_r) && (! incrHP_mergeCTmain_mask_Bool_bufchan_buf[0])))
        incrHP_mergeCTmain_mask_Bool_bufchan_buf <= incrHP_mergeCTmain_mask_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_mask_Bool,Word16#) > (mergeHP_CTmain_mask_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_CTmain_mask_Bool_bufchan_d;
  logic mergeHP_CTmain_mask_Bool_bufchan_r;
  assign mergeHP_CTmain_mask_Bool_r = ((! mergeHP_CTmain_mask_Bool_bufchan_d[0]) || mergeHP_CTmain_mask_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTmain_mask_Bool_r)
        mergeHP_CTmain_mask_Bool_bufchan_d <= mergeHP_CTmain_mask_Bool_d;
  \Word16#_t  mergeHP_CTmain_mask_Bool_bufchan_buf;
  assign mergeHP_CTmain_mask_Bool_bufchan_r = (! mergeHP_CTmain_mask_Bool_bufchan_buf[0]);
  assign mergeHP_CTmain_mask_Bool_buf_d = (mergeHP_CTmain_mask_Bool_bufchan_buf[0] ? mergeHP_CTmain_mask_Bool_bufchan_buf :
                                           mergeHP_CTmain_mask_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTmain_mask_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTmain_mask_Bool_buf_r && mergeHP_CTmain_mask_Bool_bufchan_buf[0]))
        mergeHP_CTmain_mask_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTmain_mask_Bool_buf_r) && (! mergeHP_CTmain_mask_Bool_bufchan_buf[0])))
        mergeHP_CTmain_mask_Bool_bufchan_buf <= mergeHP_CTmain_mask_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_mask_Bool_buf,Word16#) > [(forkHP1_CTmain_mask_Bool,Word16#),
                                                              (forkHP1_CTmain_mask_Boo2,Word16#),
                                                              (forkHP1_CTmain_mask_Boo3,Word16#)] */
  logic [2:0] mergeHP_CTmain_mask_Bool_buf_emitted;
  logic [2:0] mergeHP_CTmain_mask_Bool_buf_done;
  assign forkHP1_CTmain_mask_Bool_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[0]))};
  assign forkHP1_CTmain_mask_Boo2_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[1]))};
  assign forkHP1_CTmain_mask_Boo3_d = {mergeHP_CTmain_mask_Bool_buf_d[16:1],
                                       (mergeHP_CTmain_mask_Bool_buf_d[0] && (! mergeHP_CTmain_mask_Bool_buf_emitted[2]))};
  assign mergeHP_CTmain_mask_Bool_buf_done = (mergeHP_CTmain_mask_Bool_buf_emitted | ({forkHP1_CTmain_mask_Boo3_d[0],
                                                                                       forkHP1_CTmain_mask_Boo2_d[0],
                                                                                       forkHP1_CTmain_mask_Bool_d[0]} & {forkHP1_CTmain_mask_Boo3_r,
                                                                                                                         forkHP1_CTmain_mask_Boo2_r,
                                                                                                                         forkHP1_CTmain_mask_Bool_r}));
  assign mergeHP_CTmain_mask_Bool_buf_r = (& mergeHP_CTmain_mask_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTmain_mask_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_CTmain_mask_Bool_buf_emitted <= (mergeHP_CTmain_mask_Bool_buf_r ? 3'd0 :
                                               mergeHP_CTmain_mask_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_mask_Bool) : [(dconReadIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool),
                                         (dconWriteIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool)] > (memMergeChoice_CTmain_mask_Bool,C2) (memMergeIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  logic [1:0] dconReadIn_CTmain_mask_Bool_select_d;
  assign dconReadIn_CTmain_mask_Bool_select_d = ((| dconReadIn_CTmain_mask_Bool_select_q) ? dconReadIn_CTmain_mask_Bool_select_q :
                                                 (dconReadIn_CTmain_mask_Bool_d[0] ? 2'd1 :
                                                  (dconWriteIn_CTmain_mask_Bool_d[0] ? 2'd2 :
                                                   2'd0)));
  logic [1:0] dconReadIn_CTmain_mask_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Bool_select_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Bool_select_q <= (dconReadIn_CTmain_mask_Bool_done ? 2'd0 :
                                               dconReadIn_CTmain_mask_Bool_select_d);
  logic [1:0] dconReadIn_CTmain_mask_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CTmain_mask_Bool_emit_q <= 2'd0;
    else
      dconReadIn_CTmain_mask_Bool_emit_q <= (dconReadIn_CTmain_mask_Bool_done ? 2'd0 :
                                             dconReadIn_CTmain_mask_Bool_emit_d);
  logic [1:0] dconReadIn_CTmain_mask_Bool_emit_d;
  assign dconReadIn_CTmain_mask_Bool_emit_d = (dconReadIn_CTmain_mask_Bool_emit_q | ({memMergeChoice_CTmain_mask_Bool_d[0],
                                                                                      memMergeIn_CTmain_mask_Bool_d[0]} & {memMergeChoice_CTmain_mask_Bool_r,
                                                                                                                           memMergeIn_CTmain_mask_Bool_r}));
  logic dconReadIn_CTmain_mask_Bool_done;
  assign dconReadIn_CTmain_mask_Bool_done = (& dconReadIn_CTmain_mask_Bool_emit_d);
  assign {dconWriteIn_CTmain_mask_Bool_r,
          dconReadIn_CTmain_mask_Bool_r} = (dconReadIn_CTmain_mask_Bool_done ? dconReadIn_CTmain_mask_Bool_select_d :
                                            2'd0);
  assign memMergeIn_CTmain_mask_Bool_d = ((dconReadIn_CTmain_mask_Bool_select_d[0] && (! dconReadIn_CTmain_mask_Bool_emit_q[0])) ? dconReadIn_CTmain_mask_Bool_d :
                                          ((dconReadIn_CTmain_mask_Bool_select_d[1] && (! dconReadIn_CTmain_mask_Bool_emit_q[0])) ? dconWriteIn_CTmain_mask_Bool_d :
                                           {132'd0, 1'd0}));
  assign memMergeChoice_CTmain_mask_Bool_d = ((dconReadIn_CTmain_mask_Bool_select_d[0] && (! dconReadIn_CTmain_mask_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                              ((dconReadIn_CTmain_mask_Bool_select_d[1] && (! dconReadIn_CTmain_mask_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                               {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_mask_Bool,
      Ty MemOut_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool_dbuf,MemIn_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) */
  logic [114:0] memMergeIn_CTmain_mask_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTmain_mask_Bool_dbuf_address;
  logic [114:0] memMergeIn_CTmain_mask_Bool_dbuf_din;
  logic [114:0] memOut_CTmain_mask_Bool_q;
  logic memOut_CTmain_mask_Bool_valid;
  logic memMergeIn_CTmain_mask_Bool_dbuf_we;
  logic memOut_CTmain_mask_Bool_we;
  assign memMergeIn_CTmain_mask_Bool_dbuf_din = memMergeIn_CTmain_mask_Bool_dbuf_d[132:18];
  assign memMergeIn_CTmain_mask_Bool_dbuf_address = memMergeIn_CTmain_mask_Bool_dbuf_d[17:2];
  assign memMergeIn_CTmain_mask_Bool_dbuf_we = (memMergeIn_CTmain_mask_Bool_dbuf_d[1:1] && memMergeIn_CTmain_mask_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTmain_mask_Bool_we <= 1'd0;
        memOut_CTmain_mask_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_CTmain_mask_Bool_we <= memMergeIn_CTmain_mask_Bool_dbuf_we;
        memOut_CTmain_mask_Bool_valid <= memMergeIn_CTmain_mask_Bool_dbuf_d[0];
        if (memMergeIn_CTmain_mask_Bool_dbuf_we)
          begin
            memMergeIn_CTmain_mask_Bool_dbuf_mem[memMergeIn_CTmain_mask_Bool_dbuf_address] <= memMergeIn_CTmain_mask_Bool_dbuf_din;
            memOut_CTmain_mask_Bool_q <= memMergeIn_CTmain_mask_Bool_dbuf_din;
          end
        else
          memOut_CTmain_mask_Bool_q <= memMergeIn_CTmain_mask_Bool_dbuf_mem[memMergeIn_CTmain_mask_Bool_dbuf_address];
      end
  assign memOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_q,
                                      memOut_CTmain_mask_Bool_we,
                                      memOut_CTmain_mask_Bool_valid};
  assign memMergeIn_CTmain_mask_Bool_dbuf_r = ((! memOut_CTmain_mask_Bool_valid) || memOut_CTmain_mask_Bool_r);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_mask_Bool) : (memMergeChoice_CTmain_mask_Bool,C2) (memOut_CTmain_mask_Bool_dbuf,MemOut_CTmain_mask_Bool) > [(memReadOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool),
                                                                                                                                    (memWriteOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool)] */
  logic [1:0] memOut_CTmain_mask_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTmain_mask_Bool_d[0] && memOut_CTmain_mask_Bool_dbuf_d[0]))
      unique case (memMergeChoice_CTmain_mask_Bool_d[1:1])
        1'd0: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd2;
        default: memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTmain_mask_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_dbuf_d[116:1],
                                          memOut_CTmain_mask_Bool_dbuf_onehotd[0]};
  assign memWriteOut_CTmain_mask_Bool_d = {memOut_CTmain_mask_Bool_dbuf_d[116:1],
                                           memOut_CTmain_mask_Bool_dbuf_onehotd[1]};
  assign memOut_CTmain_mask_Bool_dbuf_r = (| (memOut_CTmain_mask_Bool_dbuf_onehotd & {memWriteOut_CTmain_mask_Bool_r,
                                                                                      memReadOut_CTmain_mask_Bool_r}));
  assign memMergeChoice_CTmain_mask_Bool_r = memOut_CTmain_mask_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool_rbuf,MemIn_CTmain_mask_Bool) > (memMergeIn_CTmain_mask_Bool_dbuf,MemIn_CTmain_mask_Bool) */
  assign memMergeIn_CTmain_mask_Bool_rbuf_r = ((! memMergeIn_CTmain_mask_Bool_dbuf_d[0]) || memMergeIn_CTmain_mask_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Bool_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CTmain_mask_Bool_rbuf_r)
        memMergeIn_CTmain_mask_Bool_dbuf_d <= memMergeIn_CTmain_mask_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_CTmain_mask_Bool) : (memMergeIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) > (memMergeIn_CTmain_mask_Bool_rbuf,MemIn_CTmain_mask_Bool) */
  MemIn_CTmain_mask_Bool_t memMergeIn_CTmain_mask_Bool_buf;
  assign memMergeIn_CTmain_mask_Bool_r = (! memMergeIn_CTmain_mask_Bool_buf[0]);
  assign memMergeIn_CTmain_mask_Bool_rbuf_d = (memMergeIn_CTmain_mask_Bool_buf[0] ? memMergeIn_CTmain_mask_Bool_buf :
                                               memMergeIn_CTmain_mask_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTmain_mask_Bool_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CTmain_mask_Bool_rbuf_r && memMergeIn_CTmain_mask_Bool_buf[0]))
        memMergeIn_CTmain_mask_Bool_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CTmain_mask_Bool_rbuf_r) && (! memMergeIn_CTmain_mask_Bool_buf[0])))
        memMergeIn_CTmain_mask_Bool_buf <= memMergeIn_CTmain_mask_Bool_d;
  
  /* dbuf (Ty MemOut_CTmain_mask_Bool) : (memOut_CTmain_mask_Bool_rbuf,MemOut_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool_dbuf,MemOut_CTmain_mask_Bool) */
  assign memOut_CTmain_mask_Bool_rbuf_r = ((! memOut_CTmain_mask_Bool_dbuf_d[0]) || memOut_CTmain_mask_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTmain_mask_Bool_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CTmain_mask_Bool_rbuf_r)
        memOut_CTmain_mask_Bool_dbuf_d <= memOut_CTmain_mask_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_CTmain_mask_Bool) : (memOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) > (memOut_CTmain_mask_Bool_rbuf,MemOut_CTmain_mask_Bool) */
  MemOut_CTmain_mask_Bool_t memOut_CTmain_mask_Bool_buf;
  assign memOut_CTmain_mask_Bool_r = (! memOut_CTmain_mask_Bool_buf[0]);
  assign memOut_CTmain_mask_Bool_rbuf_d = (memOut_CTmain_mask_Bool_buf[0] ? memOut_CTmain_mask_Bool_buf :
                                           memOut_CTmain_mask_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CTmain_mask_Bool_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CTmain_mask_Bool_rbuf_r && memOut_CTmain_mask_Bool_buf[0]))
        memOut_CTmain_mask_Bool_buf <= {116'd0, 1'd0};
      else if (((! memOut_CTmain_mask_Bool_rbuf_r) && (! memOut_CTmain_mask_Bool_buf[0])))
        memOut_CTmain_mask_Bool_buf <= memOut_CTmain_mask_Bool_d;
  
  /* destruct (Ty Pointer_CTmain_mask_Bool,
          Dcon Pointer_CTmain_mask_Bool) : (scfarg_0_1_1_argbuf,Pointer_CTmain_mask_Bool) > [(destructReadIn_CTmain_mask_Bool,Word16#)] */
  assign destructReadIn_CTmain_mask_Bool_d = {scfarg_0_1_1_argbuf_d[16:1],
                                              scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = destructReadIn_CTmain_mask_Bool_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Bool,
      Dcon ReadIn_CTmain_mask_Bool) : [(destructReadIn_CTmain_mask_Bool,Word16#)] > (dconReadIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  assign dconReadIn_CTmain_mask_Bool_d = ReadIn_CTmain_mask_Bool_dc((& {destructReadIn_CTmain_mask_Bool_d[0]}), destructReadIn_CTmain_mask_Bool_d);
  assign {destructReadIn_CTmain_mask_Bool_r} = {1 {(dconReadIn_CTmain_mask_Bool_r && dconReadIn_CTmain_mask_Bool_d[0])}};
  
  /* destruct (Ty MemOut_CTmain_mask_Bool,
          Dcon ReadOut_CTmain_mask_Bool) : (memReadOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) > [(readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf,CTmain_mask_Bool)] */
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d = {memReadOut_CTmain_mask_Bool_d[116:2],
                                                              memReadOut_CTmain_mask_Bool_d[0]};
  assign memReadOut_CTmain_mask_Bool_r = readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTmain_mask_Bool) : [(lizzieLet16_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet18_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet25_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet26_1_argbuf,CTmain_mask_Bool),
                                   (lizzieLet27_1_argbuf,CTmain_mask_Bool)] > (writeMerge_choice_CTmain_mask_Bool,C5) (writeMerge_data_CTmain_mask_Bool,CTmain_mask_Bool) */
  logic [4:0] lizzieLet16_1_argbuf_select_d;
  assign lizzieLet16_1_argbuf_select_d = ((| lizzieLet16_1_argbuf_select_q) ? lizzieLet16_1_argbuf_select_q :
                                          (lizzieLet16_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet18_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet25_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet26_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet27_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet16_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet16_1_argbuf_select_q <= (lizzieLet16_1_argbuf_done ? 5'd0 :
                                        lizzieLet16_1_argbuf_select_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet16_1_argbuf_emit_q <= (lizzieLet16_1_argbuf_done ? 2'd0 :
                                      lizzieLet16_1_argbuf_emit_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_d;
  assign lizzieLet16_1_argbuf_emit_d = (lizzieLet16_1_argbuf_emit_q | ({writeMerge_choice_CTmain_mask_Bool_d[0],
                                                                        writeMerge_data_CTmain_mask_Bool_d[0]} & {writeMerge_choice_CTmain_mask_Bool_r,
                                                                                                                  writeMerge_data_CTmain_mask_Bool_r}));
  logic lizzieLet16_1_argbuf_done;
  assign lizzieLet16_1_argbuf_done = (& lizzieLet16_1_argbuf_emit_d);
  assign {lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet16_1_argbuf_r} = (lizzieLet16_1_argbuf_done ? lizzieLet16_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTmain_mask_Bool_d = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                               ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                                ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                 ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                  ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                                   {115'd0, 1'd0})))));
  assign writeMerge_choice_CTmain_mask_Bool_d = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                 ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                  ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                   ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                    ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                     {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_mask_Bool) : (writeMerge_choice_CTmain_mask_Bool,C5) (demuxWriteResult_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) > [(writeCTmain_mask_BoollizzieLet16_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet18_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet25_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet26_1_argbuf,Pointer_CTmain_mask_Bool),
                                                                                                                                              (writeCTmain_mask_BoollizzieLet27_1_argbuf,Pointer_CTmain_mask_Bool)] */
  logic [4:0] demuxWriteResult_CTmain_mask_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_CTmain_mask_Bool_d[0] && demuxWriteResult_CTmain_mask_Bool_d[0]))
      unique case (writeMerge_choice_CTmain_mask_Bool_d[3:1])
        3'd0: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd16;
        default: demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTmain_mask_Bool_onehotd = 5'd0;
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[0]};
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[1]};
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[2]};
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[3]};
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_d = {demuxWriteResult_CTmain_mask_Bool_d[16:1],
                                                        demuxWriteResult_CTmain_mask_Bool_onehotd[4]};
  assign demuxWriteResult_CTmain_mask_Bool_r = (| (demuxWriteResult_CTmain_mask_Bool_onehotd & {writeCTmain_mask_BoollizzieLet27_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet26_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet25_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet18_1_argbuf_r,
                                                                                                writeCTmain_mask_BoollizzieLet16_1_argbuf_r}));
  assign writeMerge_choice_CTmain_mask_Bool_r = demuxWriteResult_CTmain_mask_Bool_r;
  
  /* dcon (Ty MemIn_CTmain_mask_Bool,
      Dcon WriteIn_CTmain_mask_Bool) : [(forkHP1_CTmain_mask_Boo2,Word16#),
                                        (writeMerge_data_CTmain_mask_Bool,CTmain_mask_Bool)] > (dconWriteIn_CTmain_mask_Bool,MemIn_CTmain_mask_Bool) */
  assign dconWriteIn_CTmain_mask_Bool_d = WriteIn_CTmain_mask_Bool_dc((& {forkHP1_CTmain_mask_Boo2_d[0],
                                                                          writeMerge_data_CTmain_mask_Bool_d[0]}), forkHP1_CTmain_mask_Boo2_d, writeMerge_data_CTmain_mask_Bool_d);
  assign {forkHP1_CTmain_mask_Boo2_r,
          writeMerge_data_CTmain_mask_Bool_r} = {2 {(dconWriteIn_CTmain_mask_Bool_r && dconWriteIn_CTmain_mask_Bool_d[0])}};
  
  /* dcon (Ty Pointer_CTmain_mask_Bool,
      Dcon Pointer_CTmain_mask_Bool) : [(forkHP1_CTmain_mask_Boo3,Word16#)] > (dconPtr_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) */
  assign dconPtr_CTmain_mask_Bool_d = Pointer_CTmain_mask_Bool_dc((& {forkHP1_CTmain_mask_Boo3_d[0]}), forkHP1_CTmain_mask_Boo3_d);
  assign {forkHP1_CTmain_mask_Boo3_r} = {1 {(dconPtr_CTmain_mask_Bool_r && dconPtr_CTmain_mask_Bool_d[0])}};
  
  /* demux (Ty MemOut_CTmain_mask_Bool,
       Ty Pointer_CTmain_mask_Bool) : (memWriteOut_CTmain_mask_Bool,MemOut_CTmain_mask_Bool) (dconPtr_CTmain_mask_Bool,Pointer_CTmain_mask_Bool) > [(_72,Pointer_CTmain_mask_Bool),
                                                                                                                                                    (demuxWriteResult_CTmain_mask_Bool,Pointer_CTmain_mask_Bool)] */
  logic [1:0] dconPtr_CTmain_mask_Bool_onehotd;
  always_comb
    if ((memWriteOut_CTmain_mask_Bool_d[0] && dconPtr_CTmain_mask_Bool_d[0]))
      unique case (memWriteOut_CTmain_mask_Bool_d[1:1])
        1'd0: dconPtr_CTmain_mask_Bool_onehotd = 2'd1;
        1'd1: dconPtr_CTmain_mask_Bool_onehotd = 2'd2;
        default: dconPtr_CTmain_mask_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_CTmain_mask_Bool_onehotd = 2'd0;
  assign _72_d = {dconPtr_CTmain_mask_Bool_d[16:1],
                  dconPtr_CTmain_mask_Bool_onehotd[0]};
  assign demuxWriteResult_CTmain_mask_Bool_d = {dconPtr_CTmain_mask_Bool_d[16:1],
                                                dconPtr_CTmain_mask_Bool_onehotd[1]};
  assign dconPtr_CTmain_mask_Bool_r = (| (dconPtr_CTmain_mask_Bool_onehotd & {demuxWriteResult_CTmain_mask_Bool_r,
                                                                              _72_r}));
  assign memWriteOut_CTmain_mask_Bool_r = dconPtr_CTmain_mask_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_MaskQTree,Go) > (initHP_MaskQTree,Word16#) */
  assign initHP_MaskQTree_d = {16'd0,
                               go_1_dummy_write_MaskQTree_d[0]};
  assign go_1_dummy_write_MaskQTree_r = initHP_MaskQTree_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_MaskQTree1,Go) > (incrHP_MaskQTree,Word16#) */
  assign incrHP_MaskQTree_d = {16'd1, incrHP_MaskQTree1_d[0]};
  assign incrHP_MaskQTree1_r = incrHP_MaskQTree_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_MaskQTree,Go),
                 (incrHP_MaskQTree2,Go)] > (incrHP_mergeMaskQTree,Go) */
  logic [1:0] incrHP_mergeMaskQTree_selected;
  logic [1:0] incrHP_mergeMaskQTree_select;
  always_comb
    begin
      incrHP_mergeMaskQTree_selected = 2'd0;
      if ((| incrHP_mergeMaskQTree_select))
        incrHP_mergeMaskQTree_selected = incrHP_mergeMaskQTree_select;
      else
        if (go_2_dummy_write_MaskQTree_d[0])
          incrHP_mergeMaskQTree_selected[0] = 1'd1;
        else if (incrHP_MaskQTree2_d[0])
          incrHP_mergeMaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_select <= 2'd0;
    else
      incrHP_mergeMaskQTree_select <= (incrHP_mergeMaskQTree_r ? 2'd0 :
                                       incrHP_mergeMaskQTree_selected);
  always_comb
    if (incrHP_mergeMaskQTree_selected[0])
      incrHP_mergeMaskQTree_d = go_2_dummy_write_MaskQTree_d;
    else if (incrHP_mergeMaskQTree_selected[1])
      incrHP_mergeMaskQTree_d = incrHP_MaskQTree2_d;
    else incrHP_mergeMaskQTree_d = 1'd0;
  assign {incrHP_MaskQTree2_r,
          go_2_dummy_write_MaskQTree_r} = (incrHP_mergeMaskQTree_r ? incrHP_mergeMaskQTree_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeMaskQTree_buf,Go) > [(incrHP_MaskQTree1,Go),
                                                 (incrHP_MaskQTree2,Go)] */
  logic [1:0] incrHP_mergeMaskQTree_buf_emitted;
  logic [1:0] incrHP_mergeMaskQTree_buf_done;
  assign incrHP_MaskQTree1_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[0]));
  assign incrHP_MaskQTree2_d = (incrHP_mergeMaskQTree_buf_d[0] && (! incrHP_mergeMaskQTree_buf_emitted[1]));
  assign incrHP_mergeMaskQTree_buf_done = (incrHP_mergeMaskQTree_buf_emitted | ({incrHP_MaskQTree2_d[0],
                                                                                 incrHP_MaskQTree1_d[0]} & {incrHP_MaskQTree2_r,
                                                                                                            incrHP_MaskQTree1_r}));
  assign incrHP_mergeMaskQTree_buf_r = (& incrHP_mergeMaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_buf_emitted <= 2'd0;
    else
      incrHP_mergeMaskQTree_buf_emitted <= (incrHP_mergeMaskQTree_buf_r ? 2'd0 :
                                            incrHP_mergeMaskQTree_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_MaskQTree,Word16#) (forkHP1_MaskQTree,Word16#) > (addHP_MaskQTree,Word16#) */
  assign addHP_MaskQTree_d = {(incrHP_MaskQTree_d[16:1] + forkHP1_MaskQTree_d[16:1]),
                              (incrHP_MaskQTree_d[0] && forkHP1_MaskQTree_d[0])};
  assign {incrHP_MaskQTree_r,
          forkHP1_MaskQTree_r} = {2 {(addHP_MaskQTree_r && addHP_MaskQTree_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_MaskQTree,Word16#),
                      (addHP_MaskQTree,Word16#)] > (mergeHP_MaskQTree,Word16#) */
  logic [1:0] mergeHP_MaskQTree_selected;
  logic [1:0] mergeHP_MaskQTree_select;
  always_comb
    begin
      mergeHP_MaskQTree_selected = 2'd0;
      if ((| mergeHP_MaskQTree_select))
        mergeHP_MaskQTree_selected = mergeHP_MaskQTree_select;
      else
        if (initHP_MaskQTree_d[0]) mergeHP_MaskQTree_selected[0] = 1'd1;
        else if (addHP_MaskQTree_d[0])
          mergeHP_MaskQTree_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_select <= 2'd0;
    else
      mergeHP_MaskQTree_select <= (mergeHP_MaskQTree_r ? 2'd0 :
                                   mergeHP_MaskQTree_selected);
  always_comb
    if (mergeHP_MaskQTree_selected[0])
      mergeHP_MaskQTree_d = initHP_MaskQTree_d;
    else if (mergeHP_MaskQTree_selected[1])
      mergeHP_MaskQTree_d = addHP_MaskQTree_d;
    else mergeHP_MaskQTree_d = {16'd0, 1'd0};
  assign {addHP_MaskQTree_r,
          initHP_MaskQTree_r} = (mergeHP_MaskQTree_r ? mergeHP_MaskQTree_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeMaskQTree,Go) > (incrHP_mergeMaskQTree_buf,Go) */
  Go_t incrHP_mergeMaskQTree_bufchan_d;
  logic incrHP_mergeMaskQTree_bufchan_r;
  assign incrHP_mergeMaskQTree_r = ((! incrHP_mergeMaskQTree_bufchan_d[0]) || incrHP_mergeMaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeMaskQTree_r)
        incrHP_mergeMaskQTree_bufchan_d <= incrHP_mergeMaskQTree_d;
  Go_t incrHP_mergeMaskQTree_bufchan_buf;
  assign incrHP_mergeMaskQTree_bufchan_r = (! incrHP_mergeMaskQTree_bufchan_buf[0]);
  assign incrHP_mergeMaskQTree_buf_d = (incrHP_mergeMaskQTree_bufchan_buf[0] ? incrHP_mergeMaskQTree_bufchan_buf :
                                        incrHP_mergeMaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeMaskQTree_buf_r && incrHP_mergeMaskQTree_bufchan_buf[0]))
        incrHP_mergeMaskQTree_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeMaskQTree_buf_r) && (! incrHP_mergeMaskQTree_bufchan_buf[0])))
        incrHP_mergeMaskQTree_bufchan_buf <= incrHP_mergeMaskQTree_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_MaskQTree,Word16#) > (mergeHP_MaskQTree_buf,Word16#) */
  \Word16#_t  mergeHP_MaskQTree_bufchan_d;
  logic mergeHP_MaskQTree_bufchan_r;
  assign mergeHP_MaskQTree_r = ((! mergeHP_MaskQTree_bufchan_d[0]) || mergeHP_MaskQTree_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_MaskQTree_r)
        mergeHP_MaskQTree_bufchan_d <= mergeHP_MaskQTree_d;
  \Word16#_t  mergeHP_MaskQTree_bufchan_buf;
  assign mergeHP_MaskQTree_bufchan_r = (! mergeHP_MaskQTree_bufchan_buf[0]);
  assign mergeHP_MaskQTree_buf_d = (mergeHP_MaskQTree_bufchan_buf[0] ? mergeHP_MaskQTree_bufchan_buf :
                                    mergeHP_MaskQTree_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_MaskQTree_buf_r && mergeHP_MaskQTree_bufchan_buf[0]))
        mergeHP_MaskQTree_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_MaskQTree_buf_r) && (! mergeHP_MaskQTree_bufchan_buf[0])))
        mergeHP_MaskQTree_bufchan_buf <= mergeHP_MaskQTree_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_MaskQTree_snk,Word16#) > */
  assign {forkHP1_MaskQTree_snk_r,
          forkHP1_MaskQTree_snk_dout} = {forkHP1_MaskQTree_snk_rout,
                                         forkHP1_MaskQTree_snk_d};
  
  /* source (Ty Go) : > (\MaskQTree_src,Go) */
  
  /* fork (Ty Go) : (\MaskQTree_src,Go) > [(go_1_dummy_write_MaskQTree,Go),
                                      (go_2_dummy_write_MaskQTree,Go)] */
  logic [1:0] \\MaskQTree_src_emitted ;
  logic [1:0] \\MaskQTree_src_done ;
  assign go_1_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [0]));
  assign go_2_dummy_write_MaskQTree_d = (\\MaskQTree_src_d [0] && (! \\MaskQTree_src_emitted [1]));
  assign \\MaskQTree_src_done  = (\\MaskQTree_src_emitted  | ({go_2_dummy_write_MaskQTree_d[0],
                                                               go_1_dummy_write_MaskQTree_d[0]} & {go_2_dummy_write_MaskQTree_r,
                                                                                                   go_1_dummy_write_MaskQTree_r}));
  assign \\MaskQTree_src_r  = (& \\MaskQTree_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\MaskQTree_src_emitted  <= 2'd0;
    else
      \\MaskQTree_src_emitted  <= (\\MaskQTree_src_r  ? 2'd0 :
                                   \\MaskQTree_src_done );
  
  /* source (Ty MaskQTree) : > (dummy_write_MaskQTree,MaskQTree) */
  
  /* sink (Ty Pointer_MaskQTree) : (dummy_write_MaskQTree_sink,Pointer_MaskQTree) > */
  assign {dummy_write_MaskQTree_sink_r,
          dummy_write_MaskQTree_sink_dout} = {dummy_write_MaskQTree_sink_rout,
                                              dummy_write_MaskQTree_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_MaskQTree_buf,Word16#) > [(forkHP1_MaskQTree,Word16#),
                                                       (forkHP1_MaskQTree_snk,Word16#),
                                                       (forkHP1_MaskQTre3,Word16#),
                                                       (forkHP1_MaskQTre4,Word16#)] */
  logic [3:0] mergeHP_MaskQTree_buf_emitted;
  logic [3:0] mergeHP_MaskQTree_buf_done;
  assign forkHP1_MaskQTree_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[0]))};
  assign forkHP1_MaskQTree_snk_d = {mergeHP_MaskQTree_buf_d[16:1],
                                    (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[1]))};
  assign forkHP1_MaskQTre3_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[2]))};
  assign forkHP1_MaskQTre4_d = {mergeHP_MaskQTree_buf_d[16:1],
                                (mergeHP_MaskQTree_buf_d[0] && (! mergeHP_MaskQTree_buf_emitted[3]))};
  assign mergeHP_MaskQTree_buf_done = (mergeHP_MaskQTree_buf_emitted | ({forkHP1_MaskQTre4_d[0],
                                                                         forkHP1_MaskQTre3_d[0],
                                                                         forkHP1_MaskQTree_snk_d[0],
                                                                         forkHP1_MaskQTree_d[0]} & {forkHP1_MaskQTre4_r,
                                                                                                    forkHP1_MaskQTre3_r,
                                                                                                    forkHP1_MaskQTree_snk_r,
                                                                                                    forkHP1_MaskQTree_r}));
  assign mergeHP_MaskQTree_buf_r = (& mergeHP_MaskQTree_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_MaskQTree_buf_emitted <= 4'd0;
    else
      mergeHP_MaskQTree_buf_emitted <= (mergeHP_MaskQTree_buf_r ? 4'd0 :
                                        mergeHP_MaskQTree_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_MaskQTree) : [(dconReadIn_MaskQTree,MemIn_MaskQTree),
                                  (dconWriteIn_MaskQTree,MemIn_MaskQTree)] > (memMergeChoice_MaskQTree,C2) (memMergeIn_MaskQTree,MemIn_MaskQTree) */
  logic [1:0] dconReadIn_MaskQTree_select_d;
  assign dconReadIn_MaskQTree_select_d = ((| dconReadIn_MaskQTree_select_q) ? dconReadIn_MaskQTree_select_q :
                                          (dconReadIn_MaskQTree_d[0] ? 2'd1 :
                                           (dconWriteIn_MaskQTree_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_MaskQTree_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_select_q <= 2'd0;
    else
      dconReadIn_MaskQTree_select_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                        dconReadIn_MaskQTree_select_d);
  logic [1:0] dconReadIn_MaskQTree_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_MaskQTree_emit_q <= 2'd0;
    else
      dconReadIn_MaskQTree_emit_q <= (dconReadIn_MaskQTree_done ? 2'd0 :
                                      dconReadIn_MaskQTree_emit_d);
  logic [1:0] dconReadIn_MaskQTree_emit_d;
  assign dconReadIn_MaskQTree_emit_d = (dconReadIn_MaskQTree_emit_q | ({memMergeChoice_MaskQTree_d[0],
                                                                        memMergeIn_MaskQTree_d[0]} & {memMergeChoice_MaskQTree_r,
                                                                                                      memMergeIn_MaskQTree_r}));
  logic dconReadIn_MaskQTree_done;
  assign dconReadIn_MaskQTree_done = (& dconReadIn_MaskQTree_emit_d);
  assign {dconWriteIn_MaskQTree_r,
          dconReadIn_MaskQTree_r} = (dconReadIn_MaskQTree_done ? dconReadIn_MaskQTree_select_d :
                                     2'd0);
  assign memMergeIn_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconReadIn_MaskQTree_d :
                                   ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[0])) ? dconWriteIn_MaskQTree_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_MaskQTree_d = ((dconReadIn_MaskQTree_select_d[0] && (! dconReadIn_MaskQTree_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_MaskQTree_select_d[1] && (! dconReadIn_MaskQTree_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_MaskQTree,
      Ty MemOut_MaskQTree) : (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) > (memOut_MaskQTree,MemOut_MaskQTree) */
  logic [65:0] memMergeIn_MaskQTree_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_MaskQTree_dbuf_address;
  logic [65:0] memMergeIn_MaskQTree_dbuf_din;
  logic [65:0] memOut_MaskQTree_q;
  logic memOut_MaskQTree_valid;
  logic memMergeIn_MaskQTree_dbuf_we;
  logic memOut_MaskQTree_we;
  assign memMergeIn_MaskQTree_dbuf_din = memMergeIn_MaskQTree_dbuf_d[83:18];
  assign memMergeIn_MaskQTree_dbuf_address = memMergeIn_MaskQTree_dbuf_d[17:2];
  assign memMergeIn_MaskQTree_dbuf_we = (memMergeIn_MaskQTree_dbuf_d[1:1] && memMergeIn_MaskQTree_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_MaskQTree_we <= 1'd0;
        memOut_MaskQTree_valid <= 1'd0;
      end
    else
      begin
        memOut_MaskQTree_we <= memMergeIn_MaskQTree_dbuf_we;
        memOut_MaskQTree_valid <= memMergeIn_MaskQTree_dbuf_d[0];
        if (memMergeIn_MaskQTree_dbuf_we)
          begin
            memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address] <= memMergeIn_MaskQTree_dbuf_din;
            memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_din;
          end
        else
          memOut_MaskQTree_q <= memMergeIn_MaskQTree_dbuf_mem[memMergeIn_MaskQTree_dbuf_address];
      end
  assign memOut_MaskQTree_d = {memOut_MaskQTree_q,
                               memOut_MaskQTree_we,
                               memOut_MaskQTree_valid};
  assign memMergeIn_MaskQTree_dbuf_r = ((! memOut_MaskQTree_valid) || memOut_MaskQTree_r);
  
  /* demux (Ty C2,
       Ty MemOut_MaskQTree) : (memMergeChoice_MaskQTree,C2) (memOut_MaskQTree_dbuf,MemOut_MaskQTree) > [(memReadOut_MaskQTree,MemOut_MaskQTree),
                                                                                                        (memWriteOut_MaskQTree,MemOut_MaskQTree)] */
  logic [1:0] memOut_MaskQTree_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_MaskQTree_d[0] && memOut_MaskQTree_dbuf_d[0]))
      unique case (memMergeChoice_MaskQTree_d[1:1])
        1'd0: memOut_MaskQTree_dbuf_onehotd = 2'd1;
        1'd1: memOut_MaskQTree_dbuf_onehotd = 2'd2;
        default: memOut_MaskQTree_dbuf_onehotd = 2'd0;
      endcase
    else memOut_MaskQTree_dbuf_onehotd = 2'd0;
  assign memReadOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                   memOut_MaskQTree_dbuf_onehotd[0]};
  assign memWriteOut_MaskQTree_d = {memOut_MaskQTree_dbuf_d[67:1],
                                    memOut_MaskQTree_dbuf_onehotd[1]};
  assign memOut_MaskQTree_dbuf_r = (| (memOut_MaskQTree_dbuf_onehotd & {memWriteOut_MaskQTree_r,
                                                                        memReadOut_MaskQTree_r}));
  assign memMergeChoice_MaskQTree_r = memOut_MaskQTree_dbuf_r;
  
  /* dbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) > (memMergeIn_MaskQTree_dbuf,MemIn_MaskQTree) */
  assign memMergeIn_MaskQTree_rbuf_r = ((! memMergeIn_MaskQTree_dbuf_d[0]) || memMergeIn_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_MaskQTree_rbuf_r)
        memMergeIn_MaskQTree_dbuf_d <= memMergeIn_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemIn_MaskQTree) : (memMergeIn_MaskQTree,MemIn_MaskQTree) > (memMergeIn_MaskQTree_rbuf,MemIn_MaskQTree) */
  MemIn_MaskQTree_t memMergeIn_MaskQTree_buf;
  assign memMergeIn_MaskQTree_r = (! memMergeIn_MaskQTree_buf[0]);
  assign memMergeIn_MaskQTree_rbuf_d = (memMergeIn_MaskQTree_buf[0] ? memMergeIn_MaskQTree_buf :
                                        memMergeIn_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_MaskQTree_rbuf_r && memMergeIn_MaskQTree_buf[0]))
        memMergeIn_MaskQTree_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_MaskQTree_rbuf_r) && (! memMergeIn_MaskQTree_buf[0])))
        memMergeIn_MaskQTree_buf <= memMergeIn_MaskQTree_d;
  
  /* dbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree_rbuf,MemOut_MaskQTree) > (memOut_MaskQTree_dbuf,MemOut_MaskQTree) */
  assign memOut_MaskQTree_rbuf_r = ((! memOut_MaskQTree_dbuf_d[0]) || memOut_MaskQTree_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_MaskQTree_rbuf_r)
        memOut_MaskQTree_dbuf_d <= memOut_MaskQTree_rbuf_d;
  
  /* rbuf (Ty MemOut_MaskQTree) : (memOut_MaskQTree,MemOut_MaskQTree) > (memOut_MaskQTree_rbuf,MemOut_MaskQTree) */
  MemOut_MaskQTree_t memOut_MaskQTree_buf;
  assign memOut_MaskQTree_r = (! memOut_MaskQTree_buf[0]);
  assign memOut_MaskQTree_rbuf_d = (memOut_MaskQTree_buf[0] ? memOut_MaskQTree_buf :
                                    memOut_MaskQTree_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_MaskQTree_buf <= {67'd0, 1'd0};
    else
      if ((memOut_MaskQTree_rbuf_r && memOut_MaskQTree_buf[0]))
        memOut_MaskQTree_buf <= {67'd0, 1'd0};
      else if (((! memOut_MaskQTree_rbuf_r) && (! memOut_MaskQTree_buf[0])))
        memOut_MaskQTree_buf <= memOut_MaskQTree_d;
  
  /* destruct (Ty Pointer_MaskQTree,
          Dcon Pointer_MaskQTree) : (mska8r_1_argbuf,Pointer_MaskQTree) > [(destructReadIn_MaskQTree,Word16#)] */
  assign destructReadIn_MaskQTree_d = {mska8r_1_argbuf_d[16:1],
                                       mska8r_1_argbuf_d[0]};
  assign mska8r_1_argbuf_r = destructReadIn_MaskQTree_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon ReadIn_MaskQTree) : [(destructReadIn_MaskQTree,Word16#)] > (dconReadIn_MaskQTree,MemIn_MaskQTree) */
  assign dconReadIn_MaskQTree_d = ReadIn_MaskQTree_dc((& {destructReadIn_MaskQTree_d[0]}), destructReadIn_MaskQTree_d);
  assign {destructReadIn_MaskQTree_r} = {1 {(dconReadIn_MaskQTree_r && dconReadIn_MaskQTree_d[0])}};
  
  /* destruct (Ty MemOut_MaskQTree,
          Dcon ReadOut_MaskQTree) : (memReadOut_MaskQTree,MemOut_MaskQTree) > [(readPointer_MaskQTreemska8r_1_argbuf,MaskQTree)] */
  assign readPointer_MaskQTreemska8r_1_argbuf_d = {memReadOut_MaskQTree_d[67:2],
                                                   memReadOut_MaskQTree_d[0]};
  assign memReadOut_MaskQTree_r = readPointer_MaskQTreemska8r_1_argbuf_r;
  
  /* dcon (Ty MemIn_MaskQTree,
      Dcon WriteIn_MaskQTree) : [(forkHP1_MaskQTre3,Word16#),
                                 (dummy_write_MaskQTree,MaskQTree)] > (dconWriteIn_MaskQTree,MemIn_MaskQTree) */
  assign dconWriteIn_MaskQTree_d = WriteIn_MaskQTree_dc((& {forkHP1_MaskQTre3_d[0],
                                                            dummy_write_MaskQTree_d[0]}), forkHP1_MaskQTre3_d, dummy_write_MaskQTree_d);
  assign {forkHP1_MaskQTre3_r,
          dummy_write_MaskQTree_r} = {2 {(dconWriteIn_MaskQTree_r && dconWriteIn_MaskQTree_d[0])}};
  
  /* dcon (Ty Pointer_MaskQTree,
      Dcon Pointer_MaskQTree) : [(forkHP1_MaskQTre4,Word16#)] > (dconPtr_MaskQTree,Pointer_MaskQTree) */
  assign dconPtr_MaskQTree_d = Pointer_MaskQTree_dc((& {forkHP1_MaskQTre4_d[0]}), forkHP1_MaskQTre4_d);
  assign {forkHP1_MaskQTre4_r} = {1 {(dconPtr_MaskQTree_r && dconPtr_MaskQTree_d[0])}};
  
  /* demux (Ty MemOut_MaskQTree,
       Ty Pointer_MaskQTree) : (memWriteOut_MaskQTree,MemOut_MaskQTree) (dconPtr_MaskQTree,Pointer_MaskQTree) > [(_71,Pointer_MaskQTree),
                                                                                                                 (dummy_write_MaskQTree_sink,Pointer_MaskQTree)] */
  logic [1:0] dconPtr_MaskQTree_onehotd;
  always_comb
    if ((memWriteOut_MaskQTree_d[0] && dconPtr_MaskQTree_d[0]))
      unique case (memWriteOut_MaskQTree_d[1:1])
        1'd0: dconPtr_MaskQTree_onehotd = 2'd1;
        1'd1: dconPtr_MaskQTree_onehotd = 2'd2;
        default: dconPtr_MaskQTree_onehotd = 2'd0;
      endcase
    else dconPtr_MaskQTree_onehotd = 2'd0;
  assign _71_d = {dconPtr_MaskQTree_d[16:1],
                  dconPtr_MaskQTree_onehotd[0]};
  assign dummy_write_MaskQTree_sink_d = {dconPtr_MaskQTree_d[16:1],
                                         dconPtr_MaskQTree_onehotd[1]};
  assign dconPtr_MaskQTree_r = (| (dconPtr_MaskQTree_onehotd & {dummy_write_MaskQTree_sink_r,
                                                                _71_r}));
  assign memWriteOut_MaskQTree_r = dconPtr_MaskQTree_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_MaskQTree) : > (m1a92_0,Pointer_MaskQTree) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m2a93_1,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m3a94_2,Pointer_QTree_Bool) */
  
  /* destruct (Ty TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) > [($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2,Go),
                                                                                                                                                                                                                                                   ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                   ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                   ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid,Pointer_QTree_Bool)] */
  logic [3:0] \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted ;
  logic [3:0] \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_d  = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [0]));
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_d  = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [1]));
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_d  = {\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [16:1],
                                                                                                     (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [2]))};
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_d  = {\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [32:17],
                                                                                                     (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted [3]))};
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done  = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  | ({\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_d [0],
                                                                                                                                                                                                     \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_d [0],
                                                                                                                                                                                                     \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_d [0],
                                                                                                                                                                                                     \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_d [0]} & {\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_r ,
                                                                                                                                                                                                                                                                                                    \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_r ,
                                                                                                                                                                                                                                                                                                    \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_r ,
                                                                                                                                                                                                                                                                                                    \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_r }));
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  = (& \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  <= 4'd0;
    else
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted  <= (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  ? 4'd0 :
                                                                                                      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done );
  
  /* fork (Ty Go) : ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2,Go) > [(go_2_1,Go),
                                                                                                           (go_2_2,Go)] */
  logic [1:0] \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted ;
  logic [1:0] \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_done ;
  assign go_2_1_d = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted [0]));
  assign go_2_2_d = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_d [0] && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted [1]));
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_done  = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted  | ({go_2_2_d[0],
                                                                                                                                                                                                         go_2_1_d[0]} & {go_2_2_r,
                                                                                                                                                                                                                         go_2_1_r}));
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_r  = (& \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted  <= 2'd0;
    else
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_emitted  <= (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_r  ? 2'd0 :
                                                                                                        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_2_done );
  
  /* buf (Ty Pointer_QTree_Bool) : ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic,Pointer_QTree_Bool) > (w1sic_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_r ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_r  = ((! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d [0]) || \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d  <= {16'd0,
                                                                                                           1'd0};
    else
      if (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_r )
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_d ;
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_r  = (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf [0]);
  assign w1sic_1_argbuf_d = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf [0] ? \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf  :
                             \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf  <= {16'd0,
                                                                                                             1'd0};
    else
      if ((w1sic_1_argbuf_r && \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf [0]))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf  <= {16'd0,
                                                                                                               1'd0};
      else if (((! w1sic_1_argbuf_r) && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf [0])))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_buf  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw1sic_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid,Pointer_QTree_Bool) > (w2sid_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_r ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_r  = ((! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d [0]) || \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d  <= {16'd0,
                                                                                                           1'd0};
    else
      if (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_r )
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_d ;
  Pointer_QTree_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_r  = (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf [0]);
  assign w2sid_1_argbuf_d = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf [0] ? \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf  :
                             \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf  <= {16'd0,
                                                                                                             1'd0};
    else
      if ((w2sid_1_argbuf_r && \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf [0]))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf  <= {16'd0,
                                                                                                               1'd0};
      else if (((! w2sid_1_argbuf_r) && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf [0])))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_buf  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolw2sid_bufchan_d ;
  
  /* buf (Ty MyDTBool_Bool_Bool) : ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib,MyDTBool_Bool_Bool) > (wsib_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d ;
  logic \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_r ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_r  = ((! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d [0]) || \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d  <= 1'd0;
    else
      if (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_r )
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_d ;
  MyDTBool_Bool_Bool_t \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf ;
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_r  = (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf [0]);
  assign wsib_1_argbuf_d = (\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf [0] ? \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf  :
                            \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf  <= 1'd0;
    else
      if ((wsib_1_argbuf_r && \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf [0]))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf  <= 1'd0;
      else if (((! wsib_1_argbuf_r) && (! \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf [0])))
        \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_buf  <= \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolwsib_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : ($wmAdd_Bool_resbuf,Pointer_QTree_Bool) > (es_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \$wmAdd_Bool_resbuf_bufchan_d ;
  logic \$wmAdd_Bool_resbuf_bufchan_r ;
  assign \$wmAdd_Bool_resbuf_r  = ((! \$wmAdd_Bool_resbuf_bufchan_d [0]) || \$wmAdd_Bool_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Bool_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\$wmAdd_Bool_resbuf_r )
        \$wmAdd_Bool_resbuf_bufchan_d  <= \$wmAdd_Bool_resbuf_d ;
  Pointer_QTree_Bool_t \$wmAdd_Bool_resbuf_bufchan_buf ;
  assign \$wmAdd_Bool_resbuf_bufchan_r  = (! \$wmAdd_Bool_resbuf_bufchan_buf [0]);
  assign es_0_1_argbuf_d = (\$wmAdd_Bool_resbuf_bufchan_buf [0] ? \$wmAdd_Bool_resbuf_bufchan_buf  :
                            \$wmAdd_Bool_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wmAdd_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && \$wmAdd_Bool_resbuf_bufchan_buf [0]))
        \$wmAdd_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! \$wmAdd_Bool_resbuf_bufchan_buf [0])))
        \$wmAdd_Bool_resbuf_bufchan_buf  <= \$wmAdd_Bool_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
          Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) > [(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0,MyDTBool_Bool_Bool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1,MyBool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done;
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[1:1],
                                                                                      (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[2:2],
                                                                                      (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[3]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted | ({applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]} & {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r ? 4'd0 :
                                                                                        applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool_Bool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0,MyDTBool_Bool_Bool) > [(arg0_1,MyDTBool_Bool_Bool),
                                                                                                                               (arg0_2,MyDTBool_Bool_Bool),
                                                                                                                               (arg0_3,MyDTBool_Bool_Bool),
                                                                                                                               (arg0_4,MyDTBool_Bool_Bool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_done;
  assign arg0_1_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted[0]));
  assign arg0_2_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted[1]));
  assign arg0_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted[2]));
  assign arg0_4_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted[3]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted | ({arg0_4_d[0],
                                                                                                                                                                             arg0_3_d[0],
                                                                                                                                                                             arg0_2_d[0],
                                                                                                                                                                             arg0_1_d[0]} & {arg0_4_r,
                                                                                                                                                                                             arg0_3_r,
                                                                                                                                                                                             arg0_2_r,
                                                                                                                                                                                             arg0_1_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_r ? 4'd0 :
                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(applyfnBool_Bool_Bool_5_resbuf,MyBool)] > (es_0_1_1QVal_Bool,QTree_Bool) */
  assign es_0_1_1QVal_Bool_d = QVal_Bool_dc((& {applyfnBool_Bool_Bool_5_resbuf_d[0]}), applyfnBool_Bool_Bool_5_resbuf_d);
  assign {applyfnBool_Bool_Bool_5_resbuf_r} = {1 {(es_0_1_1QVal_Bool_r && es_0_1_1QVal_Bool_d[0])}};
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_1,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1,MyBool) > [(arg0_1Dcon_||,MyBool)] */
  assign \arg0_1Dcon_||_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d[1:1],
                              (arg0_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_r = (\arg0_1Dcon_||_r  && (arg0_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d[0]));
  assign arg0_1_r = (\arg0_1Dcon_||_r  && (arg0_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_d[0]));
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_2,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool) > [(arg0_2Dcon_||,MyBool)] */
  assign \arg0_2Dcon_||_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[1:1],
                              (arg0_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r = (\arg0_2Dcon_||_r  && (arg0_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  assign arg0_2_r = (\arg0_2Dcon_||_r  && (arg0_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  
  /* fork (Ty MyBool) : (arg0_2Dcon_||,MyBool) > [(arg0_2Dcon_||_1,MyBool),
                                             (arg0_2Dcon_||_2,MyBool),
                                             (arg0_2Dcon_||_3,MyBool)] */
  logic [2:0] \arg0_2Dcon_||_emitted ;
  logic [2:0] \arg0_2Dcon_||_done ;
  assign \arg0_2Dcon_||_1_d  = {\arg0_2Dcon_||_d [1:1],
                                (\arg0_2Dcon_||_d [0] && (! \arg0_2Dcon_||_emitted [0]))};
  assign \arg0_2Dcon_||_2_d  = {\arg0_2Dcon_||_d [1:1],
                                (\arg0_2Dcon_||_d [0] && (! \arg0_2Dcon_||_emitted [1]))};
  assign \arg0_2Dcon_||_3_d  = {\arg0_2Dcon_||_d [1:1],
                                (\arg0_2Dcon_||_d [0] && (! \arg0_2Dcon_||_emitted [2]))};
  assign \arg0_2Dcon_||_done  = (\arg0_2Dcon_||_emitted  | ({\arg0_2Dcon_||_3_d [0],
                                                             \arg0_2Dcon_||_2_d [0],
                                                             \arg0_2Dcon_||_1_d [0]} & {\arg0_2Dcon_||_3_r ,
                                                                                        \arg0_2Dcon_||_2_r ,
                                                                                        \arg0_2Dcon_||_1_r }));
  assign \arg0_2Dcon_||_r  = (& \arg0_2Dcon_||_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2Dcon_||_emitted  <= 3'd0;
    else
      \arg0_2Dcon_||_emitted  <= (\arg0_2Dcon_||_r  ? 3'd0 :
                                  \arg0_2Dcon_||_done );
  
  /* demux (Ty MyBool,
       Ty MyBool) : (arg0_2Dcon_||_1,MyBool) (arg0_1Dcon_||,MyBool) > [(arg0_2Dcon_||_1MyFalse,MyBool),
                                                                       (_70,MyBool)] */
  logic [1:0] \arg0_1Dcon_||_onehotd ;
  always_comb
    if ((\arg0_2Dcon_||_1_d [0] && \arg0_1Dcon_||_d [0]))
      unique case (\arg0_2Dcon_||_1_d [1:1])
        1'd0: \arg0_1Dcon_||_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_||_onehotd  = 2'd2;
        default: \arg0_1Dcon_||_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_||_onehotd  = 2'd0;
  assign \arg0_2Dcon_||_1MyFalse_d  = {\arg0_1Dcon_||_d [1:1],
                                       \arg0_1Dcon_||_onehotd [0]};
  assign _70_d = {\arg0_1Dcon_||_d [1:1],
                  \arg0_1Dcon_||_onehotd [1]};
  assign \arg0_1Dcon_||_r  = (| (\arg0_1Dcon_||_onehotd  & {_70_r,
                                                            \arg0_2Dcon_||_1MyFalse_r }));
  assign \arg0_2Dcon_||_1_r  = \arg0_1Dcon_||_r ;
  
  /* buf (Ty MyBool) : (arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux,MyBool) > (applyfnBool_Bool_Bool_5_resbuf,MyBool) */
  MyBool_t \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d ;
  logic \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_r ;
  assign \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_r  = ((! \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d [0]) || \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d  <= {1'd0,
                                                                                    1'd0};
    else
      if (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_r )
        \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d  <= \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_d ;
  MyBool_t \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf ;
  assign \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_r  = (! \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf [0]);
  assign applyfnBool_Bool_Bool_5_resbuf_d = (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf [0] ? \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf  :
                                             \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf  <= {1'd0,
                                                                                      1'd0};
    else
      if ((applyfnBool_Bool_Bool_5_resbuf_r && \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf [0]))
        \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf  <= {1'd0,
                                                                                        1'd0};
      else if (((! applyfnBool_Bool_Bool_5_resbuf_r) && (! \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf [0])))
        \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_buf  <= \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_bufchan_d ;
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_2Dcon_||_2,MyBool) (arg0_3Dcon_||,Go) > [(_69,Go),
                                                               (arg0_2Dcon_||_2MyTrue,Go)] */
  logic [1:0] \arg0_3Dcon_||_onehotd ;
  always_comb
    if ((\arg0_2Dcon_||_2_d [0] && \arg0_3Dcon_||_d [0]))
      unique case (\arg0_2Dcon_||_2_d [1:1])
        1'd0: \arg0_3Dcon_||_onehotd  = 2'd1;
        1'd1: \arg0_3Dcon_||_onehotd  = 2'd2;
        default: \arg0_3Dcon_||_onehotd  = 2'd0;
      endcase
    else \arg0_3Dcon_||_onehotd  = 2'd0;
  assign _69_d = \arg0_3Dcon_||_onehotd [0];
  assign \arg0_2Dcon_||_2MyTrue_d  = \arg0_3Dcon_||_onehotd [1];
  assign \arg0_3Dcon_||_r  = (| (\arg0_3Dcon_||_onehotd  & {\arg0_2Dcon_||_2MyTrue_r ,
                                                            _69_r}));
  assign \arg0_2Dcon_||_2_r  = \arg0_3Dcon_||_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(arg0_2Dcon_||_2MyTrue,Go)] > (arg0_2Dcon_||_2MyTrue_1MyTrue,MyBool) */
  assign \arg0_2Dcon_||_2MyTrue_1MyTrue_d  = MyTrue_dc((& {\arg0_2Dcon_||_2MyTrue_d [0]}), \arg0_2Dcon_||_2MyTrue_d );
  assign {\arg0_2Dcon_||_2MyTrue_r } = {1 {(\arg0_2Dcon_||_2MyTrue_1MyTrue_r  && \arg0_2Dcon_||_2MyTrue_1MyTrue_d [0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_2Dcon_||_3,MyBool) [(arg0_2Dcon_||_1MyFalse,MyBool),
                                            (arg0_2Dcon_||_2MyTrue_1MyTrue,MyBool)] > (arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux ;
  logic [1:0] \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_onehot ;
  always_comb
    unique case (\arg0_2Dcon_||_3_d [1:1])
      1'd0:
        {\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_onehot ,
         \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux } = {2'd1,
                                                                             \arg0_2Dcon_||_1MyFalse_d };
      1'd1:
        {\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_onehot ,
         \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux } = {2'd2,
                                                                             \arg0_2Dcon_||_2MyTrue_1MyTrue_d };
      default:
        {\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_onehot ,
         \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux } = {2'd0,
                                                                             {1'd0, 1'd0}};
    endcase
  assign \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d  = {\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux [1:1],
                                                                          (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux [0] && \arg0_2Dcon_||_3_d [0])};
  assign \arg0_2Dcon_||_3_r  = (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d [0] && \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_r );
  assign {\arg0_2Dcon_||_2MyTrue_1MyTrue_r ,
          \arg0_2Dcon_||_1MyFalse_r } = (\arg0_2Dcon_||_3_r  ? \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_onehot  :
                                         2'd0);
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty Go) : (arg0_3,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go) > [(arg0_3Dcon_||,Go)] */
  assign \arg0_3Dcon_||_d  = (arg0_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]);
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r = (\arg0_3Dcon_||_r  && (arg0_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  assign arg0_3_r = (\arg0_3Dcon_||_r  && (arg0_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  
  /* mux (Ty MyDTBool_Bool_Bool,
     Ty MyBool) : (arg0_4,MyDTBool_Bool_Bool) [(arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux,MyBool)] > (arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux,MyBool) */
  assign \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_d  = {\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d [1:1],
                                                                              (arg0_4_d[0] && \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d [0])};
  assign \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_r  = (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_r  && (arg0_4_d[0] && \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d [0]));
  assign arg0_4_r = (\arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_mux_r  && (arg0_4_d[0] && \arg0_2Dcon_||_1MyFalse_1arg0_2Dcon_||_2MyTrue_1MyTrue_mux_d [0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool,
          Dcon TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool) : (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1,TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool) > [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4,Go),
                                                                                                                                                                                                                                                                                                                                (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                                (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0,Pointer_CT$wmAdd_Bool)] */
  logic [4:0] call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted;
  logic [4:0] call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_done;
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d = (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0] && (! call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted[0]));
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d = (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0] && (! call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted[1]));
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[16:1],
                                                                                                                                  (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0] && (! call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted[2]))};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[32:17],
                                                                                                                                  (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0] && (! call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted[3]))};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[48:33],
                                                                                                                               (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0] && (! call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted[4]))};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_done = (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted | ({call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d[0],
                                                                                                                                                                                                                                                           call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d[0],
                                                                                                                                                                                                                                                           call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d[0],
                                                                                                                                                                                                                                                           call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d[0],
                                                                                                                                                                                                                                                           call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d[0]} & {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_r,
                                                                                                                                                                                                                                                                                                                                                                                     call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_r,
                                                                                                                                                                                                                                                                                                                                                                                     call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_r}));
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_r = (& call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted <= 5'd0;
    else
      call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_emitted <= (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_r ? 5'd0 :
                                                                                                                                 call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_done);
  
  /* rbuf (Ty Go) : (call_$wmAdd_Bool_goConst,Go) > (call_$wmAdd_Bool_initBufi,Go) */
  Go_t call_$wmAdd_Bool_goConst_buf;
  assign call_$wmAdd_Bool_goConst_r = (! call_$wmAdd_Bool_goConst_buf[0]);
  assign call_$wmAdd_Bool_initBufi_d = (call_$wmAdd_Bool_goConst_buf[0] ? call_$wmAdd_Bool_goConst_buf :
                                        call_$wmAdd_Bool_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Bool_goConst_buf <= 1'd0;
    else
      if ((call_$wmAdd_Bool_initBufi_r && call_$wmAdd_Bool_goConst_buf[0]))
        call_$wmAdd_Bool_goConst_buf <= 1'd0;
      else if (((! call_$wmAdd_Bool_initBufi_r) && (! call_$wmAdd_Bool_goConst_buf[0])))
        call_$wmAdd_Bool_goConst_buf <= call_$wmAdd_Bool_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wmAdd_Bool_goMux1,Go),
                           (lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf,Go),
                           (lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf,Go),
                           (lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf,Go),
                           (lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf,Go)] > (go_4_goMux_choice,C5) (go_4_goMux_data,Go) */
  logic [4:0] call_$wmAdd_Bool_goMux1_select_d;
  assign call_$wmAdd_Bool_goMux1_select_d = ((| call_$wmAdd_Bool_goMux1_select_q) ? call_$wmAdd_Bool_goMux1_select_q :
                                             (call_$wmAdd_Bool_goMux1_d[0] ? 5'd1 :
                                              (lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_d[0] ? 5'd2 :
                                               (lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_d[0] ? 5'd4 :
                                                (lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_d[0] ? 5'd8 :
                                                 (lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                  5'd0))))));
  logic [4:0] call_$wmAdd_Bool_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Bool_goMux1_select_q <= 5'd0;
    else
      call_$wmAdd_Bool_goMux1_select_q <= (call_$wmAdd_Bool_goMux1_done ? 5'd0 :
                                           call_$wmAdd_Bool_goMux1_select_d);
  logic [1:0] call_$wmAdd_Bool_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Bool_goMux1_emit_q <= 2'd0;
    else
      call_$wmAdd_Bool_goMux1_emit_q <= (call_$wmAdd_Bool_goMux1_done ? 2'd0 :
                                         call_$wmAdd_Bool_goMux1_emit_d);
  logic [1:0] call_$wmAdd_Bool_goMux1_emit_d;
  assign call_$wmAdd_Bool_goMux1_emit_d = (call_$wmAdd_Bool_goMux1_emit_q | ({go_4_goMux_choice_d[0],
                                                                              go_4_goMux_data_d[0]} & {go_4_goMux_choice_r,
                                                                                                       go_4_goMux_data_r}));
  logic call_$wmAdd_Bool_goMux1_done;
  assign call_$wmAdd_Bool_goMux1_done = (& call_$wmAdd_Bool_goMux1_emit_d);
  assign {lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_r,
          lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_r,
          lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_r,
          lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_r,
          call_$wmAdd_Bool_goMux1_r} = (call_$wmAdd_Bool_goMux1_done ? call_$wmAdd_Bool_goMux1_select_d :
                                        5'd0);
  assign go_4_goMux_data_d = ((call_$wmAdd_Bool_goMux1_select_d[0] && (! call_$wmAdd_Bool_goMux1_emit_q[0])) ? call_$wmAdd_Bool_goMux1_d :
                              ((call_$wmAdd_Bool_goMux1_select_d[1] && (! call_$wmAdd_Bool_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_d :
                               ((call_$wmAdd_Bool_goMux1_select_d[2] && (! call_$wmAdd_Bool_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_d :
                                ((call_$wmAdd_Bool_goMux1_select_d[3] && (! call_$wmAdd_Bool_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_d :
                                 ((call_$wmAdd_Bool_goMux1_select_d[4] && (! call_$wmAdd_Bool_goMux1_emit_q[0])) ? lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_4_goMux_choice_d = ((call_$wmAdd_Bool_goMux1_select_d[0] && (! call_$wmAdd_Bool_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_$wmAdd_Bool_goMux1_select_d[1] && (! call_$wmAdd_Bool_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_$wmAdd_Bool_goMux1_select_d[2] && (! call_$wmAdd_Bool_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_$wmAdd_Bool_goMux1_select_d[3] && (! call_$wmAdd_Bool_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_$wmAdd_Bool_goMux1_select_d[4] && (! call_$wmAdd_Bool_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wmAdd_Bool_initBuf,Go) > [(call_$wmAdd_Bool_unlockFork1,Go),
                                                (call_$wmAdd_Bool_unlockFork2,Go),
                                                (call_$wmAdd_Bool_unlockFork3,Go),
                                                (call_$wmAdd_Bool_unlockFork4,Go),
                                                (call_$wmAdd_Bool_unlockFork5,Go)] */
  logic [4:0] call_$wmAdd_Bool_initBuf_emitted;
  logic [4:0] call_$wmAdd_Bool_initBuf_done;
  assign call_$wmAdd_Bool_unlockFork1_d = (call_$wmAdd_Bool_initBuf_d[0] && (! call_$wmAdd_Bool_initBuf_emitted[0]));
  assign call_$wmAdd_Bool_unlockFork2_d = (call_$wmAdd_Bool_initBuf_d[0] && (! call_$wmAdd_Bool_initBuf_emitted[1]));
  assign call_$wmAdd_Bool_unlockFork3_d = (call_$wmAdd_Bool_initBuf_d[0] && (! call_$wmAdd_Bool_initBuf_emitted[2]));
  assign call_$wmAdd_Bool_unlockFork4_d = (call_$wmAdd_Bool_initBuf_d[0] && (! call_$wmAdd_Bool_initBuf_emitted[3]));
  assign call_$wmAdd_Bool_unlockFork5_d = (call_$wmAdd_Bool_initBuf_d[0] && (! call_$wmAdd_Bool_initBuf_emitted[4]));
  assign call_$wmAdd_Bool_initBuf_done = (call_$wmAdd_Bool_initBuf_emitted | ({call_$wmAdd_Bool_unlockFork5_d[0],
                                                                               call_$wmAdd_Bool_unlockFork4_d[0],
                                                                               call_$wmAdd_Bool_unlockFork3_d[0],
                                                                               call_$wmAdd_Bool_unlockFork2_d[0],
                                                                               call_$wmAdd_Bool_unlockFork1_d[0]} & {call_$wmAdd_Bool_unlockFork5_r,
                                                                                                                     call_$wmAdd_Bool_unlockFork4_r,
                                                                                                                     call_$wmAdd_Bool_unlockFork3_r,
                                                                                                                     call_$wmAdd_Bool_unlockFork2_r,
                                                                                                                     call_$wmAdd_Bool_unlockFork1_r}));
  assign call_$wmAdd_Bool_initBuf_r = (& call_$wmAdd_Bool_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Bool_initBuf_emitted <= 5'd0;
    else
      call_$wmAdd_Bool_initBuf_emitted <= (call_$wmAdd_Bool_initBuf_r ? 5'd0 :
                                           call_$wmAdd_Bool_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wmAdd_Bool_initBufi,Go) > (call_$wmAdd_Bool_initBuf,Go) */
  assign call_$wmAdd_Bool_initBufi_r = ((! call_$wmAdd_Bool_initBuf_d[0]) || call_$wmAdd_Bool_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wmAdd_Bool_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wmAdd_Bool_initBufi_r)
        call_$wmAdd_Bool_initBuf_d <= call_$wmAdd_Bool_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wmAdd_Bool_unlockFork1,Go) [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4,Go)] > (call_$wmAdd_Bool_goMux1,Go) */
  assign call_$wmAdd_Bool_goMux1_d = (call_$wmAdd_Bool_unlockFork1_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d[0]);
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_r = (call_$wmAdd_Bool_goMux1_r && (call_$wmAdd_Bool_unlockFork1_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d[0]));
  assign call_$wmAdd_Bool_unlockFork1_r = (call_$wmAdd_Bool_goMux1_r && (call_$wmAdd_Bool_unlockFork1_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolgo_4_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool_Bool) : (call_$wmAdd_Bool_unlockFork2,Go) [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1,MyDTBool_Bool_Bool)] > (call_$wmAdd_Bool_goMux2,MyDTBool_Bool_Bool) */
  assign call_$wmAdd_Bool_goMux2_d = (call_$wmAdd_Bool_unlockFork2_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d[0]);
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_r = (call_$wmAdd_Bool_goMux2_r && (call_$wmAdd_Bool_unlockFork2_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d[0]));
  assign call_$wmAdd_Bool_unlockFork2_r = (call_$wmAdd_Bool_goMux2_r && (call_$wmAdd_Bool_unlockFork2_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolwsib_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_$wmAdd_Bool_unlockFork3,Go) [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1,Pointer_QTree_Bool)] > (call_$wmAdd_Bool_goMux3,Pointer_QTree_Bool) */
  assign call_$wmAdd_Bool_goMux3_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d[16:1],
                                      (call_$wmAdd_Bool_unlockFork3_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d[0])};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_r = (call_$wmAdd_Bool_goMux3_r && (call_$wmAdd_Bool_unlockFork3_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d[0]));
  assign call_$wmAdd_Bool_unlockFork3_r = (call_$wmAdd_Bool_goMux3_r && (call_$wmAdd_Bool_unlockFork3_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw1sic_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_$wmAdd_Bool_unlockFork4,Go) [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1,Pointer_QTree_Bool)] > (call_$wmAdd_Bool_goMux4,Pointer_QTree_Bool) */
  assign call_$wmAdd_Bool_goMux4_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d[16:1],
                                      (call_$wmAdd_Bool_unlockFork4_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d[0])};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_r = (call_$wmAdd_Bool_goMux4_r && (call_$wmAdd_Bool_unlockFork4_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d[0]));
  assign call_$wmAdd_Bool_unlockFork4_r = (call_$wmAdd_Bool_goMux4_r && (call_$wmAdd_Bool_unlockFork4_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolw2sid_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wmAdd_Bool) : (call_$wmAdd_Bool_unlockFork5,Go) [(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0,Pointer_CT$wmAdd_Bool)] > (call_$wmAdd_Bool_goMux5,Pointer_CT$wmAdd_Bool) */
  assign call_$wmAdd_Bool_goMux5_d = {call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d[16:1],
                                      (call_$wmAdd_Bool_unlockFork5_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d[0])};
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_r = (call_$wmAdd_Bool_goMux5_r && (call_$wmAdd_Bool_unlockFork5_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d[0]));
  assign call_$wmAdd_Bool_unlockFork5_r = (call_$wmAdd_Bool_goMux5_r && (call_$wmAdd_Bool_unlockFork5_d[0] && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Boolsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) : (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) > [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5,Go),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r,Pointer_MaskQTree),
                                                                                                                                                                                                                                                                          (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1,Pointer_CTmain_mask_Bool)] */
  logic [3:0] call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted;
  logic [3:0] call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done;
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d = (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[0]));
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[16:1],
                                                                                                               (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[1]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[32:17],
                                                                                                                 (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[2]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[48:33],
                                                                                                                 (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0] && (! call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted[3]))};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done = (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted | ({call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d[0],
                                                                                                                                                                                                                           call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]} & {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_r,
                                                                                                                                                                                                                                                                                                                                     call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r}));
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r = (& call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted <= 4'd0;
    else
      call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_emitted <= (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r ? 4'd0 :
                                                                                                                 call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_done);
  
  /* rbuf (Ty Go) : (call_main_mask_Bool_goConst,Go) > (call_main_mask_Bool_initBufi,Go) */
  Go_t call_main_mask_Bool_goConst_buf;
  assign call_main_mask_Bool_goConst_r = (! call_main_mask_Bool_goConst_buf[0]);
  assign call_main_mask_Bool_initBufi_d = (call_main_mask_Bool_goConst_buf[0] ? call_main_mask_Bool_goConst_buf :
                                           call_main_mask_Bool_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goConst_buf <= 1'd0;
    else
      if ((call_main_mask_Bool_initBufi_r && call_main_mask_Bool_goConst_buf[0]))
        call_main_mask_Bool_goConst_buf <= 1'd0;
      else if (((! call_main_mask_Bool_initBufi_r) && (! call_main_mask_Bool_goConst_buf[0])))
        call_main_mask_Bool_goConst_buf <= call_main_mask_Bool_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_mask_Bool_goMux1,Go),
                           (lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf,Go),
                           (lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf,Go),
                           (lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf,Go),
                           (lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf,Go)] > (go_5_goMux_choice,C5) (go_5_goMux_data,Go) */
  logic [4:0] call_main_mask_Bool_goMux1_select_d;
  assign call_main_mask_Bool_goMux1_select_d = ((| call_main_mask_Bool_goMux1_select_q) ? call_main_mask_Bool_goMux1_select_q :
                                                (call_main_mask_Bool_goMux1_d[0] ? 5'd1 :
                                                 (lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_d[0] ? 5'd2 :
                                                  (lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_d[0] ? 5'd4 :
                                                   (lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_d[0] ? 5'd8 :
                                                    (lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                     5'd0))))));
  logic [4:0] call_main_mask_Bool_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goMux1_select_q <= 5'd0;
    else
      call_main_mask_Bool_goMux1_select_q <= (call_main_mask_Bool_goMux1_done ? 5'd0 :
                                              call_main_mask_Bool_goMux1_select_d);
  logic [1:0] call_main_mask_Bool_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_goMux1_emit_q <= 2'd0;
    else
      call_main_mask_Bool_goMux1_emit_q <= (call_main_mask_Bool_goMux1_done ? 2'd0 :
                                            call_main_mask_Bool_goMux1_emit_d);
  logic [1:0] call_main_mask_Bool_goMux1_emit_d;
  assign call_main_mask_Bool_goMux1_emit_d = (call_main_mask_Bool_goMux1_emit_q | ({go_5_goMux_choice_d[0],
                                                                                    go_5_goMux_data_d[0]} & {go_5_goMux_choice_r,
                                                                                                             go_5_goMux_data_r}));
  logic call_main_mask_Bool_goMux1_done;
  assign call_main_mask_Bool_goMux1_done = (& call_main_mask_Bool_goMux1_emit_d);
  assign {lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_r,
          lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_r,
          lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_r,
          lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_r,
          call_main_mask_Bool_goMux1_r} = (call_main_mask_Bool_goMux1_done ? call_main_mask_Bool_goMux1_select_d :
                                           5'd0);
  assign go_5_goMux_data_d = ((call_main_mask_Bool_goMux1_select_d[0] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? call_main_mask_Bool_goMux1_d :
                              ((call_main_mask_Bool_goMux1_select_d[1] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_d :
                               ((call_main_mask_Bool_goMux1_select_d[2] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_d :
                                ((call_main_mask_Bool_goMux1_select_d[3] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_d :
                                 ((call_main_mask_Bool_goMux1_select_d[4] && (! call_main_mask_Bool_goMux1_emit_q[0])) ? lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_5_goMux_choice_d = ((call_main_mask_Bool_goMux1_select_d[0] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_main_mask_Bool_goMux1_select_d[1] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_main_mask_Bool_goMux1_select_d[2] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_main_mask_Bool_goMux1_select_d[3] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_main_mask_Bool_goMux1_select_d[4] && (! call_main_mask_Bool_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_mask_Bool_initBuf,Go) > [(call_main_mask_Bool_unlockFork1,Go),
                                                   (call_main_mask_Bool_unlockFork2,Go),
                                                   (call_main_mask_Bool_unlockFork3,Go),
                                                   (call_main_mask_Bool_unlockFork4,Go)] */
  logic [3:0] call_main_mask_Bool_initBuf_emitted;
  logic [3:0] call_main_mask_Bool_initBuf_done;
  assign call_main_mask_Bool_unlockFork1_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[0]));
  assign call_main_mask_Bool_unlockFork2_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[1]));
  assign call_main_mask_Bool_unlockFork3_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[2]));
  assign call_main_mask_Bool_unlockFork4_d = (call_main_mask_Bool_initBuf_d[0] && (! call_main_mask_Bool_initBuf_emitted[3]));
  assign call_main_mask_Bool_initBuf_done = (call_main_mask_Bool_initBuf_emitted | ({call_main_mask_Bool_unlockFork4_d[0],
                                                                                     call_main_mask_Bool_unlockFork3_d[0],
                                                                                     call_main_mask_Bool_unlockFork2_d[0],
                                                                                     call_main_mask_Bool_unlockFork1_d[0]} & {call_main_mask_Bool_unlockFork4_r,
                                                                                                                              call_main_mask_Bool_unlockFork3_r,
                                                                                                                              call_main_mask_Bool_unlockFork2_r,
                                                                                                                              call_main_mask_Bool_unlockFork1_r}));
  assign call_main_mask_Bool_initBuf_r = (& call_main_mask_Bool_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_initBuf_emitted <= 4'd0;
    else
      call_main_mask_Bool_initBuf_emitted <= (call_main_mask_Bool_initBuf_r ? 4'd0 :
                                              call_main_mask_Bool_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_mask_Bool_initBufi,Go) > (call_main_mask_Bool_initBuf,Go) */
  assign call_main_mask_Bool_initBufi_r = ((! call_main_mask_Bool_initBuf_d[0]) || call_main_mask_Bool_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_main_mask_Bool_initBuf_d <= Go_dc(1'd1);
    else
      if (call_main_mask_Bool_initBufi_r)
        call_main_mask_Bool_initBuf_d <= call_main_mask_Bool_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_mask_Bool_unlockFork1,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5,Go)] > (call_main_mask_Bool_goMux1,Go) */
  assign call_main_mask_Bool_goMux1_d = (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]);
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_r = (call_main_mask_Bool_goMux1_r && (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]));
  assign call_main_mask_Bool_unlockFork1_r = (call_main_mask_Bool_goMux1_r && (call_main_mask_Bool_unlockFork1_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolgo_5_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_main_mask_Bool_unlockFork2,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q,Pointer_QTree_Bool)] > (call_main_mask_Bool_goMux2,Pointer_QTree_Bool) */
  assign call_main_mask_Bool_goMux2_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d[16:1],
                                         (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_r = (call_main_mask_Bool_goMux2_r && (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d[0]));
  assign call_main_mask_Bool_unlockFork2_r = (call_main_mask_Bool_goMux2_r && (call_main_mask_Bool_unlockFork2_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolma8q_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_MaskQTree) : (call_main_mask_Bool_unlockFork3,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r,Pointer_MaskQTree)] > (call_main_mask_Bool_goMux3,Pointer_MaskQTree) */
  assign call_main_mask_Bool_goMux3_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d[16:1],
                                         (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_r = (call_main_mask_Bool_goMux3_r && (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d[0]));
  assign call_main_mask_Bool_unlockFork3_r = (call_main_mask_Bool_goMux3_r && (call_main_mask_Bool_unlockFork3_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolmska8r_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_mask_Bool) : (call_main_mask_Bool_unlockFork4,Go) [(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1,Pointer_CTmain_mask_Bool)] > (call_main_mask_Bool_goMux4,Pointer_CTmain_mask_Bool) */
  assign call_main_mask_Bool_goMux4_d = {call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[16:1],
                                         (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0])};
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_r = (call_main_mask_Bool_goMux4_r && (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0]));
  assign call_main_mask_Bool_unlockFork4_r = (call_main_mask_Bool_goMux4_r && (call_main_mask_Bool_unlockFork4_d[0] && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Boolsc_0_1_d[0]));
  
  /* buf (Ty QTree_Bool) : (es_0_1_1QVal_Bool,QTree_Bool) > (lizzieLet3_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_1_1QVal_Bool_bufchan_d;
  logic es_0_1_1QVal_Bool_bufchan_r;
  assign es_0_1_1QVal_Bool_r = ((! es_0_1_1QVal_Bool_bufchan_d[0]) || es_0_1_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_1QVal_Bool_r)
        es_0_1_1QVal_Bool_bufchan_d <= es_0_1_1QVal_Bool_d;
  QTree_Bool_t es_0_1_1QVal_Bool_bufchan_buf;
  assign es_0_1_1QVal_Bool_bufchan_r = (! es_0_1_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet3_1_argbuf_d = (es_0_1_1QVal_Bool_bufchan_buf[0] ? es_0_1_1QVal_Bool_bufchan_buf :
                                  es_0_1_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet3_1_argbuf_r && es_0_1_1QVal_Bool_bufchan_buf[0]))
        es_0_1_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet3_1_argbuf_r) && (! es_0_1_1QVal_Bool_bufchan_buf[0])))
        es_0_1_1QVal_Bool_bufchan_buf <= es_0_1_1QVal_Bool_bufchan_d;
  
  /* dcon (Ty MyDTBool_Bool_Bool,
      Dcon Dcon_||) : [(go_1,Go)] > (go_1Dcon_||,MyDTBool_Bool_Bool) */
  assign \go_1Dcon_||_d  = \Dcon_||_dc ((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(\go_1Dcon_||_r  && \go_1Dcon_||_d [0])}};
  
  /* buf (Ty MyDTBool_Bool_Bool) : (go_1Dcon_||,MyDTBool_Bool_Bool) > (es_2_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \go_1Dcon_||_bufchan_d ;
  logic \go_1Dcon_||_bufchan_r ;
  assign \go_1Dcon_||_r  = ((! \go_1Dcon_||_bufchan_d [0]) || \go_1Dcon_||_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_||_bufchan_d  <= 1'd0;
    else
      if (\go_1Dcon_||_r ) \go_1Dcon_||_bufchan_d  <= \go_1Dcon_||_d ;
  MyDTBool_Bool_Bool_t \go_1Dcon_||_bufchan_buf ;
  assign \go_1Dcon_||_bufchan_r  = (! \go_1Dcon_||_bufchan_buf [0]);
  assign es_2_1_argbuf_d = (\go_1Dcon_||_bufchan_buf [0] ? \go_1Dcon_||_bufchan_buf  :
                            \go_1Dcon_||_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_1Dcon_||_bufchan_buf  <= 1'd0;
    else
      if ((es_2_1_argbuf_r && \go_1Dcon_||_bufchan_buf [0]))
        \go_1Dcon_||_bufchan_buf  <= 1'd0;
      else if (((! es_2_1_argbuf_r) && (! \go_1Dcon_||_bufchan_buf [0])))
        \go_1Dcon_||_bufchan_buf  <= \go_1Dcon_||_bufchan_d ;
  
  /* buf (Ty Go) : (go_2,Go) > (go_2_argbuf,Go) */
  Go_t go_2_bufchan_d;
  logic go_2_bufchan_r;
  assign go_2_r = ((! go_2_bufchan_d[0]) || go_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_d <= 1'd0;
    else if (go_2_r) go_2_bufchan_d <= go_2_d;
  Go_t go_2_bufchan_buf;
  assign go_2_bufchan_r = (! go_2_bufchan_buf[0]);
  assign go_2_argbuf_d = (go_2_bufchan_buf[0] ? go_2_bufchan_buf :
                          go_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_bufchan_buf <= 1'd0;
    else
      if ((go_2_argbuf_r && go_2_bufchan_buf[0]))
        go_2_bufchan_buf <= 1'd0;
      else if (((! go_2_argbuf_r) && (! go_2_bufchan_buf[0])))
        go_2_bufchan_buf <= go_2_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Bool,
      Dcon L$wmAdd_Boolsbos) : [(go_2_1,Go)] > (go_2_1L$wmAdd_Boolsbos,CT$wmAdd_Bool) */
  assign go_2_1L$wmAdd_Boolsbos_d = L$wmAdd_Boolsbos_dc((& {go_2_1_d[0]}), go_2_1_d);
  assign {go_2_1_r} = {1 {(go_2_1L$wmAdd_Boolsbos_r && go_2_1L$wmAdd_Boolsbos_d[0])}};
  
  /* buf (Ty CT$wmAdd_Bool) : (go_2_1L$wmAdd_Boolsbos,CT$wmAdd_Bool) > (lizzieLet0_1_argbuf,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t go_2_1L$wmAdd_Boolsbos_bufchan_d;
  logic go_2_1L$wmAdd_Boolsbos_bufchan_r;
  assign go_2_1L$wmAdd_Boolsbos_r = ((! go_2_1L$wmAdd_Boolsbos_bufchan_d[0]) || go_2_1L$wmAdd_Boolsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_2_1L$wmAdd_Boolsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_2_1L$wmAdd_Boolsbos_r)
        go_2_1L$wmAdd_Boolsbos_bufchan_d <= go_2_1L$wmAdd_Boolsbos_d;
  CT$wmAdd_Bool_t go_2_1L$wmAdd_Boolsbos_bufchan_buf;
  assign go_2_1L$wmAdd_Boolsbos_bufchan_r = (! go_2_1L$wmAdd_Boolsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_2_1L$wmAdd_Boolsbos_bufchan_buf[0] ? go_2_1L$wmAdd_Boolsbos_bufchan_buf :
                                  go_2_1L$wmAdd_Boolsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_2_1L$wmAdd_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_2_1L$wmAdd_Boolsbos_bufchan_buf[0]))
        go_2_1L$wmAdd_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_2_1L$wmAdd_Boolsbos_bufchan_buf[0])))
        go_2_1L$wmAdd_Boolsbos_bufchan_buf <= go_2_1L$wmAdd_Boolsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_2_2,Go) > (go_2_2_argbuf,Go) */
  Go_t go_2_2_bufchan_d;
  logic go_2_2_bufchan_r;
  assign go_2_2_r = ((! go_2_2_bufchan_d[0]) || go_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_2_bufchan_d <= 1'd0;
    else if (go_2_2_r) go_2_2_bufchan_d <= go_2_2_d;
  Go_t go_2_2_bufchan_buf;
  assign go_2_2_bufchan_r = (! go_2_2_bufchan_buf[0]);
  assign go_2_2_argbuf_d = (go_2_2_bufchan_buf[0] ? go_2_2_bufchan_buf :
                            go_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2_2_bufchan_buf <= 1'd0;
    else
      if ((go_2_2_argbuf_r && go_2_2_bufchan_buf[0]))
        go_2_2_bufchan_buf <= 1'd0;
      else if (((! go_2_2_argbuf_r) && (! go_2_2_bufchan_buf[0])))
        go_2_2_bufchan_buf <= go_2_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool,
      Dcon TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool) : [(go_2_2_argbuf,Go),
                                                                                                            (wsib_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                            (w1sic_1_argbuf,Pointer_QTree_Bool),
                                                                                                            (w2sid_1_argbuf,Pointer_QTree_Bool),
                                                                                                            (lizzieLet11_1_argbuf,Pointer_CT$wmAdd_Bool)] > (call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1,TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool) */
  assign call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d = TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_dc((& {go_2_2_argbuf_d[0],
                                                                                                                                                                                                                                wsib_1_argbuf_d[0],
                                                                                                                                                                                                                                w1sic_1_argbuf_d[0],
                                                                                                                                                                                                                                w2sid_1_argbuf_d[0],
                                                                                                                                                                                                                                lizzieLet11_1_argbuf_d[0]}), go_2_2_argbuf_d, wsib_1_argbuf_d, w1sic_1_argbuf_d, w2sid_1_argbuf_d, lizzieLet11_1_argbuf_d);
  assign {go_2_2_argbuf_r,
          wsib_1_argbuf_r,
          w1sic_1_argbuf_r,
          w2sid_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = {5 {(call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_r && call_$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CT$wmAdd_Bool_1_d[0])}};
  
  /* dcon (Ty TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(go_2_argbuf,Go),
                                                                                    (es_2_1_argbuf,MyDTBool_Bool_Bool),
                                                                                    (m2a93_1,Pointer_QTree_Bool),
                                                                                    (m3a94_2,Pointer_QTree_Bool)] > ($wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d  = TupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {go_2_argbuf_d[0],
                                                                                                                                                                             es_2_1_argbuf_d[0],
                                                                                                                                                                             m2a93_1_d[0],
                                                                                                                                                                             m3a94_2_d[0]}), go_2_argbuf_d, es_2_1_argbuf_d, m2a93_1_d, m3a94_2_d);
  assign {go_2_argbuf_r,
          es_2_1_argbuf_r,
          m2a93_1_r,
          m3a94_2_r} = {4 {(\$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r  && \$wmAdd_BoolTupGo___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (go_3,Go) > (go_3_argbuf,Go) */
  Go_t go_3_bufchan_d;
  logic go_3_bufchan_r;
  assign go_3_r = ((! go_3_bufchan_d[0]) || go_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_d <= 1'd0;
    else if (go_3_r) go_3_bufchan_d <= go_3_d;
  Go_t go_3_bufchan_buf;
  assign go_3_bufchan_r = (! go_3_bufchan_buf[0]);
  assign go_3_argbuf_d = (go_3_bufchan_buf[0] ? go_3_bufchan_buf :
                          go_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_3_bufchan_buf <= 1'd0;
    else
      if ((go_3_argbuf_r && go_3_bufchan_buf[0]))
        go_3_bufchan_buf <= 1'd0;
      else if (((! go_3_argbuf_r) && (! go_3_bufchan_buf[0])))
        go_3_bufchan_buf <= go_3_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) : [(go_3_argbuf,Go),
                                                              (es_0_1_argbuf,Pointer_QTree_Bool),
                                                              (m1a92_0,Pointer_MaskQTree)] > (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) */
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d = TupGo___Pointer_QTree_Bool___Pointer_MaskQTree_dc((& {go_3_argbuf_d[0],
                                                                                                                                  es_0_1_argbuf_d[0],
                                                                                                                                  m1a92_0_d[0]}), go_3_argbuf_d, es_0_1_argbuf_d, m1a92_0_d);
  assign {go_3_argbuf_r,
          es_0_1_argbuf_r,
          m1a92_0_r} = {3 {(main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0])}};
  
  /* fork (Ty C5) : (go_4_goMux_choice,C5) > [(go_4_goMux_choice_1,C5),
                                         (go_4_goMux_choice_2,C5),
                                         (go_4_goMux_choice_3,C5),
                                         (go_4_goMux_choice_4,C5)] */
  logic [3:0] go_4_goMux_choice_emitted;
  logic [3:0] go_4_goMux_choice_done;
  assign go_4_goMux_choice_1_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[0]))};
  assign go_4_goMux_choice_2_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[1]))};
  assign go_4_goMux_choice_3_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[2]))};
  assign go_4_goMux_choice_4_d = {go_4_goMux_choice_d[3:1],
                                  (go_4_goMux_choice_d[0] && (! go_4_goMux_choice_emitted[3]))};
  assign go_4_goMux_choice_done = (go_4_goMux_choice_emitted | ({go_4_goMux_choice_4_d[0],
                                                                 go_4_goMux_choice_3_d[0],
                                                                 go_4_goMux_choice_2_d[0],
                                                                 go_4_goMux_choice_1_d[0]} & {go_4_goMux_choice_4_r,
                                                                                              go_4_goMux_choice_3_r,
                                                                                              go_4_goMux_choice_2_r,
                                                                                              go_4_goMux_choice_1_r}));
  assign go_4_goMux_choice_r = (& go_4_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4_goMux_choice_emitted <= 4'd0;
    else
      go_4_goMux_choice_emitted <= (go_4_goMux_choice_r ? 4'd0 :
                                    go_4_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool_Bool) : (go_4_goMux_choice_1,C5) [(call_$wmAdd_Bool_goMux2,MyDTBool_Bool_Bool),
                                                        (wsib_2_2_argbuf,MyDTBool_Bool_Bool),
                                                        (wsib_3_2_argbuf,MyDTBool_Bool_Bool),
                                                        (wsib_4_1_argbuf,MyDTBool_Bool_Bool),
                                                        (lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf,MyDTBool_Bool_Bool)] > (wsib_1_goMux_mux,MyDTBool_Bool_Bool) */
  logic [0:0] wsib_1_goMux_mux_mux;
  logic [4:0] wsib_1_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_1_d[3:1])
      3'd0:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd1,
                                                           call_$wmAdd_Bool_goMux2_d};
      3'd1:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd2,
                                                           wsib_2_2_argbuf_d};
      3'd2:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd4,
                                                           wsib_3_2_argbuf_d};
      3'd3:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd8,
                                                           wsib_4_1_argbuf_d};
      3'd4:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd16,
                                                           lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_d};
      default:
        {wsib_1_goMux_mux_onehot, wsib_1_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign wsib_1_goMux_mux_d = (wsib_1_goMux_mux_mux[0] && go_4_goMux_choice_1_d[0]);
  assign go_4_goMux_choice_1_r = (wsib_1_goMux_mux_d[0] && wsib_1_goMux_mux_r);
  assign {lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_r,
          wsib_4_1_argbuf_r,
          wsib_3_2_argbuf_r,
          wsib_2_2_argbuf_r,
          call_$wmAdd_Bool_goMux2_r} = (go_4_goMux_choice_1_r ? wsib_1_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_4_goMux_choice_2,C5) [(call_$wmAdd_Bool_goMux3,Pointer_QTree_Bool),
                                                        (q3a8j_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2a8i_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1a8h_3_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf,Pointer_QTree_Bool)] > (w1sic_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] w1sic_1_goMux_mux_mux;
  logic [4:0] w1sic_1_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_2_d[3:1])
      3'd0:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Bool_goMux3_d};
      3'd1:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd2,
                                                             q3a8j_1_1_argbuf_d};
      3'd2:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd4,
                                                             q2a8i_2_1_argbuf_d};
      3'd3:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd8,
                                                             q1a8h_3_1_argbuf_d};
      3'd4:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd16,
                                                             lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_d};
      default:
        {w1sic_1_goMux_mux_onehot, w1sic_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w1sic_1_goMux_mux_d = {w1sic_1_goMux_mux_mux[16:1],
                                (w1sic_1_goMux_mux_mux[0] && go_4_goMux_choice_2_d[0])};
  assign go_4_goMux_choice_2_r = (w1sic_1_goMux_mux_d[0] && w1sic_1_goMux_mux_r);
  assign {lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_r,
          q1a8h_3_1_argbuf_r,
          q2a8i_2_1_argbuf_r,
          q3a8j_1_1_argbuf_r,
          call_$wmAdd_Bool_goMux3_r} = (go_4_goMux_choice_2_r ? w1sic_1_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_4_goMux_choice_3,C5) [(call_$wmAdd_Bool_goMux4,Pointer_QTree_Bool),
                                                        (t3a8o_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8n_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8m_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4a8p_1_argbuf,Pointer_QTree_Bool)] > (w2sid_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] w2sid_1_goMux_mux_mux;
  logic [4:0] w2sid_1_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_3_d[3:1])
      3'd0:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd1,
                                                             call_$wmAdd_Bool_goMux4_d};
      3'd1:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd2,
                                                             t3a8o_1_1_argbuf_d};
      3'd2:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd4,
                                                             t2a8n_2_1_argbuf_d};
      3'd3:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd8,
                                                             t1a8m_3_1_argbuf_d};
      3'd4:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd16,
                                                             t4a8p_1_argbuf_d};
      default:
        {w2sid_1_goMux_mux_onehot, w2sid_1_goMux_mux_mux} = {5'd0,
                                                             {16'd0, 1'd0}};
    endcase
  assign w2sid_1_goMux_mux_d = {w2sid_1_goMux_mux_mux[16:1],
                                (w2sid_1_goMux_mux_mux[0] && go_4_goMux_choice_3_d[0])};
  assign go_4_goMux_choice_3_r = (w2sid_1_goMux_mux_d[0] && w2sid_1_goMux_mux_r);
  assign {t4a8p_1_argbuf_r,
          t1a8m_3_1_argbuf_r,
          t2a8n_2_1_argbuf_r,
          t3a8o_1_1_argbuf_r,
          call_$wmAdd_Bool_goMux4_r} = (go_4_goMux_choice_3_r ? w2sid_1_goMux_mux_onehot :
                                        5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wmAdd_Bool) : (go_4_goMux_choice_4,C5) [(call_$wmAdd_Bool_goMux5,Pointer_CT$wmAdd_Bool),
                                                           (sca2_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                           (sca1_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                           (sca0_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                           (sca3_1_argbuf,Pointer_CT$wmAdd_Bool)] > (sc_0_goMux_mux,Pointer_CT$wmAdd_Bool) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_4_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wmAdd_Bool_goMux5_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_4_goMux_choice_4_d[0])};
  assign go_4_goMux_choice_4_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wmAdd_Bool_goMux5_r} = (go_4_goMux_choice_4_r ? sc_0_goMux_mux_onehot :
                                        5'd0);
  
  /* fork (Ty C5) : (go_5_goMux_choice,C5) > [(go_5_goMux_choice_1,C5),
                                         (go_5_goMux_choice_2,C5),
                                         (go_5_goMux_choice_3,C5)] */
  logic [2:0] go_5_goMux_choice_emitted;
  logic [2:0] go_5_goMux_choice_done;
  assign go_5_goMux_choice_1_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[0]))};
  assign go_5_goMux_choice_2_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[1]))};
  assign go_5_goMux_choice_3_d = {go_5_goMux_choice_d[3:1],
                                  (go_5_goMux_choice_d[0] && (! go_5_goMux_choice_emitted[2]))};
  assign go_5_goMux_choice_done = (go_5_goMux_choice_emitted | ({go_5_goMux_choice_3_d[0],
                                                                 go_5_goMux_choice_2_d[0],
                                                                 go_5_goMux_choice_1_d[0]} & {go_5_goMux_choice_3_r,
                                                                                              go_5_goMux_choice_2_r,
                                                                                              go_5_goMux_choice_1_r}));
  assign go_5_goMux_choice_r = (& go_5_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_goMux_choice_emitted <= 3'd0;
    else
      go_5_goMux_choice_emitted <= (go_5_goMux_choice_r ? 3'd0 :
                                    go_5_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_5_goMux_choice_1,C5) [(call_main_mask_Bool_goMux2,Pointer_QTree_Bool),
                                                        (t3a8z_1_1_argbuf,Pointer_QTree_Bool),
                                                        (t2a8y_2_1_argbuf,Pointer_QTree_Bool),
                                                        (t1a8x_3_1_argbuf,Pointer_QTree_Bool),
                                                        (t4a8A_1_argbuf,Pointer_QTree_Bool)] > (ma8q_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] ma8q_goMux_mux_mux;
  logic [4:0] ma8q_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_1_d[3:1])
      3'd0:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd1,
                                                       call_main_mask_Bool_goMux2_d};
      3'd1:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd2,
                                                       t3a8z_1_1_argbuf_d};
      3'd2:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd4,
                                                       t2a8y_2_1_argbuf_d};
      3'd3:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd8,
                                                       t1a8x_3_1_argbuf_d};
      3'd4:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd16,
                                                       t4a8A_1_argbuf_d};
      default:
        {ma8q_goMux_mux_onehot, ma8q_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign ma8q_goMux_mux_d = {ma8q_goMux_mux_mux[16:1],
                             (ma8q_goMux_mux_mux[0] && go_5_goMux_choice_1_d[0])};
  assign go_5_goMux_choice_1_r = (ma8q_goMux_mux_d[0] && ma8q_goMux_mux_r);
  assign {t4a8A_1_argbuf_r,
          t1a8x_3_1_argbuf_r,
          t2a8y_2_1_argbuf_r,
          t3a8z_1_1_argbuf_r,
          call_main_mask_Bool_goMux2_r} = (go_5_goMux_choice_1_r ? ma8q_goMux_mux_onehot :
                                           5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_MaskQTree) : (go_5_goMux_choice_2,C5) [(call_main_mask_Bool_goMux3,Pointer_MaskQTree),
                                                       (q3a8u_1_1_argbuf,Pointer_MaskQTree),
                                                       (q2a8t_2_1_argbuf,Pointer_MaskQTree),
                                                       (q1a8s_3_1_argbuf,Pointer_MaskQTree),
                                                       (lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree)] > (mska8r_goMux_mux,Pointer_MaskQTree) */
  logic [16:0] mska8r_goMux_mux_mux;
  logic [4:0] mska8r_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_2_d[3:1])
      3'd0:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Bool_goMux3_d};
      3'd1:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd2,
                                                           q3a8u_1_1_argbuf_d};
      3'd2:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd4,
                                                           q2a8t_2_1_argbuf_d};
      3'd3:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd8,
                                                           q1a8s_3_1_argbuf_d};
      3'd4:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd16,
                                                           lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_d};
      default:
        {mska8r_goMux_mux_onehot, mska8r_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign mska8r_goMux_mux_d = {mska8r_goMux_mux_mux[16:1],
                               (mska8r_goMux_mux_mux[0] && go_5_goMux_choice_2_d[0])};
  assign go_5_goMux_choice_2_r = (mska8r_goMux_mux_d[0] && mska8r_goMux_mux_r);
  assign {lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_r,
          q1a8s_3_1_argbuf_r,
          q2a8t_2_1_argbuf_r,
          q3a8u_1_1_argbuf_r,
          call_main_mask_Bool_goMux3_r} = (go_5_goMux_choice_2_r ? mska8r_goMux_mux_onehot :
                                           5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_mask_Bool) : (go_5_goMux_choice_3,C5) [(call_main_mask_Bool_goMux4,Pointer_CTmain_mask_Bool),
                                                              (sca2_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca1_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca0_1_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sca3_1_1_argbuf,Pointer_CTmain_mask_Bool)] > (sc_0_1_goMux_mux,Pointer_CTmain_mask_Bool) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_5_goMux_choice_3_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           call_main_mask_Bool_goMux4_d};
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_5_goMux_choice_3_d[0])};
  assign go_5_goMux_choice_3_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          call_main_mask_Bool_goMux4_r} = (go_5_goMux_choice_3_r ? sc_0_1_goMux_mux_onehot :
                                           5'd0);
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lmain_mask_Boolsbos) : [(go_6_1,Go)] > (go_6_1Lmain_mask_Boolsbos,CTmain_mask_Bool) */
  assign go_6_1Lmain_mask_Boolsbos_d = Lmain_mask_Boolsbos_dc((& {go_6_1_d[0]}), go_6_1_d);
  assign {go_6_1_r} = {1 {(go_6_1Lmain_mask_Boolsbos_r && go_6_1Lmain_mask_Boolsbos_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (go_6_1Lmain_mask_Boolsbos,CTmain_mask_Bool) > (lizzieLet18_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t go_6_1Lmain_mask_Boolsbos_bufchan_d;
  logic go_6_1Lmain_mask_Boolsbos_bufchan_r;
  assign go_6_1Lmain_mask_Boolsbos_r = ((! go_6_1Lmain_mask_Boolsbos_bufchan_d[0]) || go_6_1Lmain_mask_Boolsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1Lmain_mask_Boolsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_6_1Lmain_mask_Boolsbos_r)
        go_6_1Lmain_mask_Boolsbos_bufchan_d <= go_6_1Lmain_mask_Boolsbos_d;
  CTmain_mask_Bool_t go_6_1Lmain_mask_Boolsbos_bufchan_buf;
  assign go_6_1Lmain_mask_Boolsbos_bufchan_r = (! go_6_1Lmain_mask_Boolsbos_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (go_6_1Lmain_mask_Boolsbos_bufchan_buf[0] ? go_6_1Lmain_mask_Boolsbos_bufchan_buf :
                                   go_6_1Lmain_mask_Boolsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_6_1Lmain_mask_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && go_6_1Lmain_mask_Boolsbos_bufchan_buf[0]))
        go_6_1Lmain_mask_Boolsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! go_6_1Lmain_mask_Boolsbos_bufchan_buf[0])))
        go_6_1Lmain_mask_Boolsbos_bufchan_buf <= go_6_1Lmain_mask_Boolsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_6_2,Go) > (go_6_2_argbuf,Go) */
  Go_t go_6_2_bufchan_d;
  logic go_6_2_bufchan_r;
  assign go_6_2_r = ((! go_6_2_bufchan_d[0]) || go_6_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_d <= 1'd0;
    else if (go_6_2_r) go_6_2_bufchan_d <= go_6_2_d;
  Go_t go_6_2_bufchan_buf;
  assign go_6_2_bufchan_r = (! go_6_2_bufchan_buf[0]);
  assign go_6_2_argbuf_d = (go_6_2_bufchan_buf[0] ? go_6_2_bufchan_buf :
                            go_6_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_2_bufchan_buf <= 1'd0;
    else
      if ((go_6_2_argbuf_r && go_6_2_bufchan_buf[0]))
        go_6_2_bufchan_buf <= 1'd0;
      else if (((! go_6_2_argbuf_r) && (! go_6_2_bufchan_buf[0])))
        go_6_2_bufchan_buf <= go_6_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool,
      Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) : [(go_6_2_argbuf,Go),
                                                                                         (ma8q_1_1_argbuf,Pointer_QTree_Bool),
                                                                                         (mska8r_1_1_argbuf,Pointer_MaskQTree),
                                                                                         (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Bool)] > (call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool) */
  assign call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d = TupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_dc((& {go_6_2_argbuf_d[0],
                                                                                                                                                                                             ma8q_1_1_argbuf_d[0],
                                                                                                                                                                                             mska8r_1_1_argbuf_d[0],
                                                                                                                                                                                             lizzieLet4_1_1_argbuf_d[0]}), go_6_2_argbuf_d, ma8q_1_1_argbuf_d, mska8r_1_1_argbuf_d, lizzieLet4_1_1_argbuf_d);
  assign {go_6_2_argbuf_r,
          ma8q_1_1_argbuf_r,
          mska8r_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r} = {4 {(call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_r && call_main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree___Pointer_CTmain_mask_Bool_1_d[0])}};
  
  /* fork (Ty C10) : (go_7_goMux_choice,C10) > [(go_7_goMux_choice_1,C10),
                                           (go_7_goMux_choice_2,C10)] */
  logic [1:0] go_7_goMux_choice_emitted;
  logic [1:0] go_7_goMux_choice_done;
  assign go_7_goMux_choice_1_d = {go_7_goMux_choice_d[4:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[0]))};
  assign go_7_goMux_choice_2_d = {go_7_goMux_choice_d[4:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[1]))};
  assign go_7_goMux_choice_done = (go_7_goMux_choice_emitted | ({go_7_goMux_choice_2_d[0],
                                                                 go_7_goMux_choice_1_d[0]} & {go_7_goMux_choice_2_r,
                                                                                              go_7_goMux_choice_1_r}));
  assign go_7_goMux_choice_r = (& go_7_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_goMux_choice_emitted <= 2'd0;
    else
      go_7_goMux_choice_emitted <= (go_7_goMux_choice_r ? 2'd0 :
                                    go_7_goMux_choice_done);
  
  /* mux (Ty C10,
     Ty Pointer_QTree_Bool) : (go_7_goMux_choice_1,C10) [(lizzieLet1_7QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet5_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet6_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet7_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet8_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet9_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet10_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [9:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_1_d[4:1])
      4'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet1_7QNone_Bool_1_argbuf_d};
      4'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd2,
                                                               contRet_0_1_argbuf_d};
      4'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_d};
      4'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet5_1_argbuf_d};
      4'd4:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet6_1_argbuf_d};
      4'd5:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet7_1_argbuf_d};
      4'd6:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_d};
      4'd7:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet8_1_argbuf_d};
      4'd8:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet9_1_argbuf_d};
      4'd9:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet10_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_7_goMux_choice_1_d[0])};
  assign go_7_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet10_1_argbuf_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet6_1_argbuf_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet1_7QNone_Bool_1_argbuf_r} = (go_7_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                                10'd0);
  
  /* mux (Ty C10,
     Ty Pointer_CT$wmAdd_Bool) : (go_7_goMux_choice_2,C10) [(lizzieLet1_5QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (sc_0_5_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool),
                                                            (lizzieLet1_5QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool)] > (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Bool) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [9:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_2_d[4:1])
      4'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd1,
                                                               lizzieLet1_5QNone_Bool_1_argbuf_d};
      4'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd2,
                                                               sc_0_5_1_argbuf_d};
      4'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd4,
                                                               lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_d};
      4'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd8,
                                                               lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_d};
      4'd4:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd16,
                                                               lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_d};
      4'd5:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd32,
                                                               lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_d};
      4'd6:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd64,
                                                               lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_d};
      4'd7:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd128,
                                                               lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_d};
      4'd8:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd256,
                                                               lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_d};
      4'd9:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd512,
                                                               lizzieLet1_5QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {10'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_7_goMux_choice_2_d[0])};
  assign go_7_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet1_5QError_Bool_1_argbuf_r,
          lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_r,
          lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_r,
          lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_r,
          sc_0_5_1_argbuf_r,
          lizzieLet1_5QNone_Bool_1_argbuf_r} = (go_7_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                                10'd0);
  
  /* fork (Ty C6) : (go_8_goMux_choice,C6) > [(go_8_goMux_choice_1,C6),
                                         (go_8_goMux_choice_2,C6)] */
  logic [1:0] go_8_goMux_choice_emitted;
  logic [1:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 2'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 2'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Bool) : (go_8_goMux_choice_1,C6) [(lizzieLet0_1_1_argbuf,Pointer_QTree_Bool),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet11_1_5MQVal_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [5:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet0_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet11_1_5MQVal_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet3_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0])};
  assign go_8_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r,
          lizzieLet11_1_5MQVal_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet0_1_1_argbuf_r} = (go_8_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTmain_mask_Bool) : (go_8_goMux_choice_2,C6) [(lizzieLet11_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (sc_0_9_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (lizzieLet11_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTmain_mask_Bool),
                                                              (lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf,Pointer_CTmain_mask_Bool)] > (scfarg_0_1_goMux_mux,Pointer_CTmain_mask_Bool) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [5:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet11_1_6MQNone_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   sc_0_9_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet11_1_6MQVal_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_d};
      3'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0])};
  assign go_8_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_r,
          lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_r,
          lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_r,
          lizzieLet11_1_6MQVal_1_argbuf_r,
          sc_0_9_1_argbuf_r,
          lizzieLet11_1_6MQNone_1_argbuf_r} = (go_8_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               6'd0);
  
  /* destruct (Ty MaskQTree,
          Dcon MQNode) : (lizzieLet11_1_1MQNode,MaskQTree) > [(q1a8s_destruct,Pointer_MaskQTree),
                                                              (q2a8t_destruct,Pointer_MaskQTree),
                                                              (q3a8u_destruct,Pointer_MaskQTree),
                                                              (q4a8v_destruct,Pointer_MaskQTree)] */
  logic [3:0] lizzieLet11_1_1MQNode_emitted;
  logic [3:0] lizzieLet11_1_1MQNode_done;
  assign q1a8s_destruct_d = {lizzieLet11_1_1MQNode_d[18:3],
                             (lizzieLet11_1_1MQNode_d[0] && (! lizzieLet11_1_1MQNode_emitted[0]))};
  assign q2a8t_destruct_d = {lizzieLet11_1_1MQNode_d[34:19],
                             (lizzieLet11_1_1MQNode_d[0] && (! lizzieLet11_1_1MQNode_emitted[1]))};
  assign q3a8u_destruct_d = {lizzieLet11_1_1MQNode_d[50:35],
                             (lizzieLet11_1_1MQNode_d[0] && (! lizzieLet11_1_1MQNode_emitted[2]))};
  assign q4a8v_destruct_d = {lizzieLet11_1_1MQNode_d[66:51],
                             (lizzieLet11_1_1MQNode_d[0] && (! lizzieLet11_1_1MQNode_emitted[3]))};
  assign lizzieLet11_1_1MQNode_done = (lizzieLet11_1_1MQNode_emitted | ({q4a8v_destruct_d[0],
                                                                         q3a8u_destruct_d[0],
                                                                         q2a8t_destruct_d[0],
                                                                         q1a8s_destruct_d[0]} & {q4a8v_destruct_r,
                                                                                                 q3a8u_destruct_r,
                                                                                                 q2a8t_destruct_r,
                                                                                                 q1a8s_destruct_r}));
  assign lizzieLet11_1_1MQNode_r = (& lizzieLet11_1_1MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1MQNode_emitted <= 4'd0;
    else
      lizzieLet11_1_1MQNode_emitted <= (lizzieLet11_1_1MQNode_r ? 4'd0 :
                                        lizzieLet11_1_1MQNode_done);
  
  /* demux (Ty MaskQTree,
       Ty MaskQTree) : (lizzieLet11_1_2,MaskQTree) (lizzieLet11_1_1,MaskQTree) > [(_68,MaskQTree),
                                                                                  (_67,MaskQTree),
                                                                                  (lizzieLet11_1_1MQNode,MaskQTree)] */
  logic [2:0] lizzieLet11_1_1_onehotd;
  always_comb
    if ((lizzieLet11_1_2_d[0] && lizzieLet11_1_1_d[0]))
      unique case (lizzieLet11_1_2_d[2:1])
        2'd0: lizzieLet11_1_1_onehotd = 3'd1;
        2'd1: lizzieLet11_1_1_onehotd = 3'd2;
        2'd2: lizzieLet11_1_1_onehotd = 3'd4;
        default: lizzieLet11_1_1_onehotd = 3'd0;
      endcase
    else lizzieLet11_1_1_onehotd = 3'd0;
  assign _68_d = {lizzieLet11_1_1_d[66:1],
                  lizzieLet11_1_1_onehotd[0]};
  assign _67_d = {lizzieLet11_1_1_d[66:1],
                  lizzieLet11_1_1_onehotd[1]};
  assign lizzieLet11_1_1MQNode_d = {lizzieLet11_1_1_d[66:1],
                                    lizzieLet11_1_1_onehotd[2]};
  assign lizzieLet11_1_1_r = (| (lizzieLet11_1_1_onehotd & {lizzieLet11_1_1MQNode_r,
                                                            _67_r,
                                                            _68_r}));
  assign lizzieLet11_1_2_r = lizzieLet11_1_1_r;
  
  /* demux (Ty MaskQTree,
       Ty Go) : (lizzieLet11_1_3,MaskQTree) (go_5_goMux_data,Go) > [(lizzieLet11_1_3MQNone,Go),
                                                                    (lizzieLet11_1_3MQVal,Go),
                                                                    (lizzieLet11_1_3MQNode,Go)] */
  logic [2:0] go_5_goMux_data_onehotd;
  always_comb
    if ((lizzieLet11_1_3_d[0] && go_5_goMux_data_d[0]))
      unique case (lizzieLet11_1_3_d[2:1])
        2'd0: go_5_goMux_data_onehotd = 3'd1;
        2'd1: go_5_goMux_data_onehotd = 3'd2;
        2'd2: go_5_goMux_data_onehotd = 3'd4;
        default: go_5_goMux_data_onehotd = 3'd0;
      endcase
    else go_5_goMux_data_onehotd = 3'd0;
  assign lizzieLet11_1_3MQNone_d = go_5_goMux_data_onehotd[0];
  assign lizzieLet11_1_3MQVal_d = go_5_goMux_data_onehotd[1];
  assign lizzieLet11_1_3MQNode_d = go_5_goMux_data_onehotd[2];
  assign go_5_goMux_data_r = (| (go_5_goMux_data_onehotd & {lizzieLet11_1_3MQNode_r,
                                                            lizzieLet11_1_3MQVal_r,
                                                            lizzieLet11_1_3MQNone_r}));
  assign lizzieLet11_1_3_r = go_5_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet11_1_3MQNone,Go) > [(lizzieLet11_1_3MQNone_1,Go),
                                             (lizzieLet11_1_3MQNone_2,Go)] */
  logic [1:0] lizzieLet11_1_3MQNone_emitted;
  logic [1:0] lizzieLet11_1_3MQNone_done;
  assign lizzieLet11_1_3MQNone_1_d = (lizzieLet11_1_3MQNone_d[0] && (! lizzieLet11_1_3MQNone_emitted[0]));
  assign lizzieLet11_1_3MQNone_2_d = (lizzieLet11_1_3MQNone_d[0] && (! lizzieLet11_1_3MQNone_emitted[1]));
  assign lizzieLet11_1_3MQNone_done = (lizzieLet11_1_3MQNone_emitted | ({lizzieLet11_1_3MQNone_2_d[0],
                                                                         lizzieLet11_1_3MQNone_1_d[0]} & {lizzieLet11_1_3MQNone_2_r,
                                                                                                          lizzieLet11_1_3MQNone_1_r}));
  assign lizzieLet11_1_3MQNone_r = (& lizzieLet11_1_3MQNone_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQNone_emitted <= 2'd0;
    else
      lizzieLet11_1_3MQNone_emitted <= (lizzieLet11_1_3MQNone_r ? 2'd0 :
                                        lizzieLet11_1_3MQNone_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet11_1_3MQNone_1,Go)] > (lizzieLet11_1_3MQNone_1QNone_Bool,QTree_Bool) */
  assign lizzieLet11_1_3MQNone_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet11_1_3MQNone_1_d[0]}), lizzieLet11_1_3MQNone_1_d);
  assign {lizzieLet11_1_3MQNone_1_r} = {1 {(lizzieLet11_1_3MQNone_1QNone_Bool_r && lizzieLet11_1_3MQNone_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_3MQNone_1QNone_Bool,QTree_Bool) > (lizzieLet12_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d;
  logic lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_r;
  assign lizzieLet11_1_3MQNone_1QNone_Bool_r = ((! lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d[0]) || lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet11_1_3MQNone_1QNone_Bool_r)
        lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d <= lizzieLet11_1_3MQNone_1QNone_Bool_d;
  QTree_Bool_t lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf;
  assign lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_r = (! lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf[0] ? lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf :
                                   lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf[0]))
        lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf[0])))
        lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_buf <= lizzieLet11_1_3MQNone_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_3MQNone_2,Go) > (lizzieLet11_1_3MQNone_2_argbuf,Go) */
  Go_t lizzieLet11_1_3MQNone_2_bufchan_d;
  logic lizzieLet11_1_3MQNone_2_bufchan_r;
  assign lizzieLet11_1_3MQNone_2_r = ((! lizzieLet11_1_3MQNone_2_bufchan_d[0]) || lizzieLet11_1_3MQNone_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQNone_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_3MQNone_2_r)
        lizzieLet11_1_3MQNone_2_bufchan_d <= lizzieLet11_1_3MQNone_2_d;
  Go_t lizzieLet11_1_3MQNone_2_bufchan_buf;
  assign lizzieLet11_1_3MQNone_2_bufchan_r = (! lizzieLet11_1_3MQNone_2_bufchan_buf[0]);
  assign lizzieLet11_1_3MQNone_2_argbuf_d = (lizzieLet11_1_3MQNone_2_bufchan_buf[0] ? lizzieLet11_1_3MQNone_2_bufchan_buf :
                                             lizzieLet11_1_3MQNone_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQNone_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_3MQNone_2_argbuf_r && lizzieLet11_1_3MQNone_2_bufchan_buf[0]))
        lizzieLet11_1_3MQNone_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_3MQNone_2_argbuf_r) && (! lizzieLet11_1_3MQNone_2_bufchan_buf[0])))
        lizzieLet11_1_3MQNone_2_bufchan_buf <= lizzieLet11_1_3MQNone_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet11_1_3MQNone_2_argbuf,Go),
                           (lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf,Go),
                           (lizzieLet11_1_3MQVal_1_argbuf,Go),
                           (lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf,Go),
                           (lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf,Go),
                           (lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf,Go)] > (go_8_goMux_choice,C6) (go_8_goMux_data,Go) */
  logic [5:0] lizzieLet11_1_3MQNone_2_argbuf_select_d;
  assign lizzieLet11_1_3MQNone_2_argbuf_select_d = ((| lizzieLet11_1_3MQNone_2_argbuf_select_q) ? lizzieLet11_1_3MQNone_2_argbuf_select_q :
                                                    (lizzieLet11_1_3MQNone_2_argbuf_d[0] ? 6'd1 :
                                                     (lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_d[0] ? 6'd2 :
                                                      (lizzieLet11_1_3MQVal_1_argbuf_d[0] ? 6'd4 :
                                                       (lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_d[0] ? 6'd8 :
                                                        (lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_d[0] ? 6'd16 :
                                                         (lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_d[0] ? 6'd32 :
                                                          6'd0)))))));
  logic [5:0] lizzieLet11_1_3MQNone_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_3MQNone_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet11_1_3MQNone_2_argbuf_select_q <= (lizzieLet11_1_3MQNone_2_argbuf_done ? 6'd0 :
                                                  lizzieLet11_1_3MQNone_2_argbuf_select_d);
  logic [1:0] lizzieLet11_1_3MQNone_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQNone_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_3MQNone_2_argbuf_emit_q <= (lizzieLet11_1_3MQNone_2_argbuf_done ? 2'd0 :
                                                lizzieLet11_1_3MQNone_2_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_3MQNone_2_argbuf_emit_d;
  assign lizzieLet11_1_3MQNone_2_argbuf_emit_d = (lizzieLet11_1_3MQNone_2_argbuf_emit_q | ({go_8_goMux_choice_d[0],
                                                                                            go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                                     go_8_goMux_data_r}));
  logic lizzieLet11_1_3MQNone_2_argbuf_done;
  assign lizzieLet11_1_3MQNone_2_argbuf_done = (& lizzieLet11_1_3MQNone_2_argbuf_emit_d);
  assign {lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_r,
          lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_r,
          lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_r,
          lizzieLet11_1_3MQVal_1_argbuf_r,
          lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_r,
          lizzieLet11_1_3MQNone_2_argbuf_r} = (lizzieLet11_1_3MQNone_2_argbuf_done ? lizzieLet11_1_3MQNone_2_argbuf_select_d :
                                               6'd0);
  assign go_8_goMux_data_d = ((lizzieLet11_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet11_1_3MQNone_2_argbuf_d :
                              ((lizzieLet11_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_d :
                               ((lizzieLet11_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet11_1_3MQVal_1_argbuf_d :
                                ((lizzieLet11_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_d :
                                 ((lizzieLet11_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_d :
                                  ((lizzieLet11_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[0])) ? lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_d :
                                   1'd0))))));
  assign go_8_goMux_choice_d = ((lizzieLet11_1_3MQNone_2_argbuf_select_d[0] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                ((lizzieLet11_1_3MQNone_2_argbuf_select_d[1] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                 ((lizzieLet11_1_3MQNone_2_argbuf_select_d[2] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                  ((lizzieLet11_1_3MQNone_2_argbuf_select_d[3] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                   ((lizzieLet11_1_3MQNone_2_argbuf_select_d[4] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                    ((lizzieLet11_1_3MQNone_2_argbuf_select_d[5] && (! lizzieLet11_1_3MQNone_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                     {3'd0, 1'd0}))))));
  
  /* buf (Ty Go) : (lizzieLet11_1_3MQVal,Go) > (lizzieLet11_1_3MQVal_1_argbuf,Go) */
  Go_t lizzieLet11_1_3MQVal_bufchan_d;
  logic lizzieLet11_1_3MQVal_bufchan_r;
  assign lizzieLet11_1_3MQVal_r = ((! lizzieLet11_1_3MQVal_bufchan_d[0]) || lizzieLet11_1_3MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQVal_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_3MQVal_r)
        lizzieLet11_1_3MQVal_bufchan_d <= lizzieLet11_1_3MQVal_d;
  Go_t lizzieLet11_1_3MQVal_bufchan_buf;
  assign lizzieLet11_1_3MQVal_bufchan_r = (! lizzieLet11_1_3MQVal_bufchan_buf[0]);
  assign lizzieLet11_1_3MQVal_1_argbuf_d = (lizzieLet11_1_3MQVal_bufchan_buf[0] ? lizzieLet11_1_3MQVal_bufchan_buf :
                                            lizzieLet11_1_3MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_3MQVal_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_3MQVal_1_argbuf_r && lizzieLet11_1_3MQVal_bufchan_buf[0]))
        lizzieLet11_1_3MQVal_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_3MQVal_1_argbuf_r) && (! lizzieLet11_1_3MQVal_bufchan_buf[0])))
        lizzieLet11_1_3MQVal_bufchan_buf <= lizzieLet11_1_3MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty QTree_Bool) : (lizzieLet11_1_4,MaskQTree) (readPointer_QTree_Boolma8q_1_argbuf_rwb,QTree_Bool) > [(_66,QTree_Bool),
                                                                                                            (_65,QTree_Bool),
                                                                                                            (lizzieLet11_1_4MQNode,QTree_Bool)] */
  logic [2:0] readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet11_1_4_d[0] && readPointer_QTree_Boolma8q_1_argbuf_rwb_d[0]))
      unique case (lizzieLet11_1_4_d[2:1])
        2'd0: readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd = 3'd1;
        2'd1: readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd = 3'd2;
        2'd2: readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd = 3'd4;
        default: readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd = 3'd0;
      endcase
    else readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd = 3'd0;
  assign _66_d = {readPointer_QTree_Boolma8q_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd[0]};
  assign _65_d = {readPointer_QTree_Boolma8q_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet11_1_4MQNode_d = {readPointer_QTree_Boolma8q_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd[2]};
  assign readPointer_QTree_Boolma8q_1_argbuf_rwb_r = (| (readPointer_QTree_Boolma8q_1_argbuf_rwb_onehotd & {lizzieLet11_1_4MQNode_r,
                                                                                                            _65_r,
                                                                                                            _66_r}));
  assign lizzieLet11_1_4_r = readPointer_QTree_Boolma8q_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet11_1_4MQNode,QTree_Bool) > [(lizzieLet11_1_4MQNode_1,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_2,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_3,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_4,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_5,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_6,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_7,QTree_Bool),
                                                             (lizzieLet11_1_4MQNode_8,QTree_Bool)] */
  logic [7:0] lizzieLet11_1_4MQNode_emitted;
  logic [7:0] lizzieLet11_1_4MQNode_done;
  assign lizzieLet11_1_4MQNode_1_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[0]))};
  assign lizzieLet11_1_4MQNode_2_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[1]))};
  assign lizzieLet11_1_4MQNode_3_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[2]))};
  assign lizzieLet11_1_4MQNode_4_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[3]))};
  assign lizzieLet11_1_4MQNode_5_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[4]))};
  assign lizzieLet11_1_4MQNode_6_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[5]))};
  assign lizzieLet11_1_4MQNode_7_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[6]))};
  assign lizzieLet11_1_4MQNode_8_d = {lizzieLet11_1_4MQNode_d[66:1],
                                      (lizzieLet11_1_4MQNode_d[0] && (! lizzieLet11_1_4MQNode_emitted[7]))};
  assign lizzieLet11_1_4MQNode_done = (lizzieLet11_1_4MQNode_emitted | ({lizzieLet11_1_4MQNode_8_d[0],
                                                                         lizzieLet11_1_4MQNode_7_d[0],
                                                                         lizzieLet11_1_4MQNode_6_d[0],
                                                                         lizzieLet11_1_4MQNode_5_d[0],
                                                                         lizzieLet11_1_4MQNode_4_d[0],
                                                                         lizzieLet11_1_4MQNode_3_d[0],
                                                                         lizzieLet11_1_4MQNode_2_d[0],
                                                                         lizzieLet11_1_4MQNode_1_d[0]} & {lizzieLet11_1_4MQNode_8_r,
                                                                                                          lizzieLet11_1_4MQNode_7_r,
                                                                                                          lizzieLet11_1_4MQNode_6_r,
                                                                                                          lizzieLet11_1_4MQNode_5_r,
                                                                                                          lizzieLet11_1_4MQNode_4_r,
                                                                                                          lizzieLet11_1_4MQNode_3_r,
                                                                                                          lizzieLet11_1_4MQNode_2_r,
                                                                                                          lizzieLet11_1_4MQNode_1_r}));
  assign lizzieLet11_1_4MQNode_r = (& lizzieLet11_1_4MQNode_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_4MQNode_emitted <= 8'd0;
    else
      lizzieLet11_1_4MQNode_emitted <= (lizzieLet11_1_4MQNode_r ? 8'd0 :
                                        lizzieLet11_1_4MQNode_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet11_1_4MQNode_1QNode_Bool,QTree_Bool) > [(t1a8x_destruct,Pointer_QTree_Bool),
                                                                               (t2a8y_destruct,Pointer_QTree_Bool),
                                                                               (t3a8z_destruct,Pointer_QTree_Bool),
                                                                               (t4a8A_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet11_1_4MQNode_1QNode_Bool_emitted;
  logic [3:0] lizzieLet11_1_4MQNode_1QNode_Bool_done;
  assign t1a8x_destruct_d = {lizzieLet11_1_4MQNode_1QNode_Bool_d[18:3],
                             (lizzieLet11_1_4MQNode_1QNode_Bool_d[0] && (! lizzieLet11_1_4MQNode_1QNode_Bool_emitted[0]))};
  assign t2a8y_destruct_d = {lizzieLet11_1_4MQNode_1QNode_Bool_d[34:19],
                             (lizzieLet11_1_4MQNode_1QNode_Bool_d[0] && (! lizzieLet11_1_4MQNode_1QNode_Bool_emitted[1]))};
  assign t3a8z_destruct_d = {lizzieLet11_1_4MQNode_1QNode_Bool_d[50:35],
                             (lizzieLet11_1_4MQNode_1QNode_Bool_d[0] && (! lizzieLet11_1_4MQNode_1QNode_Bool_emitted[2]))};
  assign t4a8A_destruct_d = {lizzieLet11_1_4MQNode_1QNode_Bool_d[66:51],
                             (lizzieLet11_1_4MQNode_1QNode_Bool_d[0] && (! lizzieLet11_1_4MQNode_1QNode_Bool_emitted[3]))};
  assign lizzieLet11_1_4MQNode_1QNode_Bool_done = (lizzieLet11_1_4MQNode_1QNode_Bool_emitted | ({t4a8A_destruct_d[0],
                                                                                                 t3a8z_destruct_d[0],
                                                                                                 t2a8y_destruct_d[0],
                                                                                                 t1a8x_destruct_d[0]} & {t4a8A_destruct_r,
                                                                                                                         t3a8z_destruct_r,
                                                                                                                         t2a8y_destruct_r,
                                                                                                                         t1a8x_destruct_r}));
  assign lizzieLet11_1_4MQNode_1QNode_Bool_r = (& lizzieLet11_1_4MQNode_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet11_1_4MQNode_1QNode_Bool_emitted <= (lizzieLet11_1_4MQNode_1QNode_Bool_r ? 4'd0 :
                                                    lizzieLet11_1_4MQNode_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet11_1_4MQNode_2,QTree_Bool) (lizzieLet11_1_4MQNode_1,QTree_Bool) > [(_64,QTree_Bool),
                                                                                                     (_63,QTree_Bool),
                                                                                                     (lizzieLet11_1_4MQNode_1QNode_Bool,QTree_Bool),
                                                                                                     (_62,QTree_Bool)] */
  logic [3:0] lizzieLet11_1_4MQNode_1_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_2_d[0] && lizzieLet11_1_4MQNode_1_d[0]))
      unique case (lizzieLet11_1_4MQNode_2_d[2:1])
        2'd0: lizzieLet11_1_4MQNode_1_onehotd = 4'd1;
        2'd1: lizzieLet11_1_4MQNode_1_onehotd = 4'd2;
        2'd2: lizzieLet11_1_4MQNode_1_onehotd = 4'd4;
        2'd3: lizzieLet11_1_4MQNode_1_onehotd = 4'd8;
        default: lizzieLet11_1_4MQNode_1_onehotd = 4'd0;
      endcase
    else lizzieLet11_1_4MQNode_1_onehotd = 4'd0;
  assign _64_d = {lizzieLet11_1_4MQNode_1_d[66:1],
                  lizzieLet11_1_4MQNode_1_onehotd[0]};
  assign _63_d = {lizzieLet11_1_4MQNode_1_d[66:1],
                  lizzieLet11_1_4MQNode_1_onehotd[1]};
  assign lizzieLet11_1_4MQNode_1QNode_Bool_d = {lizzieLet11_1_4MQNode_1_d[66:1],
                                                lizzieLet11_1_4MQNode_1_onehotd[2]};
  assign _62_d = {lizzieLet11_1_4MQNode_1_d[66:1],
                  lizzieLet11_1_4MQNode_1_onehotd[3]};
  assign lizzieLet11_1_4MQNode_1_r = (| (lizzieLet11_1_4MQNode_1_onehotd & {_62_r,
                                                                            lizzieLet11_1_4MQNode_1QNode_Bool_r,
                                                                            _63_r,
                                                                            _64_r}));
  assign lizzieLet11_1_4MQNode_2_r = lizzieLet11_1_4MQNode_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet11_1_4MQNode_3,QTree_Bool) (lizzieLet11_1_3MQNode,Go) > [(lizzieLet11_1_4MQNode_3QNone_Bool,Go),
                                                                                   (lizzieLet11_1_4MQNode_3QVal_Bool,Go),
                                                                                   (lizzieLet11_1_4MQNode_3QNode_Bool,Go),
                                                                                   (lizzieLet11_1_4MQNode_3QError_Bool,Go)] */
  logic [3:0] lizzieLet11_1_3MQNode_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_3_d[0] && lizzieLet11_1_3MQNode_d[0]))
      unique case (lizzieLet11_1_4MQNode_3_d[2:1])
        2'd0: lizzieLet11_1_3MQNode_onehotd = 4'd1;
        2'd1: lizzieLet11_1_3MQNode_onehotd = 4'd2;
        2'd2: lizzieLet11_1_3MQNode_onehotd = 4'd4;
        2'd3: lizzieLet11_1_3MQNode_onehotd = 4'd8;
        default: lizzieLet11_1_3MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet11_1_3MQNode_onehotd = 4'd0;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_d = lizzieLet11_1_3MQNode_onehotd[0];
  assign lizzieLet11_1_4MQNode_3QVal_Bool_d = lizzieLet11_1_3MQNode_onehotd[1];
  assign lizzieLet11_1_4MQNode_3QNode_Bool_d = lizzieLet11_1_3MQNode_onehotd[2];
  assign lizzieLet11_1_4MQNode_3QError_Bool_d = lizzieLet11_1_3MQNode_onehotd[3];
  assign lizzieLet11_1_3MQNode_r = (| (lizzieLet11_1_3MQNode_onehotd & {lizzieLet11_1_4MQNode_3QError_Bool_r,
                                                                        lizzieLet11_1_4MQNode_3QNode_Bool_r,
                                                                        lizzieLet11_1_4MQNode_3QVal_Bool_r,
                                                                        lizzieLet11_1_4MQNode_3QNone_Bool_r}));
  assign lizzieLet11_1_4MQNode_3_r = lizzieLet11_1_3MQNode_r;
  
  /* fork (Ty Go) : (lizzieLet11_1_4MQNode_3QError_Bool,Go) > [(lizzieLet11_1_4MQNode_3QError_Bool_1,Go),
                                                          (lizzieLet11_1_4MQNode_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet11_1_4MQNode_3QError_Bool_emitted;
  logic [1:0] lizzieLet11_1_4MQNode_3QError_Bool_done;
  assign lizzieLet11_1_4MQNode_3QError_Bool_1_d = (lizzieLet11_1_4MQNode_3QError_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QError_Bool_emitted[0]));
  assign lizzieLet11_1_4MQNode_3QError_Bool_2_d = (lizzieLet11_1_4MQNode_3QError_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QError_Bool_emitted[1]));
  assign lizzieLet11_1_4MQNode_3QError_Bool_done = (lizzieLet11_1_4MQNode_3QError_Bool_emitted | ({lizzieLet11_1_4MQNode_3QError_Bool_2_d[0],
                                                                                                   lizzieLet11_1_4MQNode_3QError_Bool_1_d[0]} & {lizzieLet11_1_4MQNode_3QError_Bool_2_r,
                                                                                                                                                 lizzieLet11_1_4MQNode_3QError_Bool_1_r}));
  assign lizzieLet11_1_4MQNode_3QError_Bool_r = (& lizzieLet11_1_4MQNode_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_4MQNode_3QError_Bool_emitted <= (lizzieLet11_1_4MQNode_3QError_Bool_r ? 2'd0 :
                                                     lizzieLet11_1_4MQNode_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet11_1_4MQNode_3QError_Bool_1,Go)] > (lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet11_1_4MQNode_3QError_Bool_1_d[0]}), lizzieLet11_1_4MQNode_3QError_Bool_1_d);
  assign {lizzieLet11_1_4MQNode_3QError_Bool_1_r} = {1 {(lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_r && lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet17_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_r = ((! lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_r)
        lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4MQNode_3QError_Bool_2,Go) > (lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QError_Bool_2_r = ((! lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4MQNode_3QError_Bool_2_r)
        lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d <= lizzieLet11_1_4MQNode_3QError_Bool_2_d;
  Go_t lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_r = (! lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_d = (lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf :
                                                          lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_r && lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4MQNode_3QError_Bool_2_argbuf_r) && (! lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_buf <= lizzieLet11_1_4MQNode_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4MQNode_3QNode_Bool,Go) > (lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QNode_Bool_r = ((! lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4MQNode_3QNode_Bool_r)
        lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d <= lizzieLet11_1_4MQNode_3QNode_Bool_d;
  Go_t lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_d = (lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf :
                                                         lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_r && lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4MQNode_3QNode_Bool_1_argbuf_r) && (! lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_3QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet11_1_4MQNode_3QNone_Bool,Go) > [(lizzieLet11_1_4MQNode_3QNone_Bool_1,Go),
                                                         (lizzieLet11_1_4MQNode_3QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet11_1_4MQNode_3QNone_Bool_emitted;
  logic [1:0] lizzieLet11_1_4MQNode_3QNone_Bool_done;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_1_d = (lizzieLet11_1_4MQNode_3QNone_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QNone_Bool_emitted[0]));
  assign lizzieLet11_1_4MQNode_3QNone_Bool_2_d = (lizzieLet11_1_4MQNode_3QNone_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QNone_Bool_emitted[1]));
  assign lizzieLet11_1_4MQNode_3QNone_Bool_done = (lizzieLet11_1_4MQNode_3QNone_Bool_emitted | ({lizzieLet11_1_4MQNode_3QNone_Bool_2_d[0],
                                                                                                 lizzieLet11_1_4MQNode_3QNone_Bool_1_d[0]} & {lizzieLet11_1_4MQNode_3QNone_Bool_2_r,
                                                                                                                                              lizzieLet11_1_4MQNode_3QNone_Bool_1_r}));
  assign lizzieLet11_1_4MQNode_3QNone_Bool_r = (& lizzieLet11_1_4MQNode_3QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_4MQNode_3QNone_Bool_emitted <= (lizzieLet11_1_4MQNode_3QNone_Bool_r ? 2'd0 :
                                                    lizzieLet11_1_4MQNode_3QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet11_1_4MQNode_3QNone_Bool_1,Go)] > (lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet11_1_4MQNode_3QNone_Bool_1_d[0]}), lizzieLet11_1_4MQNode_3QNone_Bool_1_d);
  assign {lizzieLet11_1_4MQNode_3QNone_Bool_1_r} = {1 {(lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_r && lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet14_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_r = ((! lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_r)
        lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf :
                                   lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_3QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4MQNode_3QNone_Bool_2,Go) > (lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_2_r = ((! lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4MQNode_3QNone_Bool_2_r)
        lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d <= lizzieLet11_1_4MQNode_3QNone_Bool_2_d;
  Go_t lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_r = (! lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_d = (lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf :
                                                         lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_r && lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4MQNode_3QNone_Bool_2_argbuf_r) && (! lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_buf <= lizzieLet11_1_4MQNode_3QNone_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet11_1_4MQNode_3QVal_Bool,Go) > [(lizzieLet11_1_4MQNode_3QVal_Bool_1,Go),
                                                        (lizzieLet11_1_4MQNode_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet11_1_4MQNode_3QVal_Bool_emitted;
  logic [1:0] lizzieLet11_1_4MQNode_3QVal_Bool_done;
  assign lizzieLet11_1_4MQNode_3QVal_Bool_1_d = (lizzieLet11_1_4MQNode_3QVal_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QVal_Bool_emitted[0]));
  assign lizzieLet11_1_4MQNode_3QVal_Bool_2_d = (lizzieLet11_1_4MQNode_3QVal_Bool_d[0] && (! lizzieLet11_1_4MQNode_3QVal_Bool_emitted[1]));
  assign lizzieLet11_1_4MQNode_3QVal_Bool_done = (lizzieLet11_1_4MQNode_3QVal_Bool_emitted | ({lizzieLet11_1_4MQNode_3QVal_Bool_2_d[0],
                                                                                               lizzieLet11_1_4MQNode_3QVal_Bool_1_d[0]} & {lizzieLet11_1_4MQNode_3QVal_Bool_2_r,
                                                                                                                                           lizzieLet11_1_4MQNode_3QVal_Bool_1_r}));
  assign lizzieLet11_1_4MQNode_3QVal_Bool_r = (& lizzieLet11_1_4MQNode_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet11_1_4MQNode_3QVal_Bool_emitted <= (lizzieLet11_1_4MQNode_3QVal_Bool_r ? 2'd0 :
                                                   lizzieLet11_1_4MQNode_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet11_1_4MQNode_3QVal_Bool_1,Go)] > (lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet11_1_4MQNode_3QVal_Bool_1_d[0]}), lizzieLet11_1_4MQNode_3QVal_Bool_1_d);
  assign {lizzieLet11_1_4MQNode_3QVal_Bool_1_r} = {1 {(lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_r && lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet15_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_r = ((! lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                  1'd0};
    else
      if (lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_r)
        lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                    1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet11_1_4MQNode_3QVal_Bool_2,Go) > (lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d;
  logic lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_r;
  assign lizzieLet11_1_4MQNode_3QVal_Bool_2_r = ((! lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d[0]) || lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet11_1_4MQNode_3QVal_Bool_2_r)
        lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d <= lizzieLet11_1_4MQNode_3QVal_Bool_2_d;
  Go_t lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_r = (! lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_d = (lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf :
                                                        lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_r && lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet11_1_4MQNode_3QVal_Bool_2_argbuf_r) && (! lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_buf <= lizzieLet11_1_4MQNode_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_4MQNode_4,QTree_Bool) (lizzieLet11_1_6MQNode,Pointer_CTmain_mask_Bool) > [(lizzieLet11_1_4MQNode_4QNone_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                               (lizzieLet11_1_4MQNode_4QVal_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                               (lizzieLet11_1_4MQNode_4QNode_Bool,Pointer_CTmain_mask_Bool),
                                                                                                                               (lizzieLet11_1_4MQNode_4QError_Bool,Pointer_CTmain_mask_Bool)] */
  logic [3:0] lizzieLet11_1_6MQNode_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_4_d[0] && lizzieLet11_1_6MQNode_d[0]))
      unique case (lizzieLet11_1_4MQNode_4_d[2:1])
        2'd0: lizzieLet11_1_6MQNode_onehotd = 4'd1;
        2'd1: lizzieLet11_1_6MQNode_onehotd = 4'd2;
        2'd2: lizzieLet11_1_6MQNode_onehotd = 4'd4;
        2'd3: lizzieLet11_1_6MQNode_onehotd = 4'd8;
        default: lizzieLet11_1_6MQNode_onehotd = 4'd0;
      endcase
    else lizzieLet11_1_6MQNode_onehotd = 4'd0;
  assign lizzieLet11_1_4MQNode_4QNone_Bool_d = {lizzieLet11_1_6MQNode_d[16:1],
                                                lizzieLet11_1_6MQNode_onehotd[0]};
  assign lizzieLet11_1_4MQNode_4QVal_Bool_d = {lizzieLet11_1_6MQNode_d[16:1],
                                               lizzieLet11_1_6MQNode_onehotd[1]};
  assign lizzieLet11_1_4MQNode_4QNode_Bool_d = {lizzieLet11_1_6MQNode_d[16:1],
                                                lizzieLet11_1_6MQNode_onehotd[2]};
  assign lizzieLet11_1_4MQNode_4QError_Bool_d = {lizzieLet11_1_6MQNode_d[16:1],
                                                 lizzieLet11_1_6MQNode_onehotd[3]};
  assign lizzieLet11_1_6MQNode_r = (| (lizzieLet11_1_6MQNode_onehotd & {lizzieLet11_1_4MQNode_4QError_Bool_r,
                                                                        lizzieLet11_1_4MQNode_4QNode_Bool_r,
                                                                        lizzieLet11_1_4MQNode_4QVal_Bool_r,
                                                                        lizzieLet11_1_4MQNode_4QNone_Bool_r}));
  assign lizzieLet11_1_4MQNode_4_r = lizzieLet11_1_6MQNode_r;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_4MQNode_4QError_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_4QError_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_4QError_Bool_r = ((! lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_4MQNode_4QError_Bool_r)
        lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d <= lizzieLet11_1_4MQNode_4QError_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_4QError_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_d = (lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf :
                                                          lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_r && lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_4MQNode_4QError_Bool_1_argbuf_r) && (! lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_4QError_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool3) : [(lizzieLet11_1_4MQNode_4QNode_Bool,Pointer_CTmain_mask_Bool),
                                     (t1a8x_destruct,Pointer_QTree_Bool),
                                     (lizzieLet11_1_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                     (t2a8y_destruct,Pointer_QTree_Bool),
                                     (lizzieLet11_1_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                     (t3a8z_destruct,Pointer_QTree_Bool),
                                     (lizzieLet11_1_4MQNode_7QNode_Bool,Pointer_MaskQTree)] > (lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3,CTmain_mask_Bool) */
  assign lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d = Lcall_main_mask_Bool3_dc((& {lizzieLet11_1_4MQNode_4QNode_Bool_d[0],
                                                                                                                                                                                                                                 t1a8x_destruct_d[0],
                                                                                                                                                                                                                                 lizzieLet11_1_4MQNode_5QNode_Bool_d[0],
                                                                                                                                                                                                                                 t2a8y_destruct_d[0],
                                                                                                                                                                                                                                 lizzieLet11_1_4MQNode_6QNode_Bool_d[0],
                                                                                                                                                                                                                                 t3a8z_destruct_d[0],
                                                                                                                                                                                                                                 lizzieLet11_1_4MQNode_7QNode_Bool_d[0]}), lizzieLet11_1_4MQNode_4QNode_Bool_d, t1a8x_destruct_d, lizzieLet11_1_4MQNode_5QNode_Bool_d, t2a8y_destruct_d, lizzieLet11_1_4MQNode_6QNode_Bool_d, t3a8z_destruct_d, lizzieLet11_1_4MQNode_7QNode_Bool_d);
  assign {lizzieLet11_1_4MQNode_4QNode_Bool_r,
          t1a8x_destruct_r,
          lizzieLet11_1_4MQNode_5QNode_Bool_r,
          t2a8y_destruct_r,
          lizzieLet11_1_4MQNode_6QNode_Bool_r,
          t3a8z_destruct_r,
          lizzieLet11_1_4MQNode_7QNode_Bool_r} = {7 {(lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r && lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3,CTmain_mask_Bool) > (lizzieLet16_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d;
  logic lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r;
  assign lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r = ((! lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d[0]) || lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d <= {115'd0,
                                                                                                                                                                                                           1'd0};
    else
      if (lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_r)
        lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d <= lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_d;
  CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf;
  assign lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_r = (! lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0] ? lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf :
                                   lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                             1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                               1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_buf <= lizzieLet11_1_4MQNode_4QNode_Bool_1t1a8x_1lizzieLet11_1_4MQNode_5QNode_Bool_1t2a8y_1lizzieLet11_1_4MQNode_6QNode_Bool_1t3a8z_1lizzieLet11_1_4MQNode_7QNode_Bool_1Lcall_main_mask_Bool3_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_4MQNode_4QNone_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_4QNone_Bool_r = ((! lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_4MQNode_4QNone_Bool_r)
        lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d <= lizzieLet11_1_4MQNode_4QNone_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_d = (lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf :
                                                         lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_r && lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_4MQNode_4QNone_Bool_1_argbuf_r) && (! lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_4MQNode_4QVal_Bool,Pointer_CTmain_mask_Bool) > (lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_4QVal_Bool_r = ((! lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_4MQNode_4QVal_Bool_r)
        lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d <= lizzieLet11_1_4MQNode_4QVal_Bool_d;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_d = (lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf :
                                                        lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_r && lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_4MQNode_4QVal_Bool_1_argbuf_r) && (! lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet11_1_4MQNode_5,QTree_Bool) (q1a8s_destruct,Pointer_MaskQTree) > [(_61,Pointer_MaskQTree),
                                                                                                          (_60,Pointer_MaskQTree),
                                                                                                          (lizzieLet11_1_4MQNode_5QNode_Bool,Pointer_MaskQTree),
                                                                                                          (_59,Pointer_MaskQTree)] */
  logic [3:0] q1a8s_destruct_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_5_d[0] && q1a8s_destruct_d[0]))
      unique case (lizzieLet11_1_4MQNode_5_d[2:1])
        2'd0: q1a8s_destruct_onehotd = 4'd1;
        2'd1: q1a8s_destruct_onehotd = 4'd2;
        2'd2: q1a8s_destruct_onehotd = 4'd4;
        2'd3: q1a8s_destruct_onehotd = 4'd8;
        default: q1a8s_destruct_onehotd = 4'd0;
      endcase
    else q1a8s_destruct_onehotd = 4'd0;
  assign _61_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[0]};
  assign _60_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[1]};
  assign lizzieLet11_1_4MQNode_5QNode_Bool_d = {q1a8s_destruct_d[16:1],
                                                q1a8s_destruct_onehotd[2]};
  assign _59_d = {q1a8s_destruct_d[16:1], q1a8s_destruct_onehotd[3]};
  assign q1a8s_destruct_r = (| (q1a8s_destruct_onehotd & {_59_r,
                                                          lizzieLet11_1_4MQNode_5QNode_Bool_r,
                                                          _60_r,
                                                          _61_r}));
  assign lizzieLet11_1_4MQNode_5_r = q1a8s_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet11_1_4MQNode_6,QTree_Bool) (q2a8t_destruct,Pointer_MaskQTree) > [(_58,Pointer_MaskQTree),
                                                                                                          (_57,Pointer_MaskQTree),
                                                                                                          (lizzieLet11_1_4MQNode_6QNode_Bool,Pointer_MaskQTree),
                                                                                                          (_56,Pointer_MaskQTree)] */
  logic [3:0] q2a8t_destruct_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_6_d[0] && q2a8t_destruct_d[0]))
      unique case (lizzieLet11_1_4MQNode_6_d[2:1])
        2'd0: q2a8t_destruct_onehotd = 4'd1;
        2'd1: q2a8t_destruct_onehotd = 4'd2;
        2'd2: q2a8t_destruct_onehotd = 4'd4;
        2'd3: q2a8t_destruct_onehotd = 4'd8;
        default: q2a8t_destruct_onehotd = 4'd0;
      endcase
    else q2a8t_destruct_onehotd = 4'd0;
  assign _58_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[0]};
  assign _57_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[1]};
  assign lizzieLet11_1_4MQNode_6QNode_Bool_d = {q2a8t_destruct_d[16:1],
                                                q2a8t_destruct_onehotd[2]};
  assign _56_d = {q2a8t_destruct_d[16:1], q2a8t_destruct_onehotd[3]};
  assign q2a8t_destruct_r = (| (q2a8t_destruct_onehotd & {_56_r,
                                                          lizzieLet11_1_4MQNode_6QNode_Bool_r,
                                                          _57_r,
                                                          _58_r}));
  assign lizzieLet11_1_4MQNode_6_r = q2a8t_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet11_1_4MQNode_7,QTree_Bool) (q3a8u_destruct,Pointer_MaskQTree) > [(_55,Pointer_MaskQTree),
                                                                                                          (_54,Pointer_MaskQTree),
                                                                                                          (lizzieLet11_1_4MQNode_7QNode_Bool,Pointer_MaskQTree),
                                                                                                          (_53,Pointer_MaskQTree)] */
  logic [3:0] q3a8u_destruct_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_7_d[0] && q3a8u_destruct_d[0]))
      unique case (lizzieLet11_1_4MQNode_7_d[2:1])
        2'd0: q3a8u_destruct_onehotd = 4'd1;
        2'd1: q3a8u_destruct_onehotd = 4'd2;
        2'd2: q3a8u_destruct_onehotd = 4'd4;
        2'd3: q3a8u_destruct_onehotd = 4'd8;
        default: q3a8u_destruct_onehotd = 4'd0;
      endcase
    else q3a8u_destruct_onehotd = 4'd0;
  assign _55_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[0]};
  assign _54_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[1]};
  assign lizzieLet11_1_4MQNode_7QNode_Bool_d = {q3a8u_destruct_d[16:1],
                                                q3a8u_destruct_onehotd[2]};
  assign _53_d = {q3a8u_destruct_d[16:1], q3a8u_destruct_onehotd[3]};
  assign q3a8u_destruct_r = (| (q3a8u_destruct_onehotd & {_53_r,
                                                          lizzieLet11_1_4MQNode_7QNode_Bool_r,
                                                          _54_r,
                                                          _55_r}));
  assign lizzieLet11_1_4MQNode_7_r = q3a8u_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_MaskQTree) : (lizzieLet11_1_4MQNode_8,QTree_Bool) (q4a8v_destruct,Pointer_MaskQTree) > [(_52,Pointer_MaskQTree),
                                                                                                          (_51,Pointer_MaskQTree),
                                                                                                          (lizzieLet11_1_4MQNode_8QNode_Bool,Pointer_MaskQTree),
                                                                                                          (_50,Pointer_MaskQTree)] */
  logic [3:0] q4a8v_destruct_onehotd;
  always_comb
    if ((lizzieLet11_1_4MQNode_8_d[0] && q4a8v_destruct_d[0]))
      unique case (lizzieLet11_1_4MQNode_8_d[2:1])
        2'd0: q4a8v_destruct_onehotd = 4'd1;
        2'd1: q4a8v_destruct_onehotd = 4'd2;
        2'd2: q4a8v_destruct_onehotd = 4'd4;
        2'd3: q4a8v_destruct_onehotd = 4'd8;
        default: q4a8v_destruct_onehotd = 4'd0;
      endcase
    else q4a8v_destruct_onehotd = 4'd0;
  assign _52_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[0]};
  assign _51_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[1]};
  assign lizzieLet11_1_4MQNode_8QNode_Bool_d = {q4a8v_destruct_d[16:1],
                                                q4a8v_destruct_onehotd[2]};
  assign _50_d = {q4a8v_destruct_d[16:1], q4a8v_destruct_onehotd[3]};
  assign q4a8v_destruct_r = (| (q4a8v_destruct_onehotd & {_50_r,
                                                          lizzieLet11_1_4MQNode_8QNode_Bool_r,
                                                          _51_r,
                                                          _52_r}));
  assign lizzieLet11_1_4MQNode_8_r = q4a8v_destruct_r;
  
  /* buf (Ty Pointer_MaskQTree) : (lizzieLet11_1_4MQNode_8QNode_Bool,Pointer_MaskQTree) > (lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d;
  logic lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_r;
  assign lizzieLet11_1_4MQNode_8QNode_Bool_r = ((! lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d[0]) || lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_4MQNode_8QNode_Bool_r)
        lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d <= lizzieLet11_1_4MQNode_8QNode_Bool_d;
  Pointer_MaskQTree_t lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf;
  assign lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_r = (! lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf[0]);
  assign lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_d = (lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf[0] ? lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf :
                                                         lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_r && lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf[0]))
        lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_4MQNode_8QNode_Bool_1_argbuf_r) && (! lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf[0])))
        lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_buf <= lizzieLet11_1_4MQNode_8QNode_Bool_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_QTree_Bool) : (lizzieLet11_1_5,MaskQTree) (ma8q_2,Pointer_QTree_Bool) > [(_49,Pointer_QTree_Bool),
                                                                                           (lizzieLet11_1_5MQVal,Pointer_QTree_Bool),
                                                                                           (_48,Pointer_QTree_Bool)] */
  logic [2:0] ma8q_2_onehotd;
  always_comb
    if ((lizzieLet11_1_5_d[0] && ma8q_2_d[0]))
      unique case (lizzieLet11_1_5_d[2:1])
        2'd0: ma8q_2_onehotd = 3'd1;
        2'd1: ma8q_2_onehotd = 3'd2;
        2'd2: ma8q_2_onehotd = 3'd4;
        default: ma8q_2_onehotd = 3'd0;
      endcase
    else ma8q_2_onehotd = 3'd0;
  assign _49_d = {ma8q_2_d[16:1], ma8q_2_onehotd[0]};
  assign lizzieLet11_1_5MQVal_d = {ma8q_2_d[16:1],
                                   ma8q_2_onehotd[1]};
  assign _48_d = {ma8q_2_d[16:1], ma8q_2_onehotd[2]};
  assign ma8q_2_r = (| (ma8q_2_onehotd & {_48_r,
                                          lizzieLet11_1_5MQVal_r,
                                          _49_r}));
  assign lizzieLet11_1_5_r = ma8q_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet11_1_5MQVal,Pointer_QTree_Bool) > (lizzieLet11_1_5MQVal_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet11_1_5MQVal_bufchan_d;
  logic lizzieLet11_1_5MQVal_bufchan_r;
  assign lizzieLet11_1_5MQVal_r = ((! lizzieLet11_1_5MQVal_bufchan_d[0]) || lizzieLet11_1_5MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_5MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_5MQVal_r)
        lizzieLet11_1_5MQVal_bufchan_d <= lizzieLet11_1_5MQVal_d;
  Pointer_QTree_Bool_t lizzieLet11_1_5MQVal_bufchan_buf;
  assign lizzieLet11_1_5MQVal_bufchan_r = (! lizzieLet11_1_5MQVal_bufchan_buf[0]);
  assign lizzieLet11_1_5MQVal_1_argbuf_d = (lizzieLet11_1_5MQVal_bufchan_buf[0] ? lizzieLet11_1_5MQVal_bufchan_buf :
                                            lizzieLet11_1_5MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_5MQVal_1_argbuf_r && lizzieLet11_1_5MQVal_bufchan_buf[0]))
        lizzieLet11_1_5MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_5MQVal_1_argbuf_r) && (! lizzieLet11_1_5MQVal_bufchan_buf[0])))
        lizzieLet11_1_5MQVal_bufchan_buf <= lizzieLet11_1_5MQVal_bufchan_d;
  
  /* demux (Ty MaskQTree,
       Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_6,MaskQTree) (sc_0_1_goMux_mux,Pointer_CTmain_mask_Bool) > [(lizzieLet11_1_6MQNone,Pointer_CTmain_mask_Bool),
                                                                                                                 (lizzieLet11_1_6MQVal,Pointer_CTmain_mask_Bool),
                                                                                                                 (lizzieLet11_1_6MQNode,Pointer_CTmain_mask_Bool)] */
  logic [2:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet11_1_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet11_1_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 3'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 3'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 3'd4;
        default: sc_0_1_goMux_mux_onehotd = 3'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 3'd0;
  assign lizzieLet11_1_6MQNone_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet11_1_6MQVal_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet11_1_6MQNode_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet11_1_6MQNode_r,
                                                              lizzieLet11_1_6MQVal_r,
                                                              lizzieLet11_1_6MQNone_r}));
  assign lizzieLet11_1_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_6MQNone,Pointer_CTmain_mask_Bool) > (lizzieLet11_1_6MQNone_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQNone_bufchan_d;
  logic lizzieLet11_1_6MQNone_bufchan_r;
  assign lizzieLet11_1_6MQNone_r = ((! lizzieLet11_1_6MQNone_bufchan_d[0]) || lizzieLet11_1_6MQNone_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6MQNone_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_6MQNone_r)
        lizzieLet11_1_6MQNone_bufchan_d <= lizzieLet11_1_6MQNone_d;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQNone_bufchan_buf;
  assign lizzieLet11_1_6MQNone_bufchan_r = (! lizzieLet11_1_6MQNone_bufchan_buf[0]);
  assign lizzieLet11_1_6MQNone_1_argbuf_d = (lizzieLet11_1_6MQNone_bufchan_buf[0] ? lizzieLet11_1_6MQNone_bufchan_buf :
                                             lizzieLet11_1_6MQNone_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_6MQNone_1_argbuf_r && lizzieLet11_1_6MQNone_bufchan_buf[0]))
        lizzieLet11_1_6MQNone_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_6MQNone_1_argbuf_r) && (! lizzieLet11_1_6MQNone_bufchan_buf[0])))
        lizzieLet11_1_6MQNone_bufchan_buf <= lizzieLet11_1_6MQNone_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (lizzieLet11_1_6MQVal,Pointer_CTmain_mask_Bool) > (lizzieLet11_1_6MQVal_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQVal_bufchan_d;
  logic lizzieLet11_1_6MQVal_bufchan_r;
  assign lizzieLet11_1_6MQVal_r = ((! lizzieLet11_1_6MQVal_bufchan_d[0]) || lizzieLet11_1_6MQVal_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6MQVal_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet11_1_6MQVal_r)
        lizzieLet11_1_6MQVal_bufchan_d <= lizzieLet11_1_6MQVal_d;
  Pointer_CTmain_mask_Bool_t lizzieLet11_1_6MQVal_bufchan_buf;
  assign lizzieLet11_1_6MQVal_bufchan_r = (! lizzieLet11_1_6MQVal_bufchan_buf[0]);
  assign lizzieLet11_1_6MQVal_1_argbuf_d = (lizzieLet11_1_6MQVal_bufchan_buf[0] ? lizzieLet11_1_6MQVal_bufchan_buf :
                                            lizzieLet11_1_6MQVal_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet11_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet11_1_6MQVal_1_argbuf_r && lizzieLet11_1_6MQVal_bufchan_buf[0]))
        lizzieLet11_1_6MQVal_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet11_1_6MQVal_1_argbuf_r) && (! lizzieLet11_1_6MQVal_bufchan_buf[0])))
        lizzieLet11_1_6MQVal_bufchan_buf <= lizzieLet11_1_6MQVal_bufchan_d;
  
  /* destruct (Ty CT$wmAdd_Bool,
          Dcon Lcall_$wmAdd_Bool0) : (lizzieLet19_1Lcall_$wmAdd_Bool0,CT$wmAdd_Bool) > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                                                        (es_3_1_destruct,Pointer_QTree_Bool),
                                                                                        (es_4_2_destruct,Pointer_QTree_Bool),
                                                                                        (sc_0_5_destruct,Pointer_CT$wmAdd_Bool)] */
  logic [3:0] lizzieLet19_1Lcall_$wmAdd_Bool0_emitted;
  logic [3:0] lizzieLet19_1Lcall_$wmAdd_Bool0_done;
  assign es_2_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool0_d[19:4],
                              (lizzieLet19_1Lcall_$wmAdd_Bool0_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool0_emitted[0]))};
  assign es_3_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool0_d[35:20],
                              (lizzieLet19_1Lcall_$wmAdd_Bool0_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool0_emitted[1]))};
  assign es_4_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool0_d[51:36],
                              (lizzieLet19_1Lcall_$wmAdd_Bool0_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool0_emitted[2]))};
  assign sc_0_5_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool0_d[67:52],
                              (lizzieLet19_1Lcall_$wmAdd_Bool0_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool0_emitted[3]))};
  assign lizzieLet19_1Lcall_$wmAdd_Bool0_done = (lizzieLet19_1Lcall_$wmAdd_Bool0_emitted | ({sc_0_5_destruct_d[0],
                                                                                             es_4_2_destruct_d[0],
                                                                                             es_3_1_destruct_d[0],
                                                                                             es_2_1_destruct_d[0]} & {sc_0_5_destruct_r,
                                                                                                                      es_4_2_destruct_r,
                                                                                                                      es_3_1_destruct_r,
                                                                                                                      es_2_1_destruct_r}));
  assign lizzieLet19_1Lcall_$wmAdd_Bool0_r = (& lizzieLet19_1Lcall_$wmAdd_Bool0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_1Lcall_$wmAdd_Bool0_emitted <= 4'd0;
    else
      lizzieLet19_1Lcall_$wmAdd_Bool0_emitted <= (lizzieLet19_1Lcall_$wmAdd_Bool0_r ? 4'd0 :
                                                  lizzieLet19_1Lcall_$wmAdd_Bool0_done);
  
  /* destruct (Ty CT$wmAdd_Bool,
          Dcon Lcall_$wmAdd_Bool1) : (lizzieLet19_1Lcall_$wmAdd_Bool1,CT$wmAdd_Bool) > [(es_3_destruct,Pointer_QTree_Bool),
                                                                                        (es_4_1_destruct,Pointer_QTree_Bool),
                                                                                        (sc_0_4_destruct,Pointer_CT$wmAdd_Bool),
                                                                                        (wsib_4_destruct,MyDTBool_Bool_Bool),
                                                                                        (q1a8h_3_destruct,Pointer_QTree_Bool),
                                                                                        (t1a8m_3_destruct,Pointer_QTree_Bool)] */
  logic [5:0] lizzieLet19_1Lcall_$wmAdd_Bool1_emitted;
  logic [5:0] lizzieLet19_1Lcall_$wmAdd_Bool1_done;
  assign es_3_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool1_d[19:4],
                            (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[0]))};
  assign es_4_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool1_d[35:20],
                              (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[1]))};
  assign sc_0_4_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool1_d[51:36],
                              (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[2]))};
  assign wsib_4_destruct_d = (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[3]));
  assign q1a8h_3_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool1_d[67:52],
                               (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[4]))};
  assign t1a8m_3_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool1_d[83:68],
                               (lizzieLet19_1Lcall_$wmAdd_Bool1_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool1_emitted[5]))};
  assign lizzieLet19_1Lcall_$wmAdd_Bool1_done = (lizzieLet19_1Lcall_$wmAdd_Bool1_emitted | ({t1a8m_3_destruct_d[0],
                                                                                             q1a8h_3_destruct_d[0],
                                                                                             wsib_4_destruct_d[0],
                                                                                             sc_0_4_destruct_d[0],
                                                                                             es_4_1_destruct_d[0],
                                                                                             es_3_destruct_d[0]} & {t1a8m_3_destruct_r,
                                                                                                                    q1a8h_3_destruct_r,
                                                                                                                    wsib_4_destruct_r,
                                                                                                                    sc_0_4_destruct_r,
                                                                                                                    es_4_1_destruct_r,
                                                                                                                    es_3_destruct_r}));
  assign lizzieLet19_1Lcall_$wmAdd_Bool1_r = (& lizzieLet19_1Lcall_$wmAdd_Bool1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_1Lcall_$wmAdd_Bool1_emitted <= 6'd0;
    else
      lizzieLet19_1Lcall_$wmAdd_Bool1_emitted <= (lizzieLet19_1Lcall_$wmAdd_Bool1_r ? 6'd0 :
                                                  lizzieLet19_1Lcall_$wmAdd_Bool1_done);
  
  /* destruct (Ty CT$wmAdd_Bool,
          Dcon Lcall_$wmAdd_Bool2) : (lizzieLet19_1Lcall_$wmAdd_Bool2,CT$wmAdd_Bool) > [(es_4_destruct,Pointer_QTree_Bool),
                                                                                        (sc_0_3_destruct,Pointer_CT$wmAdd_Bool),
                                                                                        (wsib_3_destruct,MyDTBool_Bool_Bool),
                                                                                        (q1a8h_2_destruct,Pointer_QTree_Bool),
                                                                                        (t1a8m_2_destruct,Pointer_QTree_Bool),
                                                                                        (q2a8i_2_destruct,Pointer_QTree_Bool),
                                                                                        (t2a8n_2_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet19_1Lcall_$wmAdd_Bool2_emitted;
  logic [6:0] lizzieLet19_1Lcall_$wmAdd_Bool2_done;
  assign es_4_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[19:4],
                            (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[0]))};
  assign sc_0_3_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[35:20],
                              (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[1]))};
  assign wsib_3_destruct_d = (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[2]));
  assign q1a8h_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[51:36],
                               (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[3]))};
  assign t1a8m_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[67:52],
                               (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[4]))};
  assign q2a8i_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[83:68],
                               (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[5]))};
  assign t2a8n_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool2_d[99:84],
                               (lizzieLet19_1Lcall_$wmAdd_Bool2_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool2_emitted[6]))};
  assign lizzieLet19_1Lcall_$wmAdd_Bool2_done = (lizzieLet19_1Lcall_$wmAdd_Bool2_emitted | ({t2a8n_2_destruct_d[0],
                                                                                             q2a8i_2_destruct_d[0],
                                                                                             t1a8m_2_destruct_d[0],
                                                                                             q1a8h_2_destruct_d[0],
                                                                                             wsib_3_destruct_d[0],
                                                                                             sc_0_3_destruct_d[0],
                                                                                             es_4_destruct_d[0]} & {t2a8n_2_destruct_r,
                                                                                                                    q2a8i_2_destruct_r,
                                                                                                                    t1a8m_2_destruct_r,
                                                                                                                    q1a8h_2_destruct_r,
                                                                                                                    wsib_3_destruct_r,
                                                                                                                    sc_0_3_destruct_r,
                                                                                                                    es_4_destruct_r}));
  assign lizzieLet19_1Lcall_$wmAdd_Bool2_r = (& lizzieLet19_1Lcall_$wmAdd_Bool2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_1Lcall_$wmAdd_Bool2_emitted <= 7'd0;
    else
      lizzieLet19_1Lcall_$wmAdd_Bool2_emitted <= (lizzieLet19_1Lcall_$wmAdd_Bool2_r ? 7'd0 :
                                                  lizzieLet19_1Lcall_$wmAdd_Bool2_done);
  
  /* destruct (Ty CT$wmAdd_Bool,
          Dcon Lcall_$wmAdd_Bool3) : (lizzieLet19_1Lcall_$wmAdd_Bool3,CT$wmAdd_Bool) > [(sc_0_2_destruct,Pointer_CT$wmAdd_Bool),
                                                                                        (wsib_2_destruct,MyDTBool_Bool_Bool),
                                                                                        (q1a8h_1_destruct,Pointer_QTree_Bool),
                                                                                        (t1a8m_1_destruct,Pointer_QTree_Bool),
                                                                                        (q2a8i_1_destruct,Pointer_QTree_Bool),
                                                                                        (t2a8n_1_destruct,Pointer_QTree_Bool),
                                                                                        (q3a8j_1_destruct,Pointer_QTree_Bool),
                                                                                        (t3a8o_1_destruct,Pointer_QTree_Bool)] */
  logic [7:0] lizzieLet19_1Lcall_$wmAdd_Bool3_emitted;
  logic [7:0] lizzieLet19_1Lcall_$wmAdd_Bool3_done;
  assign sc_0_2_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[19:4],
                              (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[0]))};
  assign wsib_2_destruct_d = (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[1]));
  assign q1a8h_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[35:20],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[2]))};
  assign t1a8m_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[51:36],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[3]))};
  assign q2a8i_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[67:52],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[4]))};
  assign t2a8n_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[83:68],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[5]))};
  assign q3a8j_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[99:84],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[6]))};
  assign t3a8o_1_destruct_d = {lizzieLet19_1Lcall_$wmAdd_Bool3_d[115:100],
                               (lizzieLet19_1Lcall_$wmAdd_Bool3_d[0] && (! lizzieLet19_1Lcall_$wmAdd_Bool3_emitted[7]))};
  assign lizzieLet19_1Lcall_$wmAdd_Bool3_done = (lizzieLet19_1Lcall_$wmAdd_Bool3_emitted | ({t3a8o_1_destruct_d[0],
                                                                                             q3a8j_1_destruct_d[0],
                                                                                             t2a8n_1_destruct_d[0],
                                                                                             q2a8i_1_destruct_d[0],
                                                                                             t1a8m_1_destruct_d[0],
                                                                                             q1a8h_1_destruct_d[0],
                                                                                             wsib_2_destruct_d[0],
                                                                                             sc_0_2_destruct_d[0]} & {t3a8o_1_destruct_r,
                                                                                                                      q3a8j_1_destruct_r,
                                                                                                                      t2a8n_1_destruct_r,
                                                                                                                      q2a8i_1_destruct_r,
                                                                                                                      t1a8m_1_destruct_r,
                                                                                                                      q1a8h_1_destruct_r,
                                                                                                                      wsib_2_destruct_r,
                                                                                                                      sc_0_2_destruct_r}));
  assign lizzieLet19_1Lcall_$wmAdd_Bool3_r = (& lizzieLet19_1Lcall_$wmAdd_Bool3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_1Lcall_$wmAdd_Bool3_emitted <= 8'd0;
    else
      lizzieLet19_1Lcall_$wmAdd_Bool3_emitted <= (lizzieLet19_1Lcall_$wmAdd_Bool3_r ? 8'd0 :
                                                  lizzieLet19_1Lcall_$wmAdd_Bool3_done);
  
  /* demux (Ty CT$wmAdd_Bool,
       Ty CT$wmAdd_Bool) : (lizzieLet19_2,CT$wmAdd_Bool) (lizzieLet19_1,CT$wmAdd_Bool) > [(_47,CT$wmAdd_Bool),
                                                                                          (lizzieLet19_1Lcall_$wmAdd_Bool3,CT$wmAdd_Bool),
                                                                                          (lizzieLet19_1Lcall_$wmAdd_Bool2,CT$wmAdd_Bool),
                                                                                          (lizzieLet19_1Lcall_$wmAdd_Bool1,CT$wmAdd_Bool),
                                                                                          (lizzieLet19_1Lcall_$wmAdd_Bool0,CT$wmAdd_Bool)] */
  logic [4:0] lizzieLet19_1_onehotd;
  always_comb
    if ((lizzieLet19_2_d[0] && lizzieLet19_1_d[0]))
      unique case (lizzieLet19_2_d[3:1])
        3'd0: lizzieLet19_1_onehotd = 5'd1;
        3'd1: lizzieLet19_1_onehotd = 5'd2;
        3'd2: lizzieLet19_1_onehotd = 5'd4;
        3'd3: lizzieLet19_1_onehotd = 5'd8;
        3'd4: lizzieLet19_1_onehotd = 5'd16;
        default: lizzieLet19_1_onehotd = 5'd0;
      endcase
    else lizzieLet19_1_onehotd = 5'd0;
  assign _47_d = {lizzieLet19_1_d[115:1], lizzieLet19_1_onehotd[0]};
  assign lizzieLet19_1Lcall_$wmAdd_Bool3_d = {lizzieLet19_1_d[115:1],
                                              lizzieLet19_1_onehotd[1]};
  assign lizzieLet19_1Lcall_$wmAdd_Bool2_d = {lizzieLet19_1_d[115:1],
                                              lizzieLet19_1_onehotd[2]};
  assign lizzieLet19_1Lcall_$wmAdd_Bool1_d = {lizzieLet19_1_d[115:1],
                                              lizzieLet19_1_onehotd[3]};
  assign lizzieLet19_1Lcall_$wmAdd_Bool0_d = {lizzieLet19_1_d[115:1],
                                              lizzieLet19_1_onehotd[4]};
  assign lizzieLet19_1_r = (| (lizzieLet19_1_onehotd & {lizzieLet19_1Lcall_$wmAdd_Bool0_r,
                                                        lizzieLet19_1Lcall_$wmAdd_Bool1_r,
                                                        lizzieLet19_1Lcall_$wmAdd_Bool2_r,
                                                        lizzieLet19_1Lcall_$wmAdd_Bool3_r,
                                                        _47_r}));
  assign lizzieLet19_2_r = lizzieLet19_1_r;
  
  /* demux (Ty CT$wmAdd_Bool,
       Ty Go) : (lizzieLet19_3,CT$wmAdd_Bool) (go_7_goMux_data,Go) > [(_46,Go),
                                                                      (lizzieLet19_3Lcall_$wmAdd_Bool3,Go),
                                                                      (lizzieLet19_3Lcall_$wmAdd_Bool2,Go),
                                                                      (lizzieLet19_3Lcall_$wmAdd_Bool1,Go),
                                                                      (lizzieLet19_3Lcall_$wmAdd_Bool0,Go)] */
  logic [4:0] go_7_goMux_data_onehotd;
  always_comb
    if ((lizzieLet19_3_d[0] && go_7_goMux_data_d[0]))
      unique case (lizzieLet19_3_d[3:1])
        3'd0: go_7_goMux_data_onehotd = 5'd1;
        3'd1: go_7_goMux_data_onehotd = 5'd2;
        3'd2: go_7_goMux_data_onehotd = 5'd4;
        3'd3: go_7_goMux_data_onehotd = 5'd8;
        3'd4: go_7_goMux_data_onehotd = 5'd16;
        default: go_7_goMux_data_onehotd = 5'd0;
      endcase
    else go_7_goMux_data_onehotd = 5'd0;
  assign _46_d = go_7_goMux_data_onehotd[0];
  assign lizzieLet19_3Lcall_$wmAdd_Bool3_d = go_7_goMux_data_onehotd[1];
  assign lizzieLet19_3Lcall_$wmAdd_Bool2_d = go_7_goMux_data_onehotd[2];
  assign lizzieLet19_3Lcall_$wmAdd_Bool1_d = go_7_goMux_data_onehotd[3];
  assign lizzieLet19_3Lcall_$wmAdd_Bool0_d = go_7_goMux_data_onehotd[4];
  assign go_7_goMux_data_r = (| (go_7_goMux_data_onehotd & {lizzieLet19_3Lcall_$wmAdd_Bool0_r,
                                                            lizzieLet19_3Lcall_$wmAdd_Bool1_r,
                                                            lizzieLet19_3Lcall_$wmAdd_Bool2_r,
                                                            lizzieLet19_3Lcall_$wmAdd_Bool3_r,
                                                            _46_r}));
  assign lizzieLet19_3_r = go_7_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wmAdd_Bool0,Go) > (lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_r;
  assign lizzieLet19_3Lcall_$wmAdd_Bool0_r = ((! lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d[0]) || lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wmAdd_Bool0_r)
        lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d <= lizzieLet19_3Lcall_$wmAdd_Bool0_d;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf;
  assign lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_r = (! lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_d = (lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf[0] ? lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf :
                                                       lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_r && lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_r) && (! lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_buf <= lizzieLet19_3Lcall_$wmAdd_Bool0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wmAdd_Bool1,Go) > (lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_r;
  assign lizzieLet19_3Lcall_$wmAdd_Bool1_r = ((! lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d[0]) || lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wmAdd_Bool1_r)
        lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d <= lizzieLet19_3Lcall_$wmAdd_Bool1_d;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf;
  assign lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_r = (! lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_d = (lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf[0] ? lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf :
                                                       lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_r && lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wmAdd_Bool1_1_argbuf_r) && (! lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_buf <= lizzieLet19_3Lcall_$wmAdd_Bool1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wmAdd_Bool2,Go) > (lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_r;
  assign lizzieLet19_3Lcall_$wmAdd_Bool2_r = ((! lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d[0]) || lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wmAdd_Bool2_r)
        lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d <= lizzieLet19_3Lcall_$wmAdd_Bool2_d;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf;
  assign lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_r = (! lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_d = (lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf[0] ? lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf :
                                                       lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_r && lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wmAdd_Bool2_1_argbuf_r) && (! lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_buf <= lizzieLet19_3Lcall_$wmAdd_Bool2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wmAdd_Bool3,Go) > (lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d;
  logic lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_r;
  assign lizzieLet19_3Lcall_$wmAdd_Bool3_r = ((! lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d[0]) || lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wmAdd_Bool3_r)
        lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d <= lizzieLet19_3Lcall_$wmAdd_Bool3_d;
  Go_t lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf;
  assign lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_r = (! lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_d = (lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf[0] ? lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf :
                                                       lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_r && lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wmAdd_Bool3_1_argbuf_r) && (! lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_buf <= lizzieLet19_3Lcall_$wmAdd_Bool3_bufchan_d;
  
  /* demux (Ty CT$wmAdd_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet19_4,CT$wmAdd_Bool) (srtarg_0_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet19_4L$wmAdd_Boolsbos,Pointer_QTree_Bool),
                                                                                                         (lizzieLet19_4Lcall_$wmAdd_Bool3,Pointer_QTree_Bool),
                                                                                                         (lizzieLet19_4Lcall_$wmAdd_Bool2,Pointer_QTree_Bool),
                                                                                                         (lizzieLet19_4Lcall_$wmAdd_Bool1,Pointer_QTree_Bool),
                                                                                                         (lizzieLet19_4Lcall_$wmAdd_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet19_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet19_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet19_4L$wmAdd_Boolsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                            srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet19_4Lcall_$wmAdd_Bool3_d = {srtarg_0_goMux_mux_d[16:1],
                                              srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet19_4Lcall_$wmAdd_Bool2_d = {srtarg_0_goMux_mux_d[16:1],
                                              srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet19_4Lcall_$wmAdd_Bool1_d = {srtarg_0_goMux_mux_d[16:1],
                                              srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet19_4Lcall_$wmAdd_Bool0_d = {srtarg_0_goMux_mux_d[16:1],
                                              srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet19_4Lcall_$wmAdd_Bool0_r,
                                                                  lizzieLet19_4Lcall_$wmAdd_Bool1_r,
                                                                  lizzieLet19_4Lcall_$wmAdd_Bool2_r,
                                                                  lizzieLet19_4Lcall_$wmAdd_Bool3_r,
                                                                  lizzieLet19_4L$wmAdd_Boolsbos_r}));
  assign lizzieLet19_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet19_4L$wmAdd_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                     (lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet19_4L$wmAdd_Boolsbos_emitted;
  logic [1:0] lizzieLet19_4L$wmAdd_Boolsbos_done;
  assign lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_d = {lizzieLet19_4L$wmAdd_Boolsbos_d[16:1],
                                                                 (lizzieLet19_4L$wmAdd_Boolsbos_d[0] && (! lizzieLet19_4L$wmAdd_Boolsbos_emitted[0]))};
  assign lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_d = {lizzieLet19_4L$wmAdd_Boolsbos_d[16:1],
                                                                 (lizzieLet19_4L$wmAdd_Boolsbos_d[0] && (! lizzieLet19_4L$wmAdd_Boolsbos_emitted[1]))};
  assign lizzieLet19_4L$wmAdd_Boolsbos_done = (lizzieLet19_4L$wmAdd_Boolsbos_emitted | ({lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_d[0],
                                                                                         lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_r,
                                                                                                                                                     lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet19_4L$wmAdd_Boolsbos_r = (& lizzieLet19_4L$wmAdd_Boolsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_4L$wmAdd_Boolsbos_emitted <= 2'd0;
    else
      lizzieLet19_4L$wmAdd_Boolsbos_emitted <= (lizzieLet19_4L$wmAdd_Boolsbos_r ? 2'd0 :
                                                lizzieLet19_4L$wmAdd_Boolsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_$wmAdd_Bool_goConst,Go) */
  assign call_$wmAdd_Bool_goConst_d = lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_1_r = call_$wmAdd_Bool_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > ($wmAdd_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_r = ((! lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_r)
        lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wmAdd_Bool_resbuf_d  = (lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf :
                                   lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((\$wmAdd_Bool_resbuf_r  && lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! \$wmAdd_Bool_resbuf_r ) && (! lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet19_4L$wmAdd_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet19_4Lcall_$wmAdd_Bool0,Pointer_QTree_Bool),
                          (es_2_1_destruct,Pointer_QTree_Bool),
                          (es_3_1_destruct,Pointer_QTree_Bool),
                          (es_4_2_destruct,Pointer_QTree_Bool)] > (lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool,QTree_Bool) */
  assign lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet19_4Lcall_$wmAdd_Bool0_d[0],
                                                                                                   es_2_1_destruct_d[0],
                                                                                                   es_3_1_destruct_d[0],
                                                                                                   es_4_2_destruct_d[0]}), lizzieLet19_4Lcall_$wmAdd_Bool0_d, es_2_1_destruct_d, es_3_1_destruct_d, es_4_2_destruct_d);
  assign {lizzieLet19_4Lcall_$wmAdd_Bool0_r,
          es_2_1_destruct_r,
          es_3_1_destruct_r,
          es_4_2_destruct_r} = {4 {(lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_r && lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool,QTree_Bool) > (lizzieLet23_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_r;
  assign lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_r = ((! lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d[0]) || lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                        1'd0};
    else
      if (lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_r)
        lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d <= lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_d;
  QTree_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf;
  assign lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_r = (! lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet23_1_argbuf_d = (lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf[0] ? lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf :
                                   lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                          1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf[0]))
        lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                            1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf[0])))
        lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_buf <= lizzieLet19_4Lcall_$wmAdd_Bool0_1es_2_1_1es_3_1_1es_4_2_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Bool,
      Dcon Lcall_$wmAdd_Bool0) : [(lizzieLet19_4Lcall_$wmAdd_Bool1,Pointer_QTree_Bool),
                                  (es_3_destruct,Pointer_QTree_Bool),
                                  (es_4_1_destruct,Pointer_QTree_Bool),
                                  (sc_0_4_destruct,Pointer_CT$wmAdd_Bool)] > (lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0,CT$wmAdd_Bool) */
  assign lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_d = Lcall_$wmAdd_Bool0_dc((& {lizzieLet19_4Lcall_$wmAdd_Bool1_d[0],
                                                                                                                 es_3_destruct_d[0],
                                                                                                                 es_4_1_destruct_d[0],
                                                                                                                 sc_0_4_destruct_d[0]}), lizzieLet19_4Lcall_$wmAdd_Bool1_d, es_3_destruct_d, es_4_1_destruct_d, sc_0_4_destruct_d);
  assign {lizzieLet19_4Lcall_$wmAdd_Bool1_r,
          es_3_destruct_r,
          es_4_1_destruct_r,
          sc_0_4_destruct_r} = {4 {(lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_r && lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_d[0])}};
  
  /* buf (Ty CT$wmAdd_Bool) : (lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0,CT$wmAdd_Bool) > (lizzieLet22_1_argbuf,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_r;
  assign lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_r = ((! lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d[0]) || lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_r)
        lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d <= lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_d;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf;
  assign lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_r = (! lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf[0] ? lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf :
                                   lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf[0]))
        lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf[0])))
        lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_buf <= lizzieLet19_4Lcall_$wmAdd_Bool1_1es_3_1es_4_1_1sc_0_4_1Lcall_$wmAdd_Bool0_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Bool,
      Dcon Lcall_$wmAdd_Bool1) : [(lizzieLet19_4Lcall_$wmAdd_Bool2,Pointer_QTree_Bool),
                                  (es_4_destruct,Pointer_QTree_Bool),
                                  (sc_0_3_destruct,Pointer_CT$wmAdd_Bool),
                                  (wsib_3_1,MyDTBool_Bool_Bool),
                                  (q1a8h_2_destruct,Pointer_QTree_Bool),
                                  (t1a8m_2_destruct,Pointer_QTree_Bool)] > (lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1,CT$wmAdd_Bool) */
  assign lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_d = Lcall_$wmAdd_Bool1_dc((& {lizzieLet19_4Lcall_$wmAdd_Bool2_d[0],
                                                                                                                                   es_4_destruct_d[0],
                                                                                                                                   sc_0_3_destruct_d[0],
                                                                                                                                   wsib_3_1_d[0],
                                                                                                                                   q1a8h_2_destruct_d[0],
                                                                                                                                   t1a8m_2_destruct_d[0]}), lizzieLet19_4Lcall_$wmAdd_Bool2_d, es_4_destruct_d, sc_0_3_destruct_d, wsib_3_1_d, q1a8h_2_destruct_d, t1a8m_2_destruct_d);
  assign {lizzieLet19_4Lcall_$wmAdd_Bool2_r,
          es_4_destruct_r,
          sc_0_3_destruct_r,
          wsib_3_1_r,
          q1a8h_2_destruct_r,
          t1a8m_2_destruct_r} = {6 {(lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_r && lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_d[0])}};
  
  /* buf (Ty CT$wmAdd_Bool) : (lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1,CT$wmAdd_Bool) > (lizzieLet21_1_argbuf,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_r;
  assign lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_r = ((! lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d[0]) || lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d <= {115'd0,
                                                                                                                1'd0};
    else
      if (lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_r)
        lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d <= lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_d;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf;
  assign lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_r = (! lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf[0] ? lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf :
                                   lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf <= {115'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf[0]))
        lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf <= {115'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf[0])))
        lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_buf <= lizzieLet19_4Lcall_$wmAdd_Bool2_1es_4_1sc_0_3_1wsib_3_1q1a8h_2_1t1a8m_2_1Lcall_$wmAdd_Bool1_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Bool,
      Dcon Lcall_$wmAdd_Bool2) : [(lizzieLet19_4Lcall_$wmAdd_Bool3,Pointer_QTree_Bool),
                                  (sc_0_2_destruct,Pointer_CT$wmAdd_Bool),
                                  (wsib_2_1,MyDTBool_Bool_Bool),
                                  (q1a8h_1_destruct,Pointer_QTree_Bool),
                                  (t1a8m_1_destruct,Pointer_QTree_Bool),
                                  (q2a8i_1_destruct,Pointer_QTree_Bool),
                                  (t2a8n_1_destruct,Pointer_QTree_Bool)] > (lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2,CT$wmAdd_Bool) */
  assign lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_d = Lcall_$wmAdd_Bool2_dc((& {lizzieLet19_4Lcall_$wmAdd_Bool3_d[0],
                                                                                                                                               sc_0_2_destruct_d[0],
                                                                                                                                               wsib_2_1_d[0],
                                                                                                                                               q1a8h_1_destruct_d[0],
                                                                                                                                               t1a8m_1_destruct_d[0],
                                                                                                                                               q2a8i_1_destruct_d[0],
                                                                                                                                               t2a8n_1_destruct_d[0]}), lizzieLet19_4Lcall_$wmAdd_Bool3_d, sc_0_2_destruct_d, wsib_2_1_d, q1a8h_1_destruct_d, t1a8m_1_destruct_d, q2a8i_1_destruct_d, t2a8n_1_destruct_d);
  assign {lizzieLet19_4Lcall_$wmAdd_Bool3_r,
          sc_0_2_destruct_r,
          wsib_2_1_r,
          q1a8h_1_destruct_r,
          t1a8m_1_destruct_r,
          q2a8i_1_destruct_r,
          t2a8n_1_destruct_r} = {7 {(lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_r && lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_d[0])}};
  
  /* buf (Ty CT$wmAdd_Bool) : (lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2,CT$wmAdd_Bool) > (lizzieLet20_1_argbuf,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d;
  logic lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_r;
  assign lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_r = ((! lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d[0]) || lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d <= {115'd0,
                                                                                                                            1'd0};
    else
      if (lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_r)
        lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d <= lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_d;
  CT$wmAdd_Bool_t lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf;
  assign lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_r = (! lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf[0] ? lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf :
                                   lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf <= {115'd0,
                                                                                                                              1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf[0]))
        lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf <= {115'd0,
                                                                                                                                1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf[0])))
        lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_buf <= lizzieLet19_4Lcall_$wmAdd_Bool3_1sc_0_2_1wsib_2_1q1a8h_1_1t1a8m_1_1q2a8i_1_1t2a8n_1_1Lcall_$wmAdd_Bool2_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet1_1QNode_Bool,QTree_Bool) > [(q1a8h_destruct,Pointer_QTree_Bool),
                                                                    (q2a8i_destruct,Pointer_QTree_Bool),
                                                                    (q3a8j_destruct,Pointer_QTree_Bool),
                                                                    (q4a8k_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet1_1QNode_Bool_emitted;
  logic [3:0] lizzieLet1_1QNode_Bool_done;
  assign q1a8h_destruct_d = {lizzieLet1_1QNode_Bool_d[18:3],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[0]))};
  assign q2a8i_destruct_d = {lizzieLet1_1QNode_Bool_d[34:19],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[1]))};
  assign q3a8j_destruct_d = {lizzieLet1_1QNode_Bool_d[50:35],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[2]))};
  assign q4a8k_destruct_d = {lizzieLet1_1QNode_Bool_d[66:51],
                             (lizzieLet1_1QNode_Bool_d[0] && (! lizzieLet1_1QNode_Bool_emitted[3]))};
  assign lizzieLet1_1QNode_Bool_done = (lizzieLet1_1QNode_Bool_emitted | ({q4a8k_destruct_d[0],
                                                                           q3a8j_destruct_d[0],
                                                                           q2a8i_destruct_d[0],
                                                                           q1a8h_destruct_d[0]} & {q4a8k_destruct_r,
                                                                                                   q3a8j_destruct_r,
                                                                                                   q2a8i_destruct_r,
                                                                                                   q1a8h_destruct_r}));
  assign lizzieLet1_1QNode_Bool_r = (& lizzieLet1_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet1_1QNode_Bool_emitted <= (lizzieLet1_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet1_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet1_1QVal_Bool,QTree_Bool) > [(v1a8b_destruct,MyBool)] */
  assign v1a8b_destruct_d = {lizzieLet1_1QVal_Bool_d[3:3],
                             lizzieLet1_1QVal_Bool_d[0]};
  assign lizzieLet1_1QVal_Bool_r = v1a8b_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet1_2,QTree_Bool) (lizzieLet1_1,QTree_Bool) > [(_45,QTree_Bool),
                                                                               (lizzieLet1_1QVal_Bool,QTree_Bool),
                                                                               (lizzieLet1_1QNode_Bool,QTree_Bool),
                                                                               (_44,QTree_Bool)] */
  logic [3:0] lizzieLet1_1_onehotd;
  always_comb
    if ((lizzieLet1_2_d[0] && lizzieLet1_1_d[0]))
      unique case (lizzieLet1_2_d[2:1])
        2'd0: lizzieLet1_1_onehotd = 4'd1;
        2'd1: lizzieLet1_1_onehotd = 4'd2;
        2'd2: lizzieLet1_1_onehotd = 4'd4;
        2'd3: lizzieLet1_1_onehotd = 4'd8;
        default: lizzieLet1_1_onehotd = 4'd0;
      endcase
    else lizzieLet1_1_onehotd = 4'd0;
  assign _45_d = {lizzieLet1_1_d[66:1], lizzieLet1_1_onehotd[0]};
  assign lizzieLet1_1QVal_Bool_d = {lizzieLet1_1_d[66:1],
                                    lizzieLet1_1_onehotd[1]};
  assign lizzieLet1_1QNode_Bool_d = {lizzieLet1_1_d[66:1],
                                     lizzieLet1_1_onehotd[2]};
  assign _44_d = {lizzieLet1_1_d[66:1], lizzieLet1_1_onehotd[3]};
  assign lizzieLet1_1_r = (| (lizzieLet1_1_onehotd & {_44_r,
                                                      lizzieLet1_1QNode_Bool_r,
                                                      lizzieLet1_1QVal_Bool_r,
                                                      _45_r}));
  assign lizzieLet1_2_r = lizzieLet1_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet1_3,QTree_Bool) (go_4_goMux_data,Go) > [(lizzieLet1_3QNone_Bool,Go),
                                                                  (lizzieLet1_3QVal_Bool,Go),
                                                                  (lizzieLet1_3QNode_Bool,Go),
                                                                  (lizzieLet1_3QError_Bool,Go)] */
  logic [3:0] go_4_goMux_data_onehotd;
  always_comb
    if ((lizzieLet1_3_d[0] && go_4_goMux_data_d[0]))
      unique case (lizzieLet1_3_d[2:1])
        2'd0: go_4_goMux_data_onehotd = 4'd1;
        2'd1: go_4_goMux_data_onehotd = 4'd2;
        2'd2: go_4_goMux_data_onehotd = 4'd4;
        2'd3: go_4_goMux_data_onehotd = 4'd8;
        default: go_4_goMux_data_onehotd = 4'd0;
      endcase
    else go_4_goMux_data_onehotd = 4'd0;
  assign lizzieLet1_3QNone_Bool_d = go_4_goMux_data_onehotd[0];
  assign lizzieLet1_3QVal_Bool_d = go_4_goMux_data_onehotd[1];
  assign lizzieLet1_3QNode_Bool_d = go_4_goMux_data_onehotd[2];
  assign lizzieLet1_3QError_Bool_d = go_4_goMux_data_onehotd[3];
  assign go_4_goMux_data_r = (| (go_4_goMux_data_onehotd & {lizzieLet1_3QError_Bool_r,
                                                            lizzieLet1_3QNode_Bool_r,
                                                            lizzieLet1_3QVal_Bool_r,
                                                            lizzieLet1_3QNone_Bool_r}));
  assign lizzieLet1_3_r = go_4_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet1_3QError_Bool,Go) > [(lizzieLet1_3QError_Bool_1,Go),
                                               (lizzieLet1_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet1_3QError_Bool_emitted;
  logic [1:0] lizzieLet1_3QError_Bool_done;
  assign lizzieLet1_3QError_Bool_1_d = (lizzieLet1_3QError_Bool_d[0] && (! lizzieLet1_3QError_Bool_emitted[0]));
  assign lizzieLet1_3QError_Bool_2_d = (lizzieLet1_3QError_Bool_d[0] && (! lizzieLet1_3QError_Bool_emitted[1]));
  assign lizzieLet1_3QError_Bool_done = (lizzieLet1_3QError_Bool_emitted | ({lizzieLet1_3QError_Bool_2_d[0],
                                                                             lizzieLet1_3QError_Bool_1_d[0]} & {lizzieLet1_3QError_Bool_2_r,
                                                                                                                lizzieLet1_3QError_Bool_1_r}));
  assign lizzieLet1_3QError_Bool_r = (& lizzieLet1_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet1_3QError_Bool_emitted <= (lizzieLet1_3QError_Bool_r ? 2'd0 :
                                          lizzieLet1_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet1_3QError_Bool_1,Go)] > (lizzieLet1_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet1_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet1_3QError_Bool_1_d[0]}), lizzieLet1_3QError_Bool_1_d);
  assign {lizzieLet1_3QError_Bool_1_r} = {1 {(lizzieLet1_3QError_Bool_1QError_Bool_r && lizzieLet1_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet1_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet10_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet1_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet1_3QError_Bool_1QError_Bool_r = ((! lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet1_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet1_3QError_Bool_1QError_Bool_r)
        lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet1_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet1_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf :
                                     lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet1_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet1_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QError_Bool_2,Go) > (lizzieLet1_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_3QError_Bool_2_bufchan_d;
  logic lizzieLet1_3QError_Bool_2_bufchan_r;
  assign lizzieLet1_3QError_Bool_2_r = ((! lizzieLet1_3QError_Bool_2_bufchan_d[0]) || lizzieLet1_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QError_Bool_2_r)
        lizzieLet1_3QError_Bool_2_bufchan_d <= lizzieLet1_3QError_Bool_2_d;
  Go_t lizzieLet1_3QError_Bool_2_bufchan_buf;
  assign lizzieLet1_3QError_Bool_2_bufchan_r = (! lizzieLet1_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_3QError_Bool_2_argbuf_d = (lizzieLet1_3QError_Bool_2_bufchan_buf[0] ? lizzieLet1_3QError_Bool_2_bufchan_buf :
                                               lizzieLet1_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QError_Bool_2_argbuf_r && lizzieLet1_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet1_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QError_Bool_2_argbuf_r) && (! lizzieLet1_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet1_3QError_Bool_2_bufchan_buf <= lizzieLet1_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_3QNone_Bool,Go) > (lizzieLet1_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_3QNone_Bool_bufchan_d;
  logic lizzieLet1_3QNone_Bool_bufchan_r;
  assign lizzieLet1_3QNone_Bool_r = ((! lizzieLet1_3QNone_Bool_bufchan_d[0]) || lizzieLet1_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_3QNone_Bool_r)
        lizzieLet1_3QNone_Bool_bufchan_d <= lizzieLet1_3QNone_Bool_d;
  Go_t lizzieLet1_3QNone_Bool_bufchan_buf;
  assign lizzieLet1_3QNone_Bool_bufchan_r = (! lizzieLet1_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_3QNone_Bool_1_argbuf_d = (lizzieLet1_3QNone_Bool_bufchan_buf[0] ? lizzieLet1_3QNone_Bool_bufchan_buf :
                                              lizzieLet1_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_3QNone_Bool_1_argbuf_r && lizzieLet1_3QNone_Bool_bufchan_buf[0]))
        lizzieLet1_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_3QNone_Bool_1_argbuf_r) && (! lizzieLet1_3QNone_Bool_bufchan_buf[0])))
        lizzieLet1_3QNone_Bool_bufchan_buf <= lizzieLet1_3QNone_Bool_bufchan_d;
  
  /* mergectrl (Ty C10,Ty Go) : [(lizzieLet1_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf,Go),
                            (lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf,Go),
                            (lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf,Go),
                            (lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf,Go),
                            (lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf,Go),
                            (lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf,Go),
                            (lizzieLet1_3QError_Bool_2_argbuf,Go)] > (go_7_goMux_choice,C10) (go_7_goMux_data,Go) */
  logic [9:0] lizzieLet1_3QNone_Bool_1_argbuf_select_d;
  assign lizzieLet1_3QNone_Bool_1_argbuf_select_d = ((| lizzieLet1_3QNone_Bool_1_argbuf_select_q) ? lizzieLet1_3QNone_Bool_1_argbuf_select_q :
                                                     (lizzieLet1_3QNone_Bool_1_argbuf_d[0] ? 10'd1 :
                                                      (lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_d[0] ? 10'd2 :
                                                       (lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_d[0] ? 10'd4 :
                                                        (lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_d[0] ? 10'd8 :
                                                         (lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_d[0] ? 10'd16 :
                                                          (lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_d[0] ? 10'd32 :
                                                           (lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_d[0] ? 10'd64 :
                                                            (lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_d[0] ? 10'd128 :
                                                             (lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_d[0] ? 10'd256 :
                                                              (lizzieLet1_3QError_Bool_2_argbuf_d[0] ? 10'd512 :
                                                               10'd0)))))))))));
  logic [9:0] lizzieLet1_3QNone_Bool_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_1_argbuf_select_q <= 10'd0;
    else
      lizzieLet1_3QNone_Bool_1_argbuf_select_q <= (lizzieLet1_3QNone_Bool_1_argbuf_done ? 10'd0 :
                                                   lizzieLet1_3QNone_Bool_1_argbuf_select_d);
  logic [1:0] lizzieLet1_3QNone_Bool_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_3QNone_Bool_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet1_3QNone_Bool_1_argbuf_emit_q <= (lizzieLet1_3QNone_Bool_1_argbuf_done ? 2'd0 :
                                                 lizzieLet1_3QNone_Bool_1_argbuf_emit_d);
  logic [1:0] lizzieLet1_3QNone_Bool_1_argbuf_emit_d;
  assign lizzieLet1_3QNone_Bool_1_argbuf_emit_d = (lizzieLet1_3QNone_Bool_1_argbuf_emit_q | ({go_7_goMux_choice_d[0],
                                                                                              go_7_goMux_data_d[0]} & {go_7_goMux_choice_r,
                                                                                                                       go_7_goMux_data_r}));
  logic lizzieLet1_3QNone_Bool_1_argbuf_done;
  assign lizzieLet1_3QNone_Bool_1_argbuf_done = (& lizzieLet1_3QNone_Bool_1_argbuf_emit_d);
  assign {lizzieLet1_3QError_Bool_2_argbuf_r,
          lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_r,
          lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_r,
          lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_r,
          lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_r,
          lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_r,
          lizzieLet1_3QNone_Bool_1_argbuf_r} = (lizzieLet1_3QNone_Bool_1_argbuf_done ? lizzieLet1_3QNone_Bool_1_argbuf_select_d :
                                                10'd0);
  assign go_7_goMux_data_d = ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_3QNone_Bool_1_argbuf_d :
                              ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet19_3Lcall_$wmAdd_Bool0_1_argbuf_d :
                               ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_d :
                                ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_d :
                                 ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_d :
                                  ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_d :
                                   ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_d :
                                    ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_d :
                                     ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_d :
                                      ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[0])) ? lizzieLet1_3QError_Bool_2_argbuf_d :
                                       1'd0))))))))));
  assign go_7_goMux_choice_d = ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[0] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C1_10_dc(1'd1) :
                                ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[1] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C2_10_dc(1'd1) :
                                 ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[2] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C3_10_dc(1'd1) :
                                  ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[3] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C4_10_dc(1'd1) :
                                   ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[4] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C5_10_dc(1'd1) :
                                    ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[5] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C6_10_dc(1'd1) :
                                     ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[6] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C7_10_dc(1'd1) :
                                      ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[7] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C8_10_dc(1'd1) :
                                       ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[8] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C9_10_dc(1'd1) :
                                        ((lizzieLet1_3QNone_Bool_1_argbuf_select_d[9] && (! lizzieLet1_3QNone_Bool_1_argbuf_emit_q[1])) ? C10_10_dc(1'd1) :
                                         {4'd0, 1'd0}))))))))));
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet1_4,QTree_Bool) (readPointer_QTree_Boolw2sid_1_1_argbuf_rwb,QTree_Bool) > [(_43,QTree_Bool),
                                                                                                             (lizzieLet1_4QVal_Bool,QTree_Bool),
                                                                                                             (lizzieLet1_4QNode_Bool,QTree_Bool),
                                                                                                             (_42,QTree_Bool)] */
  logic [3:0] readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet1_4_d[0] && readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d[0]))
      unique case (lizzieLet1_4_d[2:1])
        2'd0: readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd1;
        2'd1: readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd2;
        2'd2: readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd4;
        2'd3: readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd8;
        default: readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd0;
      endcase
    else readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd = 4'd0;
  assign _43_d = {readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet1_4QVal_Bool_d = {readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d[66:1],
                                    readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_d = {readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d[66:1],
                                     readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd[2]};
  assign _42_d = {readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d[66:1],
                  readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd[3]};
  assign readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_r = (| (readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_onehotd & {_42_r,
                                                                                                                  lizzieLet1_4QNode_Bool_r,
                                                                                                                  lizzieLet1_4QVal_Bool_r,
                                                                                                                  _43_r}));
  assign lizzieLet1_4_r = readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet1_4QNode_Bool,QTree_Bool) > [(lizzieLet1_4QNode_Bool_1,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_2,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_3,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_4,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_5,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_6,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_7,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_8,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_9,QTree_Bool),
                                                              (lizzieLet1_4QNode_Bool_10,QTree_Bool)] */
  logic [9:0] lizzieLet1_4QNode_Bool_emitted;
  logic [9:0] lizzieLet1_4QNode_Bool_done;
  assign lizzieLet1_4QNode_Bool_1_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[0]))};
  assign lizzieLet1_4QNode_Bool_2_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[1]))};
  assign lizzieLet1_4QNode_Bool_3_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[2]))};
  assign lizzieLet1_4QNode_Bool_4_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[3]))};
  assign lizzieLet1_4QNode_Bool_5_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[4]))};
  assign lizzieLet1_4QNode_Bool_6_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[5]))};
  assign lizzieLet1_4QNode_Bool_7_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[6]))};
  assign lizzieLet1_4QNode_Bool_8_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[7]))};
  assign lizzieLet1_4QNode_Bool_9_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                       (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[8]))};
  assign lizzieLet1_4QNode_Bool_10_d = {lizzieLet1_4QNode_Bool_d[66:1],
                                        (lizzieLet1_4QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_emitted[9]))};
  assign lizzieLet1_4QNode_Bool_done = (lizzieLet1_4QNode_Bool_emitted | ({lizzieLet1_4QNode_Bool_10_d[0],
                                                                           lizzieLet1_4QNode_Bool_9_d[0],
                                                                           lizzieLet1_4QNode_Bool_8_d[0],
                                                                           lizzieLet1_4QNode_Bool_7_d[0],
                                                                           lizzieLet1_4QNode_Bool_6_d[0],
                                                                           lizzieLet1_4QNode_Bool_5_d[0],
                                                                           lizzieLet1_4QNode_Bool_4_d[0],
                                                                           lizzieLet1_4QNode_Bool_3_d[0],
                                                                           lizzieLet1_4QNode_Bool_2_d[0],
                                                                           lizzieLet1_4QNode_Bool_1_d[0]} & {lizzieLet1_4QNode_Bool_10_r,
                                                                                                             lizzieLet1_4QNode_Bool_9_r,
                                                                                                             lizzieLet1_4QNode_Bool_8_r,
                                                                                                             lizzieLet1_4QNode_Bool_7_r,
                                                                                                             lizzieLet1_4QNode_Bool_6_r,
                                                                                                             lizzieLet1_4QNode_Bool_5_r,
                                                                                                             lizzieLet1_4QNode_Bool_4_r,
                                                                                                             lizzieLet1_4QNode_Bool_3_r,
                                                                                                             lizzieLet1_4QNode_Bool_2_r,
                                                                                                             lizzieLet1_4QNode_Bool_1_r}));
  assign lizzieLet1_4QNode_Bool_r = (& lizzieLet1_4QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_4QNode_Bool_emitted <= 10'd0;
    else
      lizzieLet1_4QNode_Bool_emitted <= (lizzieLet1_4QNode_Bool_r ? 10'd0 :
                                         lizzieLet1_4QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_10,QTree_Bool) (q4a8k_destruct,Pointer_QTree_Bool) > [(_41,Pointer_QTree_Bool),
                                                                                                              (_40,Pointer_QTree_Bool),
                                                                                                              (lizzieLet1_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool),
                                                                                                              (_39,Pointer_QTree_Bool)] */
  logic [3:0] q4a8k_destruct_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_10_d[0] && q4a8k_destruct_d[0]))
      unique case (lizzieLet1_4QNode_Bool_10_d[2:1])
        2'd0: q4a8k_destruct_onehotd = 4'd1;
        2'd1: q4a8k_destruct_onehotd = 4'd2;
        2'd2: q4a8k_destruct_onehotd = 4'd4;
        2'd3: q4a8k_destruct_onehotd = 4'd8;
        default: q4a8k_destruct_onehotd = 4'd0;
      endcase
    else q4a8k_destruct_onehotd = 4'd0;
  assign _41_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[0]};
  assign _40_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_10QNode_Bool_d = {q4a8k_destruct_d[16:1],
                                                  q4a8k_destruct_onehotd[2]};
  assign _39_d = {q4a8k_destruct_d[16:1], q4a8k_destruct_onehotd[3]};
  assign q4a8k_destruct_r = (| (q4a8k_destruct_onehotd & {_39_r,
                                                          lizzieLet1_4QNode_Bool_10QNode_Bool_r,
                                                          _40_r,
                                                          _41_r}));
  assign lizzieLet1_4QNode_Bool_10_r = q4a8k_destruct_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_10QNode_Bool,Pointer_QTree_Bool) > (lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_10QNode_Bool_r = ((! lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNode_Bool_10QNode_Bool_r)
        lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_10QNode_Bool_d;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf :
                                                           lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNode_Bool_10QNode_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_10QNode_Bool_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet1_4QNode_Bool_1QNode_Bool,QTree_Bool) > [(t1a8m_destruct,Pointer_QTree_Bool),
                                                                                (t2a8n_destruct,Pointer_QTree_Bool),
                                                                                (t3a8o_destruct,Pointer_QTree_Bool),
                                                                                (t4a8p_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet1_4QNode_Bool_1QNode_Bool_emitted;
  logic [3:0] lizzieLet1_4QNode_Bool_1QNode_Bool_done;
  assign t1a8m_destruct_d = {lizzieLet1_4QNode_Bool_1QNode_Bool_d[18:3],
                             (lizzieLet1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_1QNode_Bool_emitted[0]))};
  assign t2a8n_destruct_d = {lizzieLet1_4QNode_Bool_1QNode_Bool_d[34:19],
                             (lizzieLet1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_1QNode_Bool_emitted[1]))};
  assign t3a8o_destruct_d = {lizzieLet1_4QNode_Bool_1QNode_Bool_d[50:35],
                             (lizzieLet1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_1QNode_Bool_emitted[2]))};
  assign t4a8p_destruct_d = {lizzieLet1_4QNode_Bool_1QNode_Bool_d[66:51],
                             (lizzieLet1_4QNode_Bool_1QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_1QNode_Bool_emitted[3]))};
  assign lizzieLet1_4QNode_Bool_1QNode_Bool_done = (lizzieLet1_4QNode_Bool_1QNode_Bool_emitted | ({t4a8p_destruct_d[0],
                                                                                                   t3a8o_destruct_d[0],
                                                                                                   t2a8n_destruct_d[0],
                                                                                                   t1a8m_destruct_d[0]} & {t4a8p_destruct_r,
                                                                                                                           t3a8o_destruct_r,
                                                                                                                           t2a8n_destruct_r,
                                                                                                                           t1a8m_destruct_r}));
  assign lizzieLet1_4QNode_Bool_1QNode_Bool_r = (& lizzieLet1_4QNode_Bool_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet1_4QNode_Bool_1QNode_Bool_emitted <= (lizzieLet1_4QNode_Bool_1QNode_Bool_r ? 4'd0 :
                                                     lizzieLet1_4QNode_Bool_1QNode_Bool_done);
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet1_4QNode_Bool_2,QTree_Bool) (lizzieLet1_4QNode_Bool_1,QTree_Bool) > [(_38,QTree_Bool),
                                                                                                       (_37,QTree_Bool),
                                                                                                       (lizzieLet1_4QNode_Bool_1QNode_Bool,QTree_Bool),
                                                                                                       (_36,QTree_Bool)] */
  logic [3:0] lizzieLet1_4QNode_Bool_1_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_2_d[0] && lizzieLet1_4QNode_Bool_1_d[0]))
      unique case (lizzieLet1_4QNode_Bool_2_d[2:1])
        2'd0: lizzieLet1_4QNode_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet1_4QNode_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet1_4QNode_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet1_4QNode_Bool_1_onehotd = 4'd8;
        default: lizzieLet1_4QNode_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet1_4QNode_Bool_1_onehotd = 4'd0;
  assign _38_d = {lizzieLet1_4QNode_Bool_1_d[66:1],
                  lizzieLet1_4QNode_Bool_1_onehotd[0]};
  assign _37_d = {lizzieLet1_4QNode_Bool_1_d[66:1],
                  lizzieLet1_4QNode_Bool_1_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_1QNode_Bool_d = {lizzieLet1_4QNode_Bool_1_d[66:1],
                                                 lizzieLet1_4QNode_Bool_1_onehotd[2]};
  assign _36_d = {lizzieLet1_4QNode_Bool_1_d[66:1],
                  lizzieLet1_4QNode_Bool_1_onehotd[3]};
  assign lizzieLet1_4QNode_Bool_1_r = (| (lizzieLet1_4QNode_Bool_1_onehotd & {_36_r,
                                                                              lizzieLet1_4QNode_Bool_1QNode_Bool_r,
                                                                              _37_r,
                                                                              _38_r}));
  assign lizzieLet1_4QNode_Bool_2_r = lizzieLet1_4QNode_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet1_4QNode_Bool_3,QTree_Bool) (lizzieLet1_3QNode_Bool,Go) > [(lizzieLet1_4QNode_Bool_3QNone_Bool,Go),
                                                                                     (lizzieLet1_4QNode_Bool_3QVal_Bool,Go),
                                                                                     (lizzieLet1_4QNode_Bool_3QNode_Bool,Go),
                                                                                     (lizzieLet1_4QNode_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet1_3QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_3_d[0] && lizzieLet1_3QNode_Bool_d[0]))
      unique case (lizzieLet1_4QNode_Bool_3_d[2:1])
        2'd0: lizzieLet1_3QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_3QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_3QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_3QNode_Bool_onehotd = 4'd8;
        default: lizzieLet1_3QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_3QNode_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QNode_Bool_3QNone_Bool_d = lizzieLet1_3QNode_Bool_onehotd[0];
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_d = lizzieLet1_3QNode_Bool_onehotd[1];
  assign lizzieLet1_4QNode_Bool_3QNode_Bool_d = lizzieLet1_3QNode_Bool_onehotd[2];
  assign lizzieLet1_4QNode_Bool_3QError_Bool_d = lizzieLet1_3QNode_Bool_onehotd[3];
  assign lizzieLet1_3QNode_Bool_r = (| (lizzieLet1_3QNode_Bool_onehotd & {lizzieLet1_4QNode_Bool_3QError_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_3QNode_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_3QVal_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_3QNone_Bool_r}));
  assign lizzieLet1_4QNode_Bool_3_r = lizzieLet1_3QNode_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet1_4QNode_Bool_3QError_Bool,Go) > [(lizzieLet1_4QNode_Bool_3QError_Bool_1,Go),
                                                           (lizzieLet1_4QNode_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet1_4QNode_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet1_4QNode_Bool_3QError_Bool_done;
  assign lizzieLet1_4QNode_Bool_3QError_Bool_1_d = (lizzieLet1_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet1_4QNode_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet1_4QNode_Bool_3QError_Bool_2_d = (lizzieLet1_4QNode_Bool_3QError_Bool_d[0] && (! lizzieLet1_4QNode_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet1_4QNode_Bool_3QError_Bool_done = (lizzieLet1_4QNode_Bool_3QError_Bool_emitted | ({lizzieLet1_4QNode_Bool_3QError_Bool_2_d[0],
                                                                                                     lizzieLet1_4QNode_Bool_3QError_Bool_1_d[0]} & {lizzieLet1_4QNode_Bool_3QError_Bool_2_r,
                                                                                                                                                    lizzieLet1_4QNode_Bool_3QError_Bool_1_r}));
  assign lizzieLet1_4QNode_Bool_3QError_Bool_r = (& lizzieLet1_4QNode_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QNode_Bool_3QError_Bool_emitted <= (lizzieLet1_4QNode_Bool_3QError_Bool_r ? 2'd0 :
                                                      lizzieLet1_4QNode_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet1_4QNode_Bool_3QError_Bool_1,Go)] > (lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet1_4QNode_Bool_3QError_Bool_1_d[0]}), lizzieLet1_4QNode_Bool_3QError_Bool_1_d);
  assign {lizzieLet1_4QNode_Bool_3QError_Bool_1_r} = {1 {(lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_r && lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet9_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                     1'd0};
    else
      if (lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                    lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                         1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QNode_Bool_3QError_Bool_2,Go) > (lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QError_Bool_2_r = ((! lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QNode_Bool_3QError_Bool_2_r)
        lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d <= lizzieLet1_4QNode_Bool_3QError_Bool_2_d;
  Go_t lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_d = (lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf :
                                                           lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_r && lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QNode_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet1_4QNode_Bool_3QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QNode_Bool_3QNode_Bool,Go) > (lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QNode_Bool_r = ((! lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QNode_Bool_3QNode_Bool_r)
        lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_3QNode_Bool_d;
  Go_t lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf :
                                                          lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QNode_Bool_3QNode_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_3QNode_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QNode_Bool_3QNone_Bool,Go) > (lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QNone_Bool_r = ((! lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QNode_Bool_3QNone_Bool_r)
        lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_3QNone_Bool_d;
  Go_t lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf :
                                                          lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QNode_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_3QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet1_4QNode_Bool_3QVal_Bool,Go) > [(lizzieLet1_4QNode_Bool_3QVal_Bool_1,Go),
                                                         (lizzieLet1_4QNode_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet1_4QNode_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet1_4QNode_Bool_3QVal_Bool_done;
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_1_d = (lizzieLet1_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet1_4QNode_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_2_d = (lizzieLet1_4QNode_Bool_3QVal_Bool_d[0] && (! lizzieLet1_4QNode_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_done = (lizzieLet1_4QNode_Bool_3QVal_Bool_emitted | ({lizzieLet1_4QNode_Bool_3QVal_Bool_2_d[0],
                                                                                                 lizzieLet1_4QNode_Bool_3QVal_Bool_1_d[0]} & {lizzieLet1_4QNode_Bool_3QVal_Bool_2_r,
                                                                                                                                              lizzieLet1_4QNode_Bool_3QVal_Bool_1_r}));
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_r = (& lizzieLet1_4QNode_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QNode_Bool_3QVal_Bool_emitted <= (lizzieLet1_4QNode_Bool_3QVal_Bool_r ? 2'd0 :
                                                    lizzieLet1_4QNode_Bool_3QVal_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet1_4QNode_Bool_3QVal_Bool_1,Go)] > (lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet1_4QNode_Bool_3QVal_Bool_1_d[0]}), lizzieLet1_4QNode_Bool_3QVal_Bool_1_d);
  assign {lizzieLet1_4QNode_Bool_3QVal_Bool_1_r} = {1 {(lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_r && lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool,QTree_Bool) > (lizzieLet7_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_r = ((! lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_r)
        lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf :
                                    lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_3QVal_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QNode_Bool_3QVal_Bool_2,Go) > (lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_2_r = ((! lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QNode_Bool_3QVal_Bool_2_r)
        lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet1_4QNode_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf :
                                                         lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_r && lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QNode_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet1_4QNode_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QNode_Bool_4,QTree_Bool) (lizzieLet1_5QNode_Bool,Pointer_CT$wmAdd_Bool) > [(lizzieLet1_4QNode_Bool_4QNone_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                           (lizzieLet1_4QNode_Bool_4QVal_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                           (lizzieLet1_4QNode_Bool_4QNode_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                           (lizzieLet1_4QNode_Bool_4QError_Bool,Pointer_CT$wmAdd_Bool)] */
  logic [3:0] lizzieLet1_5QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_4_d[0] && lizzieLet1_5QNode_Bool_d[0]))
      unique case (lizzieLet1_4QNode_Bool_4_d[2:1])
        2'd0: lizzieLet1_5QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_5QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_5QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_5QNode_Bool_onehotd = 4'd8;
        default: lizzieLet1_5QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_5QNode_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QNode_Bool_4QNone_Bool_d = {lizzieLet1_5QNode_Bool_d[16:1],
                                                 lizzieLet1_5QNode_Bool_onehotd[0]};
  assign lizzieLet1_4QNode_Bool_4QVal_Bool_d = {lizzieLet1_5QNode_Bool_d[16:1],
                                                lizzieLet1_5QNode_Bool_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_4QNode_Bool_d = {lizzieLet1_5QNode_Bool_d[16:1],
                                                 lizzieLet1_5QNode_Bool_onehotd[2]};
  assign lizzieLet1_4QNode_Bool_4QError_Bool_d = {lizzieLet1_5QNode_Bool_d[16:1],
                                                  lizzieLet1_5QNode_Bool_onehotd[3]};
  assign lizzieLet1_5QNode_Bool_r = (| (lizzieLet1_5QNode_Bool_onehotd & {lizzieLet1_4QNode_Bool_4QError_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_4QNode_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_4QVal_Bool_r,
                                                                          lizzieLet1_4QNode_Bool_4QNone_Bool_r}));
  assign lizzieLet1_4QNode_Bool_4_r = lizzieLet1_5QNode_Bool_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QNode_Bool_4QError_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_4QError_Bool_r = ((! lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNode_Bool_4QError_Bool_r)
        lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_4QError_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf :
                                                           lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNode_Bool_4QError_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_4QError_Bool_bufchan_d;
  
  /* dcon (Ty CT$wmAdd_Bool,
      Dcon Lcall_$wmAdd_Bool3) : [(lizzieLet1_4QNode_Bool_4QNode_Bool,Pointer_CT$wmAdd_Bool),
                                  (lizzieLet1_4QNode_Bool_6QNode_Bool_1,MyDTBool_Bool_Bool),
                                  (lizzieLet1_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                  (t1a8m_destruct,Pointer_QTree_Bool),
                                  (lizzieLet1_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                  (t2a8n_destruct,Pointer_QTree_Bool),
                                  (lizzieLet1_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                  (t3a8o_destruct,Pointer_QTree_Bool)] > (lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3,CT$wmAdd_Bool) */
  assign lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_d = Lcall_$wmAdd_Bool3_dc((& {lizzieLet1_4QNode_Bool_4QNode_Bool_d[0],
                                                                                                                                                                                                                                                                   lizzieLet1_4QNode_Bool_6QNode_Bool_1_d[0],
                                                                                                                                                                                                                                                                   lizzieLet1_4QNode_Bool_7QNode_Bool_d[0],
                                                                                                                                                                                                                                                                   t1a8m_destruct_d[0],
                                                                                                                                                                                                                                                                   lizzieLet1_4QNode_Bool_8QNode_Bool_d[0],
                                                                                                                                                                                                                                                                   t2a8n_destruct_d[0],
                                                                                                                                                                                                                                                                   lizzieLet1_4QNode_Bool_9QNode_Bool_d[0],
                                                                                                                                                                                                                                                                   t3a8o_destruct_d[0]}), lizzieLet1_4QNode_Bool_4QNode_Bool_d, lizzieLet1_4QNode_Bool_6QNode_Bool_1_d, lizzieLet1_4QNode_Bool_7QNode_Bool_d, t1a8m_destruct_d, lizzieLet1_4QNode_Bool_8QNode_Bool_d, t2a8n_destruct_d, lizzieLet1_4QNode_Bool_9QNode_Bool_d, t3a8o_destruct_d);
  assign {lizzieLet1_4QNode_Bool_4QNode_Bool_r,
          lizzieLet1_4QNode_Bool_6QNode_Bool_1_r,
          lizzieLet1_4QNode_Bool_7QNode_Bool_r,
          t1a8m_destruct_r,
          lizzieLet1_4QNode_Bool_8QNode_Bool_r,
          t2a8n_destruct_r,
          lizzieLet1_4QNode_Bool_9QNode_Bool_r,
          t3a8o_destruct_r} = {8 {(lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_r && lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_d[0])}};
  
  /* buf (Ty CT$wmAdd_Bool) : (lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3,CT$wmAdd_Bool) > (lizzieLet8_1_1_argbuf,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d;
  logic lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_r;
  assign lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_r = ((! lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d[0]) || lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d <= {115'd0,
                                                                                                                                                                                                                                                1'd0};
    else
      if (lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_r)
        lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d <= lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_d;
  CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_r = (! lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf :
                                    lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                                  1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf <= {115'd0,
                                                                                                                                                                                                                                                    1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_buf <= lizzieLet1_4QNode_Bool_4QNode_Bool_1lizzieLet1_4QNode_Bool_6QNode_Bool_1lizzieLet1_4QNode_Bool_7QNode_Bool_1t1a8m_1lizzieLet1_4QNode_Bool_8QNode_Bool_1t2a8n_1lizzieLet1_4QNode_Bool_9QNode_Bool_1t3a8o_1Lcall_$wmAdd_Bool3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QNode_Bool_4QNone_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_4QNone_Bool_r = ((! lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNode_Bool_4QNone_Bool_r)
        lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_4QNone_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf :
                                                          lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNode_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QNode_Bool_4QVal_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_4QVal_Bool_r = ((! lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNode_Bool_4QVal_Bool_r)
        lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_4QVal_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf :
                                                         lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNode_Bool_4QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_5,QTree_Bool) (lizzieLet1_6QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet1_4QNode_Bool_5QNone_Bool,Pointer_QTree_Bool),
                                                                                                                     (_35,Pointer_QTree_Bool),
                                                                                                                     (_34,Pointer_QTree_Bool),
                                                                                                                     (_33,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet1_6QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_5_d[0] && lizzieLet1_6QNode_Bool_d[0]))
      unique case (lizzieLet1_4QNode_Bool_5_d[2:1])
        2'd0: lizzieLet1_6QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_6QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_6QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_6QNode_Bool_onehotd = 4'd8;
        default: lizzieLet1_6QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_6QNode_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QNode_Bool_5QNone_Bool_d = {lizzieLet1_6QNode_Bool_d[16:1],
                                                 lizzieLet1_6QNode_Bool_onehotd[0]};
  assign _35_d = {lizzieLet1_6QNode_Bool_d[16:1],
                  lizzieLet1_6QNode_Bool_onehotd[1]};
  assign _34_d = {lizzieLet1_6QNode_Bool_d[16:1],
                  lizzieLet1_6QNode_Bool_onehotd[2]};
  assign _33_d = {lizzieLet1_6QNode_Bool_d[16:1],
                  lizzieLet1_6QNode_Bool_onehotd[3]};
  assign lizzieLet1_6QNode_Bool_r = (| (lizzieLet1_6QNode_Bool_onehotd & {_33_r,
                                                                          _34_r,
                                                                          _35_r,
                                                                          lizzieLet1_4QNode_Bool_5QNone_Bool_r}));
  assign lizzieLet1_4QNode_Bool_5_r = lizzieLet1_6QNode_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_5QNone_Bool,Pointer_QTree_Bool) > (lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet1_4QNode_Bool_5QNone_Bool_r = ((! lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QNode_Bool_5QNone_Bool_r)
        lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d <= lizzieLet1_4QNode_Bool_5QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_r = (! lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf :
                                                          lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_r && lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QNode_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_buf <= lizzieLet1_4QNode_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet1_4QNode_Bool_6,QTree_Bool) (lizzieLet1_8QNode_Bool,MyDTBool_Bool_Bool) > [(_32,MyDTBool_Bool_Bool),
                                                                                                                     (_31,MyDTBool_Bool_Bool),
                                                                                                                     (lizzieLet1_4QNode_Bool_6QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                                     (_30,MyDTBool_Bool_Bool)] */
  logic [3:0] lizzieLet1_8QNode_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_6_d[0] && lizzieLet1_8QNode_Bool_d[0]))
      unique case (lizzieLet1_4QNode_Bool_6_d[2:1])
        2'd0: lizzieLet1_8QNode_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_8QNode_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_8QNode_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_8QNode_Bool_onehotd = 4'd8;
        default: lizzieLet1_8QNode_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_8QNode_Bool_onehotd = 4'd0;
  assign _32_d = lizzieLet1_8QNode_Bool_onehotd[0];
  assign _31_d = lizzieLet1_8QNode_Bool_onehotd[1];
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_d = lizzieLet1_8QNode_Bool_onehotd[2];
  assign _30_d = lizzieLet1_8QNode_Bool_onehotd[3];
  assign lizzieLet1_8QNode_Bool_r = (| (lizzieLet1_8QNode_Bool_onehotd & {_30_r,
                                                                          lizzieLet1_4QNode_Bool_6QNode_Bool_r,
                                                                          _31_r,
                                                                          _32_r}));
  assign lizzieLet1_4QNode_Bool_6_r = lizzieLet1_8QNode_Bool_r;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (lizzieLet1_4QNode_Bool_6QNode_Bool,MyDTBool_Bool_Bool) > [(lizzieLet1_4QNode_Bool_6QNode_Bool_1,MyDTBool_Bool_Bool),
                                                                                          (lizzieLet1_4QNode_Bool_6QNode_Bool_2,MyDTBool_Bool_Bool)] */
  logic [1:0] lizzieLet1_4QNode_Bool_6QNode_Bool_emitted;
  logic [1:0] lizzieLet1_4QNode_Bool_6QNode_Bool_done;
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_1_d = (lizzieLet1_4QNode_Bool_6QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_6QNode_Bool_emitted[0]));
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_2_d = (lizzieLet1_4QNode_Bool_6QNode_Bool_d[0] && (! lizzieLet1_4QNode_Bool_6QNode_Bool_emitted[1]));
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_done = (lizzieLet1_4QNode_Bool_6QNode_Bool_emitted | ({lizzieLet1_4QNode_Bool_6QNode_Bool_2_d[0],
                                                                                                   lizzieLet1_4QNode_Bool_6QNode_Bool_1_d[0]} & {lizzieLet1_4QNode_Bool_6QNode_Bool_2_r,
                                                                                                                                                 lizzieLet1_4QNode_Bool_6QNode_Bool_1_r}));
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_r = (& lizzieLet1_4QNode_Bool_6QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_6QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QNode_Bool_6QNode_Bool_emitted <= (lizzieLet1_4QNode_Bool_6QNode_Bool_r ? 2'd0 :
                                                     lizzieLet1_4QNode_Bool_6QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet1_4QNode_Bool_6QNode_Bool_2,MyDTBool_Bool_Bool) > (lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d;
  logic lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_r;
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_2_r = ((! lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d[0]) || lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QNode_Bool_6QNode_Bool_2_r)
        lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d <= lizzieLet1_4QNode_Bool_6QNode_Bool_2_d;
  MyDTBool_Bool_Bool_t lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf;
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_r = (! lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_d = (lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf[0] ? lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf :
                                                          lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_r && lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QNode_Bool_6QNode_Bool_2_argbuf_r) && (! lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_buf <= lizzieLet1_4QNode_Bool_6QNode_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_7,QTree_Bool) (q1a8h_destruct,Pointer_QTree_Bool) > [(_29,Pointer_QTree_Bool),
                                                                                                             (_28,Pointer_QTree_Bool),
                                                                                                             (lizzieLet1_4QNode_Bool_7QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_27,Pointer_QTree_Bool)] */
  logic [3:0] q1a8h_destruct_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_7_d[0] && q1a8h_destruct_d[0]))
      unique case (lizzieLet1_4QNode_Bool_7_d[2:1])
        2'd0: q1a8h_destruct_onehotd = 4'd1;
        2'd1: q1a8h_destruct_onehotd = 4'd2;
        2'd2: q1a8h_destruct_onehotd = 4'd4;
        2'd3: q1a8h_destruct_onehotd = 4'd8;
        default: q1a8h_destruct_onehotd = 4'd0;
      endcase
    else q1a8h_destruct_onehotd = 4'd0;
  assign _29_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[0]};
  assign _28_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_7QNode_Bool_d = {q1a8h_destruct_d[16:1],
                                                 q1a8h_destruct_onehotd[2]};
  assign _27_d = {q1a8h_destruct_d[16:1], q1a8h_destruct_onehotd[3]};
  assign q1a8h_destruct_r = (| (q1a8h_destruct_onehotd & {_27_r,
                                                          lizzieLet1_4QNode_Bool_7QNode_Bool_r,
                                                          _28_r,
                                                          _29_r}));
  assign lizzieLet1_4QNode_Bool_7_r = q1a8h_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_8,QTree_Bool) (q2a8i_destruct,Pointer_QTree_Bool) > [(_26,Pointer_QTree_Bool),
                                                                                                             (_25,Pointer_QTree_Bool),
                                                                                                             (lizzieLet1_4QNode_Bool_8QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_24,Pointer_QTree_Bool)] */
  logic [3:0] q2a8i_destruct_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_8_d[0] && q2a8i_destruct_d[0]))
      unique case (lizzieLet1_4QNode_Bool_8_d[2:1])
        2'd0: q2a8i_destruct_onehotd = 4'd1;
        2'd1: q2a8i_destruct_onehotd = 4'd2;
        2'd2: q2a8i_destruct_onehotd = 4'd4;
        2'd3: q2a8i_destruct_onehotd = 4'd8;
        default: q2a8i_destruct_onehotd = 4'd0;
      endcase
    else q2a8i_destruct_onehotd = 4'd0;
  assign _26_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[0]};
  assign _25_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_8QNode_Bool_d = {q2a8i_destruct_d[16:1],
                                                 q2a8i_destruct_onehotd[2]};
  assign _24_d = {q2a8i_destruct_d[16:1], q2a8i_destruct_onehotd[3]};
  assign q2a8i_destruct_r = (| (q2a8i_destruct_onehotd & {_24_r,
                                                          lizzieLet1_4QNode_Bool_8QNode_Bool_r,
                                                          _25_r,
                                                          _26_r}));
  assign lizzieLet1_4QNode_Bool_8_r = q2a8i_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QNode_Bool_9,QTree_Bool) (q3a8j_destruct,Pointer_QTree_Bool) > [(_23,Pointer_QTree_Bool),
                                                                                                             (_22,Pointer_QTree_Bool),
                                                                                                             (lizzieLet1_4QNode_Bool_9QNode_Bool,Pointer_QTree_Bool),
                                                                                                             (_21,Pointer_QTree_Bool)] */
  logic [3:0] q3a8j_destruct_onehotd;
  always_comb
    if ((lizzieLet1_4QNode_Bool_9_d[0] && q3a8j_destruct_d[0]))
      unique case (lizzieLet1_4QNode_Bool_9_d[2:1])
        2'd0: q3a8j_destruct_onehotd = 4'd1;
        2'd1: q3a8j_destruct_onehotd = 4'd2;
        2'd2: q3a8j_destruct_onehotd = 4'd4;
        2'd3: q3a8j_destruct_onehotd = 4'd8;
        default: q3a8j_destruct_onehotd = 4'd0;
      endcase
    else q3a8j_destruct_onehotd = 4'd0;
  assign _23_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[0]};
  assign _22_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[1]};
  assign lizzieLet1_4QNode_Bool_9QNode_Bool_d = {q3a8j_destruct_d[16:1],
                                                 q3a8j_destruct_onehotd[2]};
  assign _21_d = {q3a8j_destruct_d[16:1], q3a8j_destruct_onehotd[3]};
  assign q3a8j_destruct_r = (| (q3a8j_destruct_onehotd & {_21_r,
                                                          lizzieLet1_4QNode_Bool_9QNode_Bool_r,
                                                          _22_r,
                                                          _23_r}));
  assign lizzieLet1_4QNode_Bool_9_r = q3a8j_destruct_r;
  
  /* fork (Ty QTree_Bool) : (lizzieLet1_4QVal_Bool,QTree_Bool) > [(lizzieLet1_4QVal_Bool_1,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_2,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_3,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_4,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_5,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_6,QTree_Bool),
                                                             (lizzieLet1_4QVal_Bool_7,QTree_Bool)] */
  logic [6:0] lizzieLet1_4QVal_Bool_emitted;
  logic [6:0] lizzieLet1_4QVal_Bool_done;
  assign lizzieLet1_4QVal_Bool_1_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[0]))};
  assign lizzieLet1_4QVal_Bool_2_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[1]))};
  assign lizzieLet1_4QVal_Bool_3_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[2]))};
  assign lizzieLet1_4QVal_Bool_4_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[3]))};
  assign lizzieLet1_4QVal_Bool_5_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[4]))};
  assign lizzieLet1_4QVal_Bool_6_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[5]))};
  assign lizzieLet1_4QVal_Bool_7_d = {lizzieLet1_4QVal_Bool_d[66:1],
                                      (lizzieLet1_4QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_emitted[6]))};
  assign lizzieLet1_4QVal_Bool_done = (lizzieLet1_4QVal_Bool_emitted | ({lizzieLet1_4QVal_Bool_7_d[0],
                                                                         lizzieLet1_4QVal_Bool_6_d[0],
                                                                         lizzieLet1_4QVal_Bool_5_d[0],
                                                                         lizzieLet1_4QVal_Bool_4_d[0],
                                                                         lizzieLet1_4QVal_Bool_3_d[0],
                                                                         lizzieLet1_4QVal_Bool_2_d[0],
                                                                         lizzieLet1_4QVal_Bool_1_d[0]} & {lizzieLet1_4QVal_Bool_7_r,
                                                                                                          lizzieLet1_4QVal_Bool_6_r,
                                                                                                          lizzieLet1_4QVal_Bool_5_r,
                                                                                                          lizzieLet1_4QVal_Bool_4_r,
                                                                                                          lizzieLet1_4QVal_Bool_3_r,
                                                                                                          lizzieLet1_4QVal_Bool_2_r,
                                                                                                          lizzieLet1_4QVal_Bool_1_r}));
  assign lizzieLet1_4QVal_Bool_r = (& lizzieLet1_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet1_4QVal_Bool_emitted <= 7'd0;
    else
      lizzieLet1_4QVal_Bool_emitted <= (lizzieLet1_4QVal_Bool_r ? 7'd0 :
                                        lizzieLet1_4QVal_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet1_4QVal_Bool_1QVal_Bool,QTree_Bool) > [(va8c_destruct,MyBool)] */
  assign va8c_destruct_d = {lizzieLet1_4QVal_Bool_1QVal_Bool_d[3:3],
                            lizzieLet1_4QVal_Bool_1QVal_Bool_d[0]};
  assign lizzieLet1_4QVal_Bool_1QVal_Bool_r = va8c_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet1_4QVal_Bool_2,QTree_Bool) (lizzieLet1_4QVal_Bool_1,QTree_Bool) > [(_20,QTree_Bool),
                                                                                                     (lizzieLet1_4QVal_Bool_1QVal_Bool,QTree_Bool),
                                                                                                     (_19,QTree_Bool),
                                                                                                     (_18,QTree_Bool)] */
  logic [3:0] lizzieLet1_4QVal_Bool_1_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_2_d[0] && lizzieLet1_4QVal_Bool_1_d[0]))
      unique case (lizzieLet1_4QVal_Bool_2_d[2:1])
        2'd0: lizzieLet1_4QVal_Bool_1_onehotd = 4'd1;
        2'd1: lizzieLet1_4QVal_Bool_1_onehotd = 4'd2;
        2'd2: lizzieLet1_4QVal_Bool_1_onehotd = 4'd4;
        2'd3: lizzieLet1_4QVal_Bool_1_onehotd = 4'd8;
        default: lizzieLet1_4QVal_Bool_1_onehotd = 4'd0;
      endcase
    else lizzieLet1_4QVal_Bool_1_onehotd = 4'd0;
  assign _20_d = {lizzieLet1_4QVal_Bool_1_d[66:1],
                  lizzieLet1_4QVal_Bool_1_onehotd[0]};
  assign lizzieLet1_4QVal_Bool_1QVal_Bool_d = {lizzieLet1_4QVal_Bool_1_d[66:1],
                                               lizzieLet1_4QVal_Bool_1_onehotd[1]};
  assign _19_d = {lizzieLet1_4QVal_Bool_1_d[66:1],
                  lizzieLet1_4QVal_Bool_1_onehotd[2]};
  assign _18_d = {lizzieLet1_4QVal_Bool_1_d[66:1],
                  lizzieLet1_4QVal_Bool_1_onehotd[3]};
  assign lizzieLet1_4QVal_Bool_1_r = (| (lizzieLet1_4QVal_Bool_1_onehotd & {_18_r,
                                                                            _19_r,
                                                                            lizzieLet1_4QVal_Bool_1QVal_Bool_r,
                                                                            _20_r}));
  assign lizzieLet1_4QVal_Bool_2_r = lizzieLet1_4QVal_Bool_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet1_4QVal_Bool_3,QTree_Bool) (lizzieLet1_3QVal_Bool,Go) > [(lizzieLet1_4QVal_Bool_3QNone_Bool,Go),
                                                                                   (lizzieLet1_4QVal_Bool_3QVal_Bool,Go),
                                                                                   (lizzieLet1_4QVal_Bool_3QNode_Bool,Go),
                                                                                   (lizzieLet1_4QVal_Bool_3QError_Bool,Go)] */
  logic [3:0] lizzieLet1_3QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_3_d[0] && lizzieLet1_3QVal_Bool_d[0]))
      unique case (lizzieLet1_4QVal_Bool_3_d[2:1])
        2'd0: lizzieLet1_3QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_3QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_3QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_3QVal_Bool_onehotd = 4'd8;
        default: lizzieLet1_3QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_3QVal_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QVal_Bool_3QNone_Bool_d = lizzieLet1_3QVal_Bool_onehotd[0];
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_d = lizzieLet1_3QVal_Bool_onehotd[1];
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_d = lizzieLet1_3QVal_Bool_onehotd[2];
  assign lizzieLet1_4QVal_Bool_3QError_Bool_d = lizzieLet1_3QVal_Bool_onehotd[3];
  assign lizzieLet1_3QVal_Bool_r = (| (lizzieLet1_3QVal_Bool_onehotd & {lizzieLet1_4QVal_Bool_3QError_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_3QNode_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_3QVal_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_3QNone_Bool_r}));
  assign lizzieLet1_4QVal_Bool_3_r = lizzieLet1_3QVal_Bool_r;
  
  /* fork (Ty Go) : (lizzieLet1_4QVal_Bool_3QError_Bool,Go) > [(lizzieLet1_4QVal_Bool_3QError_Bool_1,Go),
                                                          (lizzieLet1_4QVal_Bool_3QError_Bool_2,Go)] */
  logic [1:0] lizzieLet1_4QVal_Bool_3QError_Bool_emitted;
  logic [1:0] lizzieLet1_4QVal_Bool_3QError_Bool_done;
  assign lizzieLet1_4QVal_Bool_3QError_Bool_1_d = (lizzieLet1_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QError_Bool_emitted[0]));
  assign lizzieLet1_4QVal_Bool_3QError_Bool_2_d = (lizzieLet1_4QVal_Bool_3QError_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QError_Bool_emitted[1]));
  assign lizzieLet1_4QVal_Bool_3QError_Bool_done = (lizzieLet1_4QVal_Bool_3QError_Bool_emitted | ({lizzieLet1_4QVal_Bool_3QError_Bool_2_d[0],
                                                                                                   lizzieLet1_4QVal_Bool_3QError_Bool_1_d[0]} & {lizzieLet1_4QVal_Bool_3QError_Bool_2_r,
                                                                                                                                                 lizzieLet1_4QVal_Bool_3QError_Bool_1_r}));
  assign lizzieLet1_4QVal_Bool_3QError_Bool_r = (& lizzieLet1_4QVal_Bool_3QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QError_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QVal_Bool_3QError_Bool_emitted <= (lizzieLet1_4QVal_Bool_3QError_Bool_r ? 2'd0 :
                                                     lizzieLet1_4QVal_Bool_3QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet1_4QVal_Bool_3QError_Bool_1,Go)] > (lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet1_4QVal_Bool_3QError_Bool_1_d[0]}), lizzieLet1_4QVal_Bool_3QError_Bool_1_d);
  assign {lizzieLet1_4QVal_Bool_3QError_Bool_1_r} = {1 {(lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_r && lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet5_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_r = ((! lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                    1'd0};
    else
      if (lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_r)
        lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf :
                                    lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                      1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                        1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_3QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QVal_Bool_3QError_Bool_2,Go) > (lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QError_Bool_2_r = ((! lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_3QError_Bool_2_r)
        lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d <= lizzieLet1_4QVal_Bool_3QError_Bool_2_d;
  Go_t lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_r = (! lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_d = (lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf :
                                                          lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_r && lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_3QError_Bool_2_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_buf <= lizzieLet1_4QVal_Bool_3QError_Bool_2_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet1_4QVal_Bool_3QNode_Bool,Go) > [(lizzieLet1_4QVal_Bool_3QNode_Bool_1,Go),
                                                         (lizzieLet1_4QVal_Bool_3QNode_Bool_2,Go)] */
  logic [1:0] lizzieLet1_4QVal_Bool_3QNode_Bool_emitted;
  logic [1:0] lizzieLet1_4QVal_Bool_3QNode_Bool_done;
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_1_d = (lizzieLet1_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QNode_Bool_emitted[0]));
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_2_d = (lizzieLet1_4QVal_Bool_3QNode_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QNode_Bool_emitted[1]));
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_done = (lizzieLet1_4QVal_Bool_3QNode_Bool_emitted | ({lizzieLet1_4QVal_Bool_3QNode_Bool_2_d[0],
                                                                                                 lizzieLet1_4QVal_Bool_3QNode_Bool_1_d[0]} & {lizzieLet1_4QVal_Bool_3QNode_Bool_2_r,
                                                                                                                                              lizzieLet1_4QVal_Bool_3QNode_Bool_1_r}));
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_r = (& lizzieLet1_4QVal_Bool_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QVal_Bool_3QNode_Bool_emitted <= (lizzieLet1_4QVal_Bool_3QNode_Bool_r ? 2'd0 :
                                                    lizzieLet1_4QVal_Bool_3QNode_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet1_4QVal_Bool_3QNode_Bool_1,Go)] > (lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet1_4QVal_Bool_3QNode_Bool_1_d[0]}), lizzieLet1_4QVal_Bool_3QNode_Bool_1_d);
  assign {lizzieLet1_4QVal_Bool_3QNode_Bool_1_r} = {1 {(lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_r && lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool,QTree_Bool) > (lizzieLet4_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_r = ((! lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= {66'd0,
                                                                   1'd0};
    else
      if (lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_r)
        lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet4_1_argbuf_d = (lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                     1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                       1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_3QNode_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QVal_Bool_3QNode_Bool_2,Go) > (lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_2_r = ((! lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_3QNode_Bool_2_r)
        lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d <= lizzieLet1_4QVal_Bool_3QNode_Bool_2_d;
  Go_t lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_r = (! lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_d = (lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf :
                                                         lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_r && lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_3QNode_Bool_2_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_buf <= lizzieLet1_4QVal_Bool_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet1_4QVal_Bool_3QNone_Bool,Go) > (lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QNone_Bool_r = ((! lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_3QNone_Bool_r)
        lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_3QNone_Bool_d;
  Go_t lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf :
                                                         lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_3QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_3QNone_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet1_4QVal_Bool_3QVal_Bool,Go) > [(lizzieLet1_4QVal_Bool_3QVal_Bool_1,Go),
                                                        (lizzieLet1_4QVal_Bool_3QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet1_4QVal_Bool_3QVal_Bool_emitted;
  logic [1:0] lizzieLet1_4QVal_Bool_3QVal_Bool_done;
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_1_d = (lizzieLet1_4QVal_Bool_3QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QVal_Bool_emitted[0]));
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_2_d = (lizzieLet1_4QVal_Bool_3QVal_Bool_d[0] && (! lizzieLet1_4QVal_Bool_3QVal_Bool_emitted[1]));
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_done = (lizzieLet1_4QVal_Bool_3QVal_Bool_emitted | ({lizzieLet1_4QVal_Bool_3QVal_Bool_2_d[0],
                                                                                               lizzieLet1_4QVal_Bool_3QVal_Bool_1_d[0]} & {lizzieLet1_4QVal_Bool_3QVal_Bool_2_r,
                                                                                                                                           lizzieLet1_4QVal_Bool_3QVal_Bool_1_r}));
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_r = (& lizzieLet1_4QVal_Bool_3QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet1_4QVal_Bool_3QVal_Bool_emitted <= (lizzieLet1_4QVal_Bool_3QVal_Bool_r ? 2'd0 :
                                                   lizzieLet1_4QVal_Bool_3QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet1_4QVal_Bool_3QVal_Bool_1,Go) > (lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_1_r = ((! lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_3QVal_Bool_1_r)
        lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d <= lizzieLet1_4QVal_Bool_3QVal_Bool_1_d;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_r = (! lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf :
                                                        lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_buf <= lizzieLet1_4QVal_Bool_3QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
      Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : [(lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf,Go),
                                                            (lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf,MyDTBool_Bool_Bool),
                                                            (lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf,MyBool),
                                                            (va8c_1_argbuf,MyBool)] > (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) */
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d = TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_dc((& {lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_d[0],
                                                                                                                                       va8c_1_argbuf_d[0]}), lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_d, lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_d, lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_d, va8c_1_argbuf_d);
  assign {lizzieLet1_4QVal_Bool_3QVal_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_r,
          lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_r,
          va8c_1_argbuf_r} = {4 {(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet1_4QVal_Bool_3QVal_Bool_2,Go) > (lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d;
  logic lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_r;
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_2_r = ((! lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d[0]) || lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_3QVal_Bool_2_r)
        lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d <= lizzieLet1_4QVal_Bool_3QVal_Bool_2_d;
  Go_t lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_r = (! lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_d = (lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf :
                                                        lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_r && lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_3QVal_Bool_2_argbuf_r) && (! lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_buf <= lizzieLet1_4QVal_Bool_3QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QVal_Bool_4,QTree_Bool) (lizzieLet1_5QVal_Bool,Pointer_CT$wmAdd_Bool) > [(lizzieLet1_4QVal_Bool_4QNone_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                         (lizzieLet1_4QVal_Bool_4QVal_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                         (lizzieLet1_4QVal_Bool_4QNode_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                                         (lizzieLet1_4QVal_Bool_4QError_Bool,Pointer_CT$wmAdd_Bool)] */
  logic [3:0] lizzieLet1_5QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_4_d[0] && lizzieLet1_5QVal_Bool_d[0]))
      unique case (lizzieLet1_4QVal_Bool_4_d[2:1])
        2'd0: lizzieLet1_5QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_5QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_5QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_5QVal_Bool_onehotd = 4'd8;
        default: lizzieLet1_5QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_5QVal_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QVal_Bool_4QNone_Bool_d = {lizzieLet1_5QVal_Bool_d[16:1],
                                                lizzieLet1_5QVal_Bool_onehotd[0]};
  assign lizzieLet1_4QVal_Bool_4QVal_Bool_d = {lizzieLet1_5QVal_Bool_d[16:1],
                                               lizzieLet1_5QVal_Bool_onehotd[1]};
  assign lizzieLet1_4QVal_Bool_4QNode_Bool_d = {lizzieLet1_5QVal_Bool_d[16:1],
                                                lizzieLet1_5QVal_Bool_onehotd[2]};
  assign lizzieLet1_4QVal_Bool_4QError_Bool_d = {lizzieLet1_5QVal_Bool_d[16:1],
                                                 lizzieLet1_5QVal_Bool_onehotd[3]};
  assign lizzieLet1_5QVal_Bool_r = (| (lizzieLet1_5QVal_Bool_onehotd & {lizzieLet1_4QVal_Bool_4QError_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_4QNode_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_4QVal_Bool_r,
                                                                        lizzieLet1_4QVal_Bool_4QNone_Bool_r}));
  assign lizzieLet1_4QVal_Bool_4_r = lizzieLet1_5QVal_Bool_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QVal_Bool_4QError_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_4QError_Bool_r = ((! lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_4QError_Bool_r)
        lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_4QError_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf :
                                                          lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_4QError_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_4QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QVal_Bool_4QNode_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_4QNode_Bool_r = ((! lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_4QNode_Bool_r)
        lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_4QNode_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf :
                                                         lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_4QNode_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_4QNode_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QVal_Bool_4QNone_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_4QNone_Bool_r = ((! lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_4QNone_Bool_r)
        lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_4QNone_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf :
                                                         lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_4QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_4QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_4QVal_Bool_4QVal_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_4QVal_Bool_r = ((! lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_4QVal_Bool_r)
        lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_4QVal_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf :
                                                        lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_4QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_4QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_4QVal_Bool_5,QTree_Bool) (lizzieLet1_6QVal_Bool,Pointer_QTree_Bool) > [(lizzieLet1_4QVal_Bool_5QNone_Bool,Pointer_QTree_Bool),
                                                                                                                   (_17,Pointer_QTree_Bool),
                                                                                                                   (_16,Pointer_QTree_Bool),
                                                                                                                   (_15,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet1_6QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_5_d[0] && lizzieLet1_6QVal_Bool_d[0]))
      unique case (lizzieLet1_4QVal_Bool_5_d[2:1])
        2'd0: lizzieLet1_6QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_6QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_6QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_6QVal_Bool_onehotd = 4'd8;
        default: lizzieLet1_6QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_6QVal_Bool_onehotd = 4'd0;
  assign lizzieLet1_4QVal_Bool_5QNone_Bool_d = {lizzieLet1_6QVal_Bool_d[16:1],
                                                lizzieLet1_6QVal_Bool_onehotd[0]};
  assign _17_d = {lizzieLet1_6QVal_Bool_d[16:1],
                  lizzieLet1_6QVal_Bool_onehotd[1]};
  assign _16_d = {lizzieLet1_6QVal_Bool_d[16:1],
                  lizzieLet1_6QVal_Bool_onehotd[2]};
  assign _15_d = {lizzieLet1_6QVal_Bool_d[16:1],
                  lizzieLet1_6QVal_Bool_onehotd[3]};
  assign lizzieLet1_6QVal_Bool_r = (| (lizzieLet1_6QVal_Bool_onehotd & {_15_r,
                                                                        _16_r,
                                                                        _17_r,
                                                                        lizzieLet1_4QVal_Bool_5QNone_Bool_r}));
  assign lizzieLet1_4QVal_Bool_5_r = lizzieLet1_6QVal_Bool_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet1_4QVal_Bool_5QNone_Bool,Pointer_QTree_Bool) > (lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_5QNone_Bool_r = ((! lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_5QNone_Bool_r)
        lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_5QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf :
                                                         lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_5QNone_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet1_4QVal_Bool_6,QTree_Bool) (lizzieLet1_8QVal_Bool,MyDTBool_Bool_Bool) > [(_14,MyDTBool_Bool_Bool),
                                                                                                                   (lizzieLet1_4QVal_Bool_6QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                                   (_13,MyDTBool_Bool_Bool),
                                                                                                                   (_12,MyDTBool_Bool_Bool)] */
  logic [3:0] lizzieLet1_8QVal_Bool_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_6_d[0] && lizzieLet1_8QVal_Bool_d[0]))
      unique case (lizzieLet1_4QVal_Bool_6_d[2:1])
        2'd0: lizzieLet1_8QVal_Bool_onehotd = 4'd1;
        2'd1: lizzieLet1_8QVal_Bool_onehotd = 4'd2;
        2'd2: lizzieLet1_8QVal_Bool_onehotd = 4'd4;
        2'd3: lizzieLet1_8QVal_Bool_onehotd = 4'd8;
        default: lizzieLet1_8QVal_Bool_onehotd = 4'd0;
      endcase
    else lizzieLet1_8QVal_Bool_onehotd = 4'd0;
  assign _14_d = lizzieLet1_8QVal_Bool_onehotd[0];
  assign lizzieLet1_4QVal_Bool_6QVal_Bool_d = lizzieLet1_8QVal_Bool_onehotd[1];
  assign _13_d = lizzieLet1_8QVal_Bool_onehotd[2];
  assign _12_d = lizzieLet1_8QVal_Bool_onehotd[3];
  assign lizzieLet1_8QVal_Bool_r = (| (lizzieLet1_8QVal_Bool_onehotd & {_12_r,
                                                                        _13_r,
                                                                        lizzieLet1_4QVal_Bool_6QVal_Bool_r,
                                                                        _14_r}));
  assign lizzieLet1_4QVal_Bool_6_r = lizzieLet1_8QVal_Bool_r;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet1_4QVal_Bool_6QVal_Bool,MyDTBool_Bool_Bool) > (lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_6QVal_Bool_r = ((! lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet1_4QVal_Bool_6QVal_Bool_r)
        lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_6QVal_Bool_d;
  MyDTBool_Bool_Bool_t lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf :
                                                        lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet1_4QVal_Bool_6QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_6QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet1_4QVal_Bool_7,QTree_Bool) (v1a8b_destruct,MyBool) > [(_11,MyBool),
                                                                                    (lizzieLet1_4QVal_Bool_7QVal_Bool,MyBool),
                                                                                    (_10,MyBool),
                                                                                    (_9,MyBool)] */
  logic [3:0] v1a8b_destruct_onehotd;
  always_comb
    if ((lizzieLet1_4QVal_Bool_7_d[0] && v1a8b_destruct_d[0]))
      unique case (lizzieLet1_4QVal_Bool_7_d[2:1])
        2'd0: v1a8b_destruct_onehotd = 4'd1;
        2'd1: v1a8b_destruct_onehotd = 4'd2;
        2'd2: v1a8b_destruct_onehotd = 4'd4;
        2'd3: v1a8b_destruct_onehotd = 4'd8;
        default: v1a8b_destruct_onehotd = 4'd0;
      endcase
    else v1a8b_destruct_onehotd = 4'd0;
  assign _11_d = {v1a8b_destruct_d[1:1], v1a8b_destruct_onehotd[0]};
  assign lizzieLet1_4QVal_Bool_7QVal_Bool_d = {v1a8b_destruct_d[1:1],
                                               v1a8b_destruct_onehotd[1]};
  assign _10_d = {v1a8b_destruct_d[1:1], v1a8b_destruct_onehotd[2]};
  assign _9_d = {v1a8b_destruct_d[1:1], v1a8b_destruct_onehotd[3]};
  assign v1a8b_destruct_r = (| (v1a8b_destruct_onehotd & {_9_r,
                                                          _10_r,
                                                          lizzieLet1_4QVal_Bool_7QVal_Bool_r,
                                                          _11_r}));
  assign lizzieLet1_4QVal_Bool_7_r = v1a8b_destruct_r;
  
  /* buf (Ty MyBool) : (lizzieLet1_4QVal_Bool_7QVal_Bool,MyBool) > (lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf,MyBool) */
  MyBool_t lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d;
  logic lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_r;
  assign lizzieLet1_4QVal_Bool_7QVal_Bool_r = ((! lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d[0]) || lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_4QVal_Bool_7QVal_Bool_r)
        lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d <= lizzieLet1_4QVal_Bool_7QVal_Bool_d;
  MyBool_t lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf;
  assign lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_r = (! lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf[0]);
  assign lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_d = (lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf[0] ? lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf :
                                                        lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_r && lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf[0]))
        lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet1_4QVal_Bool_7QVal_Bool_1_argbuf_r) && (! lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf[0])))
        lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_buf <= lizzieLet1_4QVal_Bool_7QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_5,QTree_Bool) (sc_0_goMux_mux,Pointer_CT$wmAdd_Bool) > [(lizzieLet1_5QNone_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                       (lizzieLet1_5QVal_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                       (lizzieLet1_5QNode_Bool,Pointer_CT$wmAdd_Bool),
                                                                                                       (lizzieLet1_5QError_Bool,Pointer_CT$wmAdd_Bool)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet1_5_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet1_5_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet1_5QNone_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet1_5QVal_Bool_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet1_5QNode_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet1_5QError_Bool_d = {sc_0_goMux_mux_d[16:1],
                                      sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet1_5QError_Bool_r,
                                                          lizzieLet1_5QNode_Bool_r,
                                                          lizzieLet1_5QVal_Bool_r,
                                                          lizzieLet1_5QNone_Bool_r}));
  assign lizzieLet1_5_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_5QError_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_5QError_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QError_Bool_bufchan_d;
  logic lizzieLet1_5QError_Bool_bufchan_r;
  assign lizzieLet1_5QError_Bool_r = ((! lizzieLet1_5QError_Bool_bufchan_d[0]) || lizzieLet1_5QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_5QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_5QError_Bool_r)
        lizzieLet1_5QError_Bool_bufchan_d <= lizzieLet1_5QError_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QError_Bool_bufchan_buf;
  assign lizzieLet1_5QError_Bool_bufchan_r = (! lizzieLet1_5QError_Bool_bufchan_buf[0]);
  assign lizzieLet1_5QError_Bool_1_argbuf_d = (lizzieLet1_5QError_Bool_bufchan_buf[0] ? lizzieLet1_5QError_Bool_bufchan_buf :
                                               lizzieLet1_5QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_5QError_Bool_1_argbuf_r && lizzieLet1_5QError_Bool_bufchan_buf[0]))
        lizzieLet1_5QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_5QError_Bool_1_argbuf_r) && (! lizzieLet1_5QError_Bool_bufchan_buf[0])))
        lizzieLet1_5QError_Bool_bufchan_buf <= lizzieLet1_5QError_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (lizzieLet1_5QNone_Bool,Pointer_CT$wmAdd_Bool) > (lizzieLet1_5QNone_Bool_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QNone_Bool_bufchan_d;
  logic lizzieLet1_5QNone_Bool_bufchan_r;
  assign lizzieLet1_5QNone_Bool_r = ((! lizzieLet1_5QNone_Bool_bufchan_d[0]) || lizzieLet1_5QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_5QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_5QNone_Bool_r)
        lizzieLet1_5QNone_Bool_bufchan_d <= lizzieLet1_5QNone_Bool_d;
  Pointer_CT$wmAdd_Bool_t lizzieLet1_5QNone_Bool_bufchan_buf;
  assign lizzieLet1_5QNone_Bool_bufchan_r = (! lizzieLet1_5QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_5QNone_Bool_1_argbuf_d = (lizzieLet1_5QNone_Bool_bufchan_buf[0] ? lizzieLet1_5QNone_Bool_bufchan_buf :
                                              lizzieLet1_5QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_5QNone_Bool_1_argbuf_r && lizzieLet1_5QNone_Bool_bufchan_buf[0]))
        lizzieLet1_5QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_5QNone_Bool_1_argbuf_r) && (! lizzieLet1_5QNone_Bool_bufchan_buf[0])))
        lizzieLet1_5QNone_Bool_bufchan_buf <= lizzieLet1_5QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_6,QTree_Bool) (w1sic_1_2,Pointer_QTree_Bool) > [(_8,Pointer_QTree_Bool),
                                                                                            (lizzieLet1_6QVal_Bool,Pointer_QTree_Bool),
                                                                                            (lizzieLet1_6QNode_Bool,Pointer_QTree_Bool),
                                                                                            (_7,Pointer_QTree_Bool)] */
  logic [3:0] w1sic_1_2_onehotd;
  always_comb
    if ((lizzieLet1_6_d[0] && w1sic_1_2_d[0]))
      unique case (lizzieLet1_6_d[2:1])
        2'd0: w1sic_1_2_onehotd = 4'd1;
        2'd1: w1sic_1_2_onehotd = 4'd2;
        2'd2: w1sic_1_2_onehotd = 4'd4;
        2'd3: w1sic_1_2_onehotd = 4'd8;
        default: w1sic_1_2_onehotd = 4'd0;
      endcase
    else w1sic_1_2_onehotd = 4'd0;
  assign _8_d = {w1sic_1_2_d[16:1], w1sic_1_2_onehotd[0]};
  assign lizzieLet1_6QVal_Bool_d = {w1sic_1_2_d[16:1],
                                    w1sic_1_2_onehotd[1]};
  assign lizzieLet1_6QNode_Bool_d = {w1sic_1_2_d[16:1],
                                     w1sic_1_2_onehotd[2]};
  assign _7_d = {w1sic_1_2_d[16:1], w1sic_1_2_onehotd[3]};
  assign w1sic_1_2_r = (| (w1sic_1_2_onehotd & {_7_r,
                                                lizzieLet1_6QNode_Bool_r,
                                                lizzieLet1_6QVal_Bool_r,
                                                _8_r}));
  assign lizzieLet1_6_r = w1sic_1_2_r;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet1_7,QTree_Bool) (w2sid_1_2,Pointer_QTree_Bool) > [(lizzieLet1_7QNone_Bool,Pointer_QTree_Bool),
                                                                                            (_6,Pointer_QTree_Bool),
                                                                                            (_5,Pointer_QTree_Bool),
                                                                                            (_4,Pointer_QTree_Bool)] */
  logic [3:0] w2sid_1_2_onehotd;
  always_comb
    if ((lizzieLet1_7_d[0] && w2sid_1_2_d[0]))
      unique case (lizzieLet1_7_d[2:1])
        2'd0: w2sid_1_2_onehotd = 4'd1;
        2'd1: w2sid_1_2_onehotd = 4'd2;
        2'd2: w2sid_1_2_onehotd = 4'd4;
        2'd3: w2sid_1_2_onehotd = 4'd8;
        default: w2sid_1_2_onehotd = 4'd0;
      endcase
    else w2sid_1_2_onehotd = 4'd0;
  assign lizzieLet1_7QNone_Bool_d = {w2sid_1_2_d[16:1],
                                     w2sid_1_2_onehotd[0]};
  assign _6_d = {w2sid_1_2_d[16:1], w2sid_1_2_onehotd[1]};
  assign _5_d = {w2sid_1_2_d[16:1], w2sid_1_2_onehotd[2]};
  assign _4_d = {w2sid_1_2_d[16:1], w2sid_1_2_onehotd[3]};
  assign w2sid_1_2_r = (| (w2sid_1_2_onehotd & {_4_r,
                                                _5_r,
                                                _6_r,
                                                lizzieLet1_7QNone_Bool_r}));
  assign lizzieLet1_7_r = w2sid_1_2_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet1_7QNone_Bool,Pointer_QTree_Bool) > (lizzieLet1_7QNone_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet1_7QNone_Bool_bufchan_d;
  logic lizzieLet1_7QNone_Bool_bufchan_r;
  assign lizzieLet1_7QNone_Bool_r = ((! lizzieLet1_7QNone_Bool_bufchan_d[0]) || lizzieLet1_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet1_7QNone_Bool_r)
        lizzieLet1_7QNone_Bool_bufchan_d <= lizzieLet1_7QNone_Bool_d;
  Pointer_QTree_Bool_t lizzieLet1_7QNone_Bool_bufchan_buf;
  assign lizzieLet1_7QNone_Bool_bufchan_r = (! lizzieLet1_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet1_7QNone_Bool_1_argbuf_d = (lizzieLet1_7QNone_Bool_bufchan_buf[0] ? lizzieLet1_7QNone_Bool_bufchan_buf :
                                              lizzieLet1_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_7QNone_Bool_1_argbuf_r && lizzieLet1_7QNone_Bool_bufchan_buf[0]))
        lizzieLet1_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_7QNone_Bool_1_argbuf_r) && (! lizzieLet1_7QNone_Bool_bufchan_buf[0])))
        lizzieLet1_7QNone_Bool_bufchan_buf <= lizzieLet1_7QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet1_8,QTree_Bool) (wsib_1_goMux_mux,MyDTBool_Bool_Bool) > [(_3,MyDTBool_Bool_Bool),
                                                                                                   (lizzieLet1_8QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                   (lizzieLet1_8QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                   (_2,MyDTBool_Bool_Bool)] */
  logic [3:0] wsib_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet1_8_d[0] && wsib_1_goMux_mux_d[0]))
      unique case (lizzieLet1_8_d[2:1])
        2'd0: wsib_1_goMux_mux_onehotd = 4'd1;
        2'd1: wsib_1_goMux_mux_onehotd = 4'd2;
        2'd2: wsib_1_goMux_mux_onehotd = 4'd4;
        2'd3: wsib_1_goMux_mux_onehotd = 4'd8;
        default: wsib_1_goMux_mux_onehotd = 4'd0;
      endcase
    else wsib_1_goMux_mux_onehotd = 4'd0;
  assign _3_d = wsib_1_goMux_mux_onehotd[0];
  assign lizzieLet1_8QVal_Bool_d = wsib_1_goMux_mux_onehotd[1];
  assign lizzieLet1_8QNode_Bool_d = wsib_1_goMux_mux_onehotd[2];
  assign _2_d = wsib_1_goMux_mux_onehotd[3];
  assign wsib_1_goMux_mux_r = (| (wsib_1_goMux_mux_onehotd & {_2_r,
                                                              lizzieLet1_8QNode_Bool_r,
                                                              lizzieLet1_8QVal_Bool_r,
                                                              _3_r}));
  assign lizzieLet1_8_r = wsib_1_goMux_mux_r;
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool0) : (lizzieLet24_1Lcall_main_mask_Bool0,CTmain_mask_Bool) > [(es_1_destruct,Pointer_QTree_Bool),
                                                                                                 (es_2_3_destruct,Pointer_QTree_Bool),
                                                                                                 (es_3_4_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_9_destruct,Pointer_CTmain_mask_Bool)] */
  logic [3:0] lizzieLet24_1Lcall_main_mask_Bool0_emitted;
  logic [3:0] lizzieLet24_1Lcall_main_mask_Bool0_done;
  assign es_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool0_d[19:4],
                            (lizzieLet24_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool0_emitted[0]))};
  assign es_2_3_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool0_d[35:20],
                              (lizzieLet24_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool0_emitted[1]))};
  assign es_3_4_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool0_d[51:36],
                              (lizzieLet24_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool0_emitted[2]))};
  assign sc_0_9_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool0_d[67:52],
                              (lizzieLet24_1Lcall_main_mask_Bool0_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool0_emitted[3]))};
  assign lizzieLet24_1Lcall_main_mask_Bool0_done = (lizzieLet24_1Lcall_main_mask_Bool0_emitted | ({sc_0_9_destruct_d[0],
                                                                                                   es_3_4_destruct_d[0],
                                                                                                   es_2_3_destruct_d[0],
                                                                                                   es_1_destruct_d[0]} & {sc_0_9_destruct_r,
                                                                                                                          es_3_4_destruct_r,
                                                                                                                          es_2_3_destruct_r,
                                                                                                                          es_1_destruct_r}));
  assign lizzieLet24_1Lcall_main_mask_Bool0_r = (& lizzieLet24_1Lcall_main_mask_Bool0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_main_mask_Bool0_emitted <= 4'd0;
    else
      lizzieLet24_1Lcall_main_mask_Bool0_emitted <= (lizzieLet24_1Lcall_main_mask_Bool0_r ? 4'd0 :
                                                     lizzieLet24_1Lcall_main_mask_Bool0_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool1) : (lizzieLet24_1Lcall_main_mask_Bool1,CTmain_mask_Bool) > [(es_2_2_destruct,Pointer_QTree_Bool),
                                                                                                 (es_3_3_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_8_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1a8x_3_destruct,Pointer_QTree_Bool),
                                                                                                 (q1a8s_3_destruct,Pointer_MaskQTree)] */
  logic [4:0] lizzieLet24_1Lcall_main_mask_Bool1_emitted;
  logic [4:0] lizzieLet24_1Lcall_main_mask_Bool1_done;
  assign es_2_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool1_d[19:4],
                              (lizzieLet24_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool1_emitted[0]))};
  assign es_3_3_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool1_d[35:20],
                              (lizzieLet24_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool1_emitted[1]))};
  assign sc_0_8_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool1_d[51:36],
                              (lizzieLet24_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool1_emitted[2]))};
  assign t1a8x_3_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool1_d[67:52],
                               (lizzieLet24_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool1_emitted[3]))};
  assign q1a8s_3_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool1_d[83:68],
                               (lizzieLet24_1Lcall_main_mask_Bool1_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool1_emitted[4]))};
  assign lizzieLet24_1Lcall_main_mask_Bool1_done = (lizzieLet24_1Lcall_main_mask_Bool1_emitted | ({q1a8s_3_destruct_d[0],
                                                                                                   t1a8x_3_destruct_d[0],
                                                                                                   sc_0_8_destruct_d[0],
                                                                                                   es_3_3_destruct_d[0],
                                                                                                   es_2_2_destruct_d[0]} & {q1a8s_3_destruct_r,
                                                                                                                            t1a8x_3_destruct_r,
                                                                                                                            sc_0_8_destruct_r,
                                                                                                                            es_3_3_destruct_r,
                                                                                                                            es_2_2_destruct_r}));
  assign lizzieLet24_1Lcall_main_mask_Bool1_r = (& lizzieLet24_1Lcall_main_mask_Bool1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_main_mask_Bool1_emitted <= 5'd0;
    else
      lizzieLet24_1Lcall_main_mask_Bool1_emitted <= (lizzieLet24_1Lcall_main_mask_Bool1_r ? 5'd0 :
                                                     lizzieLet24_1Lcall_main_mask_Bool1_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool2) : (lizzieLet24_1Lcall_main_mask_Bool2,CTmain_mask_Bool) > [(es_3_2_destruct,Pointer_QTree_Bool),
                                                                                                 (sc_0_7_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1a8x_2_destruct,Pointer_QTree_Bool),
                                                                                                 (q1a8s_2_destruct,Pointer_MaskQTree),
                                                                                                 (t2a8y_2_destruct,Pointer_QTree_Bool),
                                                                                                 (q2a8t_2_destruct,Pointer_MaskQTree)] */
  logic [5:0] lizzieLet24_1Lcall_main_mask_Bool2_emitted;
  logic [5:0] lizzieLet24_1Lcall_main_mask_Bool2_done;
  assign es_3_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[19:4],
                              (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[0]))};
  assign sc_0_7_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[35:20],
                              (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[1]))};
  assign t1a8x_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[51:36],
                               (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[2]))};
  assign q1a8s_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[67:52],
                               (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[3]))};
  assign t2a8y_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[83:68],
                               (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[4]))};
  assign q2a8t_2_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool2_d[99:84],
                               (lizzieLet24_1Lcall_main_mask_Bool2_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool2_emitted[5]))};
  assign lizzieLet24_1Lcall_main_mask_Bool2_done = (lizzieLet24_1Lcall_main_mask_Bool2_emitted | ({q2a8t_2_destruct_d[0],
                                                                                                   t2a8y_2_destruct_d[0],
                                                                                                   q1a8s_2_destruct_d[0],
                                                                                                   t1a8x_2_destruct_d[0],
                                                                                                   sc_0_7_destruct_d[0],
                                                                                                   es_3_2_destruct_d[0]} & {q2a8t_2_destruct_r,
                                                                                                                            t2a8y_2_destruct_r,
                                                                                                                            q1a8s_2_destruct_r,
                                                                                                                            t1a8x_2_destruct_r,
                                                                                                                            sc_0_7_destruct_r,
                                                                                                                            es_3_2_destruct_r}));
  assign lizzieLet24_1Lcall_main_mask_Bool2_r = (& lizzieLet24_1Lcall_main_mask_Bool2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_main_mask_Bool2_emitted <= 6'd0;
    else
      lizzieLet24_1Lcall_main_mask_Bool2_emitted <= (lizzieLet24_1Lcall_main_mask_Bool2_r ? 6'd0 :
                                                     lizzieLet24_1Lcall_main_mask_Bool2_done);
  
  /* destruct (Ty CTmain_mask_Bool,
          Dcon Lcall_main_mask_Bool3) : (lizzieLet24_1Lcall_main_mask_Bool3,CTmain_mask_Bool) > [(sc_0_6_destruct,Pointer_CTmain_mask_Bool),
                                                                                                 (t1a8x_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q1a8s_1_destruct,Pointer_MaskQTree),
                                                                                                 (t2a8y_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q2a8t_1_destruct,Pointer_MaskQTree),
                                                                                                 (t3a8z_1_destruct,Pointer_QTree_Bool),
                                                                                                 (q3a8u_1_destruct,Pointer_MaskQTree)] */
  logic [6:0] lizzieLet24_1Lcall_main_mask_Bool3_emitted;
  logic [6:0] lizzieLet24_1Lcall_main_mask_Bool3_done;
  assign sc_0_6_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[19:4],
                              (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[0]))};
  assign t1a8x_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[35:20],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[1]))};
  assign q1a8s_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[51:36],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[2]))};
  assign t2a8y_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[67:52],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[3]))};
  assign q2a8t_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[83:68],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[4]))};
  assign t3a8z_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[99:84],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[5]))};
  assign q3a8u_1_destruct_d = {lizzieLet24_1Lcall_main_mask_Bool3_d[115:100],
                               (lizzieLet24_1Lcall_main_mask_Bool3_d[0] && (! lizzieLet24_1Lcall_main_mask_Bool3_emitted[6]))};
  assign lizzieLet24_1Lcall_main_mask_Bool3_done = (lizzieLet24_1Lcall_main_mask_Bool3_emitted | ({q3a8u_1_destruct_d[0],
                                                                                                   t3a8z_1_destruct_d[0],
                                                                                                   q2a8t_1_destruct_d[0],
                                                                                                   t2a8y_1_destruct_d[0],
                                                                                                   q1a8s_1_destruct_d[0],
                                                                                                   t1a8x_1_destruct_d[0],
                                                                                                   sc_0_6_destruct_d[0]} & {q3a8u_1_destruct_r,
                                                                                                                            t3a8z_1_destruct_r,
                                                                                                                            q2a8t_1_destruct_r,
                                                                                                                            t2a8y_1_destruct_r,
                                                                                                                            q1a8s_1_destruct_r,
                                                                                                                            t1a8x_1_destruct_r,
                                                                                                                            sc_0_6_destruct_r}));
  assign lizzieLet24_1Lcall_main_mask_Bool3_r = (& lizzieLet24_1Lcall_main_mask_Bool3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_main_mask_Bool3_emitted <= 7'd0;
    else
      lizzieLet24_1Lcall_main_mask_Bool3_emitted <= (lizzieLet24_1Lcall_main_mask_Bool3_r ? 7'd0 :
                                                     lizzieLet24_1Lcall_main_mask_Bool3_done);
  
  /* demux (Ty CTmain_mask_Bool,
       Ty CTmain_mask_Bool) : (lizzieLet24_2,CTmain_mask_Bool) (lizzieLet24_1,CTmain_mask_Bool) > [(_1,CTmain_mask_Bool),
                                                                                                   (lizzieLet24_1Lcall_main_mask_Bool3,CTmain_mask_Bool),
                                                                                                   (lizzieLet24_1Lcall_main_mask_Bool2,CTmain_mask_Bool),
                                                                                                   (lizzieLet24_1Lcall_main_mask_Bool1,CTmain_mask_Bool),
                                                                                                   (lizzieLet24_1Lcall_main_mask_Bool0,CTmain_mask_Bool)] */
  logic [4:0] lizzieLet24_1_onehotd;
  always_comb
    if ((lizzieLet24_2_d[0] && lizzieLet24_1_d[0]))
      unique case (lizzieLet24_2_d[3:1])
        3'd0: lizzieLet24_1_onehotd = 5'd1;
        3'd1: lizzieLet24_1_onehotd = 5'd2;
        3'd2: lizzieLet24_1_onehotd = 5'd4;
        3'd3: lizzieLet24_1_onehotd = 5'd8;
        3'd4: lizzieLet24_1_onehotd = 5'd16;
        default: lizzieLet24_1_onehotd = 5'd0;
      endcase
    else lizzieLet24_1_onehotd = 5'd0;
  assign _1_d = {lizzieLet24_1_d[115:1], lizzieLet24_1_onehotd[0]};
  assign lizzieLet24_1Lcall_main_mask_Bool3_d = {lizzieLet24_1_d[115:1],
                                                 lizzieLet24_1_onehotd[1]};
  assign lizzieLet24_1Lcall_main_mask_Bool2_d = {lizzieLet24_1_d[115:1],
                                                 lizzieLet24_1_onehotd[2]};
  assign lizzieLet24_1Lcall_main_mask_Bool1_d = {lizzieLet24_1_d[115:1],
                                                 lizzieLet24_1_onehotd[3]};
  assign lizzieLet24_1Lcall_main_mask_Bool0_d = {lizzieLet24_1_d[115:1],
                                                 lizzieLet24_1_onehotd[4]};
  assign lizzieLet24_1_r = (| (lizzieLet24_1_onehotd & {lizzieLet24_1Lcall_main_mask_Bool0_r,
                                                        lizzieLet24_1Lcall_main_mask_Bool1_r,
                                                        lizzieLet24_1Lcall_main_mask_Bool2_r,
                                                        lizzieLet24_1Lcall_main_mask_Bool3_r,
                                                        _1_r}));
  assign lizzieLet24_2_r = lizzieLet24_1_r;
  
  /* demux (Ty CTmain_mask_Bool,
       Ty Go) : (lizzieLet24_3,CTmain_mask_Bool) (go_8_goMux_data,Go) > [(_0,Go),
                                                                         (lizzieLet24_3Lcall_main_mask_Bool3,Go),
                                                                         (lizzieLet24_3Lcall_main_mask_Bool2,Go),
                                                                         (lizzieLet24_3Lcall_main_mask_Bool1,Go),
                                                                         (lizzieLet24_3Lcall_main_mask_Bool0,Go)] */
  logic [4:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet24_3_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet24_3_d[3:1])
        3'd0: go_8_goMux_data_onehotd = 5'd1;
        3'd1: go_8_goMux_data_onehotd = 5'd2;
        3'd2: go_8_goMux_data_onehotd = 5'd4;
        3'd3: go_8_goMux_data_onehotd = 5'd8;
        3'd4: go_8_goMux_data_onehotd = 5'd16;
        default: go_8_goMux_data_onehotd = 5'd0;
      endcase
    else go_8_goMux_data_onehotd = 5'd0;
  assign _0_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet24_3Lcall_main_mask_Bool3_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet24_3Lcall_main_mask_Bool2_d = go_8_goMux_data_onehotd[2];
  assign lizzieLet24_3Lcall_main_mask_Bool1_d = go_8_goMux_data_onehotd[3];
  assign lizzieLet24_3Lcall_main_mask_Bool0_d = go_8_goMux_data_onehotd[4];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet24_3Lcall_main_mask_Bool0_r,
                                                            lizzieLet24_3Lcall_main_mask_Bool1_r,
                                                            lizzieLet24_3Lcall_main_mask_Bool2_r,
                                                            lizzieLet24_3Lcall_main_mask_Bool3_r,
                                                            _0_r}));
  assign lizzieLet24_3_r = go_8_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_main_mask_Bool0,Go) > (lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d;
  logic lizzieLet24_3Lcall_main_mask_Bool0_bufchan_r;
  assign lizzieLet24_3Lcall_main_mask_Bool0_r = ((! lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d[0]) || lizzieLet24_3Lcall_main_mask_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_main_mask_Bool0_r)
        lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d <= lizzieLet24_3Lcall_main_mask_Bool0_d;
  Go_t lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf;
  assign lizzieLet24_3Lcall_main_mask_Bool0_bufchan_r = (! lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_d = (lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf[0] ? lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf :
                                                          lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_r && lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf[0]))
        lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_main_mask_Bool0_1_argbuf_r) && (! lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf[0])))
        lizzieLet24_3Lcall_main_mask_Bool0_bufchan_buf <= lizzieLet24_3Lcall_main_mask_Bool0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_main_mask_Bool1,Go) > (lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d;
  logic lizzieLet24_3Lcall_main_mask_Bool1_bufchan_r;
  assign lizzieLet24_3Lcall_main_mask_Bool1_r = ((! lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d[0]) || lizzieLet24_3Lcall_main_mask_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_main_mask_Bool1_r)
        lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d <= lizzieLet24_3Lcall_main_mask_Bool1_d;
  Go_t lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf;
  assign lizzieLet24_3Lcall_main_mask_Bool1_bufchan_r = (! lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_d = (lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf[0] ? lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf :
                                                          lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_r && lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf[0]))
        lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_main_mask_Bool1_1_argbuf_r) && (! lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf[0])))
        lizzieLet24_3Lcall_main_mask_Bool1_bufchan_buf <= lizzieLet24_3Lcall_main_mask_Bool1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_main_mask_Bool2,Go) > (lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d;
  logic lizzieLet24_3Lcall_main_mask_Bool2_bufchan_r;
  assign lizzieLet24_3Lcall_main_mask_Bool2_r = ((! lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d[0]) || lizzieLet24_3Lcall_main_mask_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_main_mask_Bool2_r)
        lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d <= lizzieLet24_3Lcall_main_mask_Bool2_d;
  Go_t lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf;
  assign lizzieLet24_3Lcall_main_mask_Bool2_bufchan_r = (! lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_d = (lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf[0] ? lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf :
                                                          lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_r && lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf[0]))
        lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_main_mask_Bool2_1_argbuf_r) && (! lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf[0])))
        lizzieLet24_3Lcall_main_mask_Bool2_bufchan_buf <= lizzieLet24_3Lcall_main_mask_Bool2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_main_mask_Bool3,Go) > (lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d;
  logic lizzieLet24_3Lcall_main_mask_Bool3_bufchan_r;
  assign lizzieLet24_3Lcall_main_mask_Bool3_r = ((! lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d[0]) || lizzieLet24_3Lcall_main_mask_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_main_mask_Bool3_r)
        lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d <= lizzieLet24_3Lcall_main_mask_Bool3_d;
  Go_t lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf;
  assign lizzieLet24_3Lcall_main_mask_Bool3_bufchan_r = (! lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_d = (lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf[0] ? lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf :
                                                          lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_r && lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf[0]))
        lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_main_mask_Bool3_1_argbuf_r) && (! lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf[0])))
        lizzieLet24_3Lcall_main_mask_Bool3_bufchan_buf <= lizzieLet24_3Lcall_main_mask_Bool3_bufchan_d;
  
  /* demux (Ty CTmain_mask_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet24_4,CTmain_mask_Bool) (srtarg_0_1_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet24_4Lmain_mask_Boolsbos,Pointer_QTree_Bool),
                                                                                                              (lizzieLet24_4Lcall_main_mask_Bool3,Pointer_QTree_Bool),
                                                                                                              (lizzieLet24_4Lcall_main_mask_Bool2,Pointer_QTree_Bool),
                                                                                                              (lizzieLet24_4Lcall_main_mask_Bool1,Pointer_QTree_Bool),
                                                                                                              (lizzieLet24_4Lcall_main_mask_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet24_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign lizzieLet24_4Lmain_mask_Boolsbos_d = {srtarg_0_1_goMux_mux_d[16:1],
                                               srtarg_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet24_4Lcall_main_mask_Bool3_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet24_4Lcall_main_mask_Bool2_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet24_4Lcall_main_mask_Bool1_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[3]};
  assign lizzieLet24_4Lcall_main_mask_Bool0_d = {srtarg_0_1_goMux_mux_d[16:1],
                                                 srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {lizzieLet24_4Lcall_main_mask_Bool0_r,
                                                                      lizzieLet24_4Lcall_main_mask_Bool1_r,
                                                                      lizzieLet24_4Lcall_main_mask_Bool2_r,
                                                                      lizzieLet24_4Lcall_main_mask_Bool3_r,
                                                                      lizzieLet24_4Lmain_mask_Boolsbos_r}));
  assign lizzieLet24_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet24_4Lcall_main_mask_Bool0,Pointer_QTree_Bool),
                          (es_1_destruct,Pointer_QTree_Bool),
                          (es_2_3_destruct,Pointer_QTree_Bool),
                          (es_3_4_destruct,Pointer_QTree_Bool)] > (lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool,QTree_Bool) */
  assign lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet24_4Lcall_main_mask_Bool0_d[0],
                                                                                                    es_1_destruct_d[0],
                                                                                                    es_2_3_destruct_d[0],
                                                                                                    es_3_4_destruct_d[0]}), lizzieLet24_4Lcall_main_mask_Bool0_d, es_1_destruct_d, es_2_3_destruct_d, es_3_4_destruct_d);
  assign {lizzieLet24_4Lcall_main_mask_Bool0_r,
          es_1_destruct_r,
          es_2_3_destruct_r,
          es_3_4_destruct_r} = {4 {(lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_r && lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool,QTree_Bool) > (lizzieLet28_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d;
  logic lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_r;
  assign lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_r = ((! lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d[0]) || lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                         1'd0};
    else
      if (lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_r)
        lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d <= lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_d;
  QTree_Bool_t lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf;
  assign lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_r = (! lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf[0] ? lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf :
                                   lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                           1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf[0]))
        lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                             1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf[0])))
        lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_buf <= lizzieLet24_4Lcall_main_mask_Bool0_1es_1_1es_2_3_1es_3_4_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool0) : [(lizzieLet24_4Lcall_main_mask_Bool1,Pointer_QTree_Bool),
                                     (es_2_2_destruct,Pointer_QTree_Bool),
                                     (es_3_3_destruct,Pointer_QTree_Bool),
                                     (sc_0_8_destruct,Pointer_CTmain_mask_Bool)] > (lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0,CTmain_mask_Bool) */
  assign lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_d = Lcall_main_mask_Bool0_dc((& {lizzieLet24_4Lcall_main_mask_Bool1_d[0],
                                                                                                                            es_2_2_destruct_d[0],
                                                                                                                            es_3_3_destruct_d[0],
                                                                                                                            sc_0_8_destruct_d[0]}), lizzieLet24_4Lcall_main_mask_Bool1_d, es_2_2_destruct_d, es_3_3_destruct_d, sc_0_8_destruct_d);
  assign {lizzieLet24_4Lcall_main_mask_Bool1_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r,
          sc_0_8_destruct_r} = {4 {(lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_r && lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0,CTmain_mask_Bool) > (lizzieLet27_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d;
  logic lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_r;
  assign lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_r = ((! lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d[0]) || lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d <= {115'd0,
                                                                                                      1'd0};
    else
      if (lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_r)
        lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d <= lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_d;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf;
  assign lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_r = (! lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf[0] ? lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf :
                                   lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf <= {115'd0,
                                                                                                        1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf[0]))
        lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf <= {115'd0,
                                                                                                          1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf[0])))
        lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_buf <= lizzieLet24_4Lcall_main_mask_Bool1_1es_2_2_1es_3_3_1sc_0_8_1Lcall_main_mask_Bool0_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool1) : [(lizzieLet24_4Lcall_main_mask_Bool2,Pointer_QTree_Bool),
                                     (es_3_2_destruct,Pointer_QTree_Bool),
                                     (sc_0_7_destruct,Pointer_CTmain_mask_Bool),
                                     (t1a8x_2_destruct,Pointer_QTree_Bool),
                                     (q1a8s_2_destruct,Pointer_MaskQTree)] > (lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1,CTmain_mask_Bool) */
  assign lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_d = Lcall_main_mask_Bool1_dc((& {lizzieLet24_4Lcall_main_mask_Bool2_d[0],
                                                                                                                                      es_3_2_destruct_d[0],
                                                                                                                                      sc_0_7_destruct_d[0],
                                                                                                                                      t1a8x_2_destruct_d[0],
                                                                                                                                      q1a8s_2_destruct_d[0]}), lizzieLet24_4Lcall_main_mask_Bool2_d, es_3_2_destruct_d, sc_0_7_destruct_d, t1a8x_2_destruct_d, q1a8s_2_destruct_d);
  assign {lizzieLet24_4Lcall_main_mask_Bool2_r,
          es_3_2_destruct_r,
          sc_0_7_destruct_r,
          t1a8x_2_destruct_r,
          q1a8s_2_destruct_r} = {5 {(lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_r && lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1,CTmain_mask_Bool) > (lizzieLet26_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d;
  logic lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_r;
  assign lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_r = ((! lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d[0]) || lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d <= {115'd0,
                                                                                                                1'd0};
    else
      if (lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_r)
        lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d <= lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_d;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf;
  assign lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_r = (! lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf[0] ? lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf :
                                   lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf <= {115'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf[0]))
        lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf <= {115'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf[0])))
        lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_buf <= lizzieLet24_4Lcall_main_mask_Bool2_1es_3_2_1sc_0_7_1t1a8x_2_1q1a8s_2_1Lcall_main_mask_Bool1_bufchan_d;
  
  /* dcon (Ty CTmain_mask_Bool,
      Dcon Lcall_main_mask_Bool2) : [(lizzieLet24_4Lcall_main_mask_Bool3,Pointer_QTree_Bool),
                                     (sc_0_6_destruct,Pointer_CTmain_mask_Bool),
                                     (t1a8x_1_destruct,Pointer_QTree_Bool),
                                     (q1a8s_1_destruct,Pointer_MaskQTree),
                                     (t2a8y_1_destruct,Pointer_QTree_Bool),
                                     (q2a8t_1_destruct,Pointer_MaskQTree)] > (lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2,CTmain_mask_Bool) */
  assign lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_d = Lcall_main_mask_Bool2_dc((& {lizzieLet24_4Lcall_main_mask_Bool3_d[0],
                                                                                                                                                sc_0_6_destruct_d[0],
                                                                                                                                                t1a8x_1_destruct_d[0],
                                                                                                                                                q1a8s_1_destruct_d[0],
                                                                                                                                                t2a8y_1_destruct_d[0],
                                                                                                                                                q2a8t_1_destruct_d[0]}), lizzieLet24_4Lcall_main_mask_Bool3_d, sc_0_6_destruct_d, t1a8x_1_destruct_d, q1a8s_1_destruct_d, t2a8y_1_destruct_d, q2a8t_1_destruct_d);
  assign {lizzieLet24_4Lcall_main_mask_Bool3_r,
          sc_0_6_destruct_r,
          t1a8x_1_destruct_r,
          q1a8s_1_destruct_r,
          t2a8y_1_destruct_r,
          q2a8t_1_destruct_r} = {6 {(lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_r && lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_d[0])}};
  
  /* buf (Ty CTmain_mask_Bool) : (lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2,CTmain_mask_Bool) > (lizzieLet25_1_argbuf,CTmain_mask_Bool) */
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d;
  logic lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_r;
  assign lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_r = ((! lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d[0]) || lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d <= {115'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_r)
        lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d <= lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_d;
  CTmain_mask_Bool_t lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf;
  assign lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_r = (! lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf[0] ? lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf :
                                   lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf <= {115'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf[0]))
        lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf <= {115'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf[0])))
        lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_buf <= lizzieLet24_4Lcall_main_mask_Bool3_1sc_0_6_1t1a8x_1_1q1a8s_1_1t2a8y_1_1q2a8t_1_1Lcall_main_mask_Bool2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lmain_mask_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                        (lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet24_4Lmain_mask_Boolsbos_emitted;
  logic [1:0] lizzieLet24_4Lmain_mask_Boolsbos_done;
  assign lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d = {lizzieLet24_4Lmain_mask_Boolsbos_d[16:1],
                                                                    (lizzieLet24_4Lmain_mask_Boolsbos_d[0] && (! lizzieLet24_4Lmain_mask_Boolsbos_emitted[0]))};
  assign lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d = {lizzieLet24_4Lmain_mask_Boolsbos_d[16:1],
                                                                    (lizzieLet24_4Lmain_mask_Boolsbos_d[0] && (! lizzieLet24_4Lmain_mask_Boolsbos_emitted[1]))};
  assign lizzieLet24_4Lmain_mask_Boolsbos_done = (lizzieLet24_4Lmain_mask_Boolsbos_emitted | ({lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d[0],
                                                                                               lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r,
                                                                                                                                                              lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet24_4Lmain_mask_Boolsbos_r = (& lizzieLet24_4Lmain_mask_Boolsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lmain_mask_Boolsbos_emitted <= 2'd0;
    else
      lizzieLet24_4Lmain_mask_Boolsbos_emitted <= (lizzieLet24_4Lmain_mask_Boolsbos_r ? 2'd0 :
                                                   lizzieLet24_4Lmain_mask_Boolsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_main_mask_Bool_goConst,Go) */
  assign call_main_mask_Bool_goConst_d = lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_1_r = call_main_mask_Bool_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (main_mask_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r = ((! lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                          1'd0};
    else
      if (lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_r)
        lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign main_mask_Bool_resbuf_d = (lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf :
                                    lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                            1'd0};
    else
      if ((main_mask_Bool_resbuf_r && lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                              1'd0};
      else if (((! main_mask_Bool_resbuf_r) && (! lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet24_4Lmain_mask_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (ma8q_1,Pointer_QTree_Bool) > (ma8q_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t ma8q_1_bufchan_d;
  logic ma8q_1_bufchan_r;
  assign ma8q_1_r = ((! ma8q_1_bufchan_d[0]) || ma8q_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_bufchan_d <= {16'd0, 1'd0};
    else if (ma8q_1_r) ma8q_1_bufchan_d <= ma8q_1_d;
  Pointer_QTree_Bool_t ma8q_1_bufchan_buf;
  assign ma8q_1_bufchan_r = (! ma8q_1_bufchan_buf[0]);
  assign ma8q_1_argbuf_d = (ma8q_1_bufchan_buf[0] ? ma8q_1_bufchan_buf :
                            ma8q_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((ma8q_1_argbuf_r && ma8q_1_bufchan_buf[0]))
        ma8q_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! ma8q_1_argbuf_r) && (! ma8q_1_bufchan_buf[0])))
        ma8q_1_bufchan_buf <= ma8q_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (ma8q_goMux_mux,Pointer_QTree_Bool) > [(ma8q_1,Pointer_QTree_Bool),
                                                                      (ma8q_2,Pointer_QTree_Bool)] */
  logic [1:0] ma8q_goMux_mux_emitted;
  logic [1:0] ma8q_goMux_mux_done;
  assign ma8q_1_d = {ma8q_goMux_mux_d[16:1],
                     (ma8q_goMux_mux_d[0] && (! ma8q_goMux_mux_emitted[0]))};
  assign ma8q_2_d = {ma8q_goMux_mux_d[16:1],
                     (ma8q_goMux_mux_d[0] && (! ma8q_goMux_mux_emitted[1]))};
  assign ma8q_goMux_mux_done = (ma8q_goMux_mux_emitted | ({ma8q_2_d[0],
                                                           ma8q_1_d[0]} & {ma8q_2_r, ma8q_1_r}));
  assign ma8q_goMux_mux_r = (& ma8q_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) ma8q_goMux_mux_emitted <= 2'd0;
    else
      ma8q_goMux_mux_emitted <= (ma8q_goMux_mux_r ? 2'd0 :
                                 ma8q_goMux_mux_done);
  
  /* destruct (Ty TupGo___Pointer_QTree_Bool___Pointer_MaskQTree,
          Dcon TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1,TupGo___Pointer_QTree_Bool___Pointer_MaskQTree) > [(main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6,Go),
                                                                                                                                                                                    (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1,Pointer_QTree_Bool),
                                                                                                                                                                                    (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1,Pointer_MaskQTree)] */
  logic [2:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted;
  logic [2:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[0]));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_d = {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[16:1],
                                                                                 (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[1]))};
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_d = {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[32:17],
                                                                                   (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted[2]))};
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted | ({main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_d[0],
                                                                                                                                                           main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_d[0],
                                                                                                                                                           main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_d[0]} & {main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_r,
                                                                                                                                                                                                                                     main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_r,
                                                                                                                                                                                                                                     main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_r}));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r = (& main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted <= 3'd0;
    else
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_emitted <= (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_r ? 3'd0 :
                                                                                 main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTree_1_done);
  
  /* fork (Ty Go) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6,Go) > [(go_6_1,Go),
                                                                                        (go_6_2,Go)] */
  logic [1:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted;
  logic [1:0] main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_done;
  assign go_6_1_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted[0]));
  assign go_6_2_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_d[0] && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted[1]));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_done = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted | ({go_6_2_d[0],
                                                                                                                                                               go_6_1_d[0]} & {go_6_2_r,
                                                                                                                                                                               go_6_1_r}));
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_r = (& main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted <= 2'd0;
    else
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_emitted <= (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_r ? 2'd0 :
                                                                                   main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreego_6_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1,Pointer_QTree_Bool) > (ma8q_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_r;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_r = ((! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d[0]) || main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d <= {16'd0,
                                                                                       1'd0};
    else
      if (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_r)
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_d;
  Pointer_QTree_Bool_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_r = (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf[0]);
  assign ma8q_1_1_argbuf_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf[0] ? main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf :
                              main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf <= {16'd0,
                                                                                         1'd0};
    else
      if ((ma8q_1_1_argbuf_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf[0]))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
      else if (((! ma8q_1_1_argbuf_r) && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf[0])))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_buf <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreema8q_1_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1,Pointer_MaskQTree) > (mska8r_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d;
  logic main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_r;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_r = ((! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d[0]) || main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d <= {16'd0,
                                                                                         1'd0};
    else
      if (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_r)
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_d;
  Pointer_MaskQTree_t main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf;
  assign main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_r = (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf[0]);
  assign mska8r_1_1_argbuf_d = (main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf[0] ? main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf :
                                main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf <= {16'd0,
                                                                                           1'd0};
    else
      if ((mska8r_1_1_argbuf_r && main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf[0]))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf <= {16'd0,
                                                                                             1'd0};
      else if (((! mska8r_1_1_argbuf_r) && (! main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf[0])))
        main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_buf <= main_mask_BoolTupGo___Pointer_QTree_Bool___Pointer_MaskQTreemska8r_1_bufchan_d;
  
  /* sink (Ty Pointer_QTree_Bool) : (main_mask_Bool_resbuf,Pointer_QTree_Bool) > */
  assign {main_mask_Bool_resbuf_r,
          main_mask_Bool_resbuf_dout} = {main_mask_Bool_resbuf_rout,
                                         main_mask_Bool_resbuf_d};
  
  /* buf (Ty Pointer_MaskQTree) : (mska8r_goMux_mux,Pointer_MaskQTree) > (mska8r_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t mska8r_goMux_mux_bufchan_d;
  logic mska8r_goMux_mux_bufchan_r;
  assign mska8r_goMux_mux_r = ((! mska8r_goMux_mux_bufchan_d[0]) || mska8r_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mska8r_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (mska8r_goMux_mux_r)
        mska8r_goMux_mux_bufchan_d <= mska8r_goMux_mux_d;
  Pointer_MaskQTree_t mska8r_goMux_mux_bufchan_buf;
  assign mska8r_goMux_mux_bufchan_r = (! mska8r_goMux_mux_bufchan_buf[0]);
  assign mska8r_1_argbuf_d = (mska8r_goMux_mux_bufchan_buf[0] ? mska8r_goMux_mux_bufchan_buf :
                              mska8r_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mska8r_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mska8r_1_argbuf_r && mska8r_goMux_mux_bufchan_buf[0]))
        mska8r_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mska8r_1_argbuf_r) && (! mska8r_goMux_mux_bufchan_buf[0])))
        mska8r_goMux_mux_bufchan_buf <= mska8r_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1a8h_3_destruct,Pointer_QTree_Bool) > (q1a8h_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1a8h_3_destruct_bufchan_d;
  logic q1a8h_3_destruct_bufchan_r;
  assign q1a8h_3_destruct_r = ((! q1a8h_3_destruct_bufchan_d[0]) || q1a8h_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8h_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8h_3_destruct_r)
        q1a8h_3_destruct_bufchan_d <= q1a8h_3_destruct_d;
  Pointer_QTree_Bool_t q1a8h_3_destruct_bufchan_buf;
  assign q1a8h_3_destruct_bufchan_r = (! q1a8h_3_destruct_bufchan_buf[0]);
  assign q1a8h_3_1_argbuf_d = (q1a8h_3_destruct_bufchan_buf[0] ? q1a8h_3_destruct_bufchan_buf :
                               q1a8h_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8h_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8h_3_1_argbuf_r && q1a8h_3_destruct_bufchan_buf[0]))
        q1a8h_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8h_3_1_argbuf_r) && (! q1a8h_3_destruct_bufchan_buf[0])))
        q1a8h_3_destruct_bufchan_buf <= q1a8h_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q1a8s_3_destruct,Pointer_MaskQTree) > (q1a8s_3_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q1a8s_3_destruct_bufchan_d;
  logic q1a8s_3_destruct_bufchan_r;
  assign q1a8s_3_destruct_r = ((! q1a8s_3_destruct_bufchan_d[0]) || q1a8s_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8s_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1a8s_3_destruct_r)
        q1a8s_3_destruct_bufchan_d <= q1a8s_3_destruct_d;
  Pointer_MaskQTree_t q1a8s_3_destruct_bufchan_buf;
  assign q1a8s_3_destruct_bufchan_r = (! q1a8s_3_destruct_bufchan_buf[0]);
  assign q1a8s_3_1_argbuf_d = (q1a8s_3_destruct_bufchan_buf[0] ? q1a8s_3_destruct_bufchan_buf :
                               q1a8s_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1a8s_3_1_argbuf_r && q1a8s_3_destruct_bufchan_buf[0]))
        q1a8s_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1a8s_3_1_argbuf_r) && (! q1a8s_3_destruct_bufchan_buf[0])))
        q1a8s_3_destruct_bufchan_buf <= q1a8s_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2a8i_2_destruct,Pointer_QTree_Bool) > (q2a8i_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2a8i_2_destruct_bufchan_d;
  logic q2a8i_2_destruct_bufchan_r;
  assign q2a8i_2_destruct_r = ((! q2a8i_2_destruct_bufchan_d[0]) || q2a8i_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8i_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8i_2_destruct_r)
        q2a8i_2_destruct_bufchan_d <= q2a8i_2_destruct_d;
  Pointer_QTree_Bool_t q2a8i_2_destruct_bufchan_buf;
  assign q2a8i_2_destruct_bufchan_r = (! q2a8i_2_destruct_bufchan_buf[0]);
  assign q2a8i_2_1_argbuf_d = (q2a8i_2_destruct_bufchan_buf[0] ? q2a8i_2_destruct_bufchan_buf :
                               q2a8i_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8i_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8i_2_1_argbuf_r && q2a8i_2_destruct_bufchan_buf[0]))
        q2a8i_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8i_2_1_argbuf_r) && (! q2a8i_2_destruct_bufchan_buf[0])))
        q2a8i_2_destruct_bufchan_buf <= q2a8i_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q2a8t_2_destruct,Pointer_MaskQTree) > (q2a8t_2_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q2a8t_2_destruct_bufchan_d;
  logic q2a8t_2_destruct_bufchan_r;
  assign q2a8t_2_destruct_r = ((! q2a8t_2_destruct_bufchan_d[0]) || q2a8t_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8t_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2a8t_2_destruct_r)
        q2a8t_2_destruct_bufchan_d <= q2a8t_2_destruct_d;
  Pointer_MaskQTree_t q2a8t_2_destruct_bufchan_buf;
  assign q2a8t_2_destruct_bufchan_r = (! q2a8t_2_destruct_bufchan_buf[0]);
  assign q2a8t_2_1_argbuf_d = (q2a8t_2_destruct_bufchan_buf[0] ? q2a8t_2_destruct_bufchan_buf :
                               q2a8t_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2a8t_2_1_argbuf_r && q2a8t_2_destruct_bufchan_buf[0]))
        q2a8t_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2a8t_2_1_argbuf_r) && (! q2a8t_2_destruct_bufchan_buf[0])))
        q2a8t_2_destruct_bufchan_buf <= q2a8t_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3a8j_1_destruct,Pointer_QTree_Bool) > (q3a8j_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3a8j_1_destruct_bufchan_d;
  logic q3a8j_1_destruct_bufchan_r;
  assign q3a8j_1_destruct_r = ((! q3a8j_1_destruct_bufchan_d[0]) || q3a8j_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8j_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8j_1_destruct_r)
        q3a8j_1_destruct_bufchan_d <= q3a8j_1_destruct_d;
  Pointer_QTree_Bool_t q3a8j_1_destruct_bufchan_buf;
  assign q3a8j_1_destruct_bufchan_r = (! q3a8j_1_destruct_bufchan_buf[0]);
  assign q3a8j_1_1_argbuf_d = (q3a8j_1_destruct_bufchan_buf[0] ? q3a8j_1_destruct_bufchan_buf :
                               q3a8j_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8j_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8j_1_1_argbuf_r && q3a8j_1_destruct_bufchan_buf[0]))
        q3a8j_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8j_1_1_argbuf_r) && (! q3a8j_1_destruct_bufchan_buf[0])))
        q3a8j_1_destruct_bufchan_buf <= q3a8j_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_MaskQTree) : (q3a8u_1_destruct,Pointer_MaskQTree) > (q3a8u_1_1_argbuf,Pointer_MaskQTree) */
  Pointer_MaskQTree_t q3a8u_1_destruct_bufchan_d;
  logic q3a8u_1_destruct_bufchan_r;
  assign q3a8u_1_destruct_r = ((! q3a8u_1_destruct_bufchan_d[0]) || q3a8u_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8u_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3a8u_1_destruct_r)
        q3a8u_1_destruct_bufchan_d <= q3a8u_1_destruct_d;
  Pointer_MaskQTree_t q3a8u_1_destruct_bufchan_buf;
  assign q3a8u_1_destruct_bufchan_r = (! q3a8u_1_destruct_bufchan_buf[0]);
  assign q3a8u_1_1_argbuf_d = (q3a8u_1_destruct_bufchan_buf[0] ? q3a8u_1_destruct_bufchan_buf :
                               q3a8u_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3a8u_1_1_argbuf_r && q3a8u_1_destruct_bufchan_buf[0]))
        q3a8u_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3a8u_1_1_argbuf_r) && (! q3a8u_1_destruct_bufchan_buf[0])))
        q3a8u_1_destruct_bufchan_buf <= q3a8u_1_destruct_bufchan_d;
  
  /* buf (Ty CT$wmAdd_Bool) : (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf,CT$wmAdd_Bool) > (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb,CT$wmAdd_Bool) */
  CT$wmAdd_Bool_t readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_r = ((! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                               1'd0};
    else
      if (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_r)
        readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_d;
  CT$wmAdd_Bool_t readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf :
                                                             readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
    else
      if ((readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_r && readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                   1'd0};
      else if (((! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wmAdd_Bool) : (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb,CT$wmAdd_Bool) > [(lizzieLet19_1,CT$wmAdd_Bool),
                                                                                            (lizzieLet19_2,CT$wmAdd_Bool),
                                                                                            (lizzieLet19_3,CT$wmAdd_Bool),
                                                                                            (lizzieLet19_4,CT$wmAdd_Bool)] */
  logic [3:0] readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet19_1_d = {readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet19_2_d = {readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet19_3_d = {readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet19_4_d = {readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet19_4_d[0],
                                                                                                                           lizzieLet19_3_d[0],
                                                                                                                           lizzieLet19_2_d[0],
                                                                                                                           lizzieLet19_1_d[0]} & {lizzieLet19_4_r,
                                                                                                                                                  lizzieLet19_3_r,
                                                                                                                                                  lizzieLet19_2_r,
                                                                                                                                                  lizzieLet19_1_r}));
  assign readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                                 readPointer_CT$wmAdd_Boolscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_mask_Bool) : (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf,CTmain_mask_Bool) > (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb,CTmain_mask_Bool) */
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d;
  logic readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r;
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r = ((! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d[0]) || readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d <= {115'd0,
                                                                    1'd0};
    else
      if (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_r)
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d <= readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_d;
  CTmain_mask_Bool_t readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf;
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_r = (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d = (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0] ? readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf :
                                                                  readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                      1'd0};
    else
      if ((readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r && readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0]))
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= {115'd0,
                                                                        1'd0};
      else if (((! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r) && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf[0])))
        readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_buf <= readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_bufchan_d;
  
  /* fork (Ty CTmain_mask_Bool) : (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb,CTmain_mask_Bool) > [(lizzieLet24_1,CTmain_mask_Bool),
                                                                                                       (lizzieLet24_2,CTmain_mask_Bool),
                                                                                                       (lizzieLet24_3,CTmain_mask_Bool),
                                                                                                       (lizzieLet24_4,CTmain_mask_Bool)] */
  logic [3:0] readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done;
  assign lizzieLet24_1_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet24_2_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet24_3_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet24_4_d = {readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[115:1],
                            (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_d[0] && (! readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done = (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted | ({lizzieLet24_4_d[0],
                                                                                                                                     lizzieLet24_3_d[0],
                                                                                                                                     lizzieLet24_2_d[0],
                                                                                                                                     lizzieLet24_1_d[0]} & {lizzieLet24_4_r,
                                                                                                                                                            lizzieLet24_3_r,
                                                                                                                                                            lizzieLet24_2_r,
                                                                                                                                                            lizzieLet24_1_r}));
  assign readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r = (& readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_emitted <= (readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_r ? 4'd0 :
                                                                      readPointer_CTmain_mask_Boolscfarg_0_1_1_argbuf_rwb_done);
  
  /* buf (Ty MaskQTree) : (readPointer_MaskQTreemska8r_1_argbuf,MaskQTree) > (readPointer_MaskQTreemska8r_1_argbuf_rwb,MaskQTree) */
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_bufchan_d;
  logic readPointer_MaskQTreemska8r_1_argbuf_bufchan_r;
  assign readPointer_MaskQTreemska8r_1_argbuf_r = ((! readPointer_MaskQTreemska8r_1_argbuf_bufchan_d[0]) || readPointer_MaskQTreemska8r_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_MaskQTreemska8r_1_argbuf_r)
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_d <= readPointer_MaskQTreemska8r_1_argbuf_d;
  MaskQTree_t readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf;
  assign readPointer_MaskQTreemska8r_1_argbuf_bufchan_r = (! readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0]);
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_d = (readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0] ? readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf :
                                                       readPointer_MaskQTreemska8r_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_MaskQTreemska8r_1_argbuf_rwb_r && readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0]))
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_MaskQTreemska8r_1_argbuf_rwb_r) && (! readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf[0])))
        readPointer_MaskQTreemska8r_1_argbuf_bufchan_buf <= readPointer_MaskQTreemska8r_1_argbuf_bufchan_d;
  
  /* fork (Ty MaskQTree) : (readPointer_MaskQTreemska8r_1_argbuf_rwb,MaskQTree) > [(lizzieLet11_1_1,MaskQTree),
                                                                              (lizzieLet11_1_2,MaskQTree),
                                                                              (lizzieLet11_1_3,MaskQTree),
                                                                              (lizzieLet11_1_4,MaskQTree),
                                                                              (lizzieLet11_1_5,MaskQTree),
                                                                              (lizzieLet11_1_6,MaskQTree)] */
  logic [5:0] readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_MaskQTreemska8r_1_argbuf_rwb_done;
  assign lizzieLet11_1_1_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet11_1_2_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet11_1_3_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet11_1_4_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet11_1_5_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet11_1_6_d = {readPointer_MaskQTreemska8r_1_argbuf_rwb_d[66:1],
                              (readPointer_MaskQTreemska8r_1_argbuf_rwb_d[0] && (! readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted[5]))};
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_done = (readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted | ({lizzieLet11_1_6_d[0],
                                                                                                               lizzieLet11_1_5_d[0],
                                                                                                               lizzieLet11_1_4_d[0],
                                                                                                               lizzieLet11_1_3_d[0],
                                                                                                               lizzieLet11_1_2_d[0],
                                                                                                               lizzieLet11_1_1_d[0]} & {lizzieLet11_1_6_r,
                                                                                                                                        lizzieLet11_1_5_r,
                                                                                                                                        lizzieLet11_1_4_r,
                                                                                                                                        lizzieLet11_1_3_r,
                                                                                                                                        lizzieLet11_1_2_r,
                                                                                                                                        lizzieLet11_1_1_r}));
  assign readPointer_MaskQTreemska8r_1_argbuf_rwb_r = (& readPointer_MaskQTreemska8r_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_MaskQTreemska8r_1_argbuf_rwb_emitted <= (readPointer_MaskQTreemska8r_1_argbuf_rwb_r ? 6'd0 :
                                                           readPointer_MaskQTreemska8r_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolma8q_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolma8q_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolma8q_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolma8q_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolma8q_1_argbuf_r = ((! readPointer_QTree_Boolma8q_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolma8q_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolma8q_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolma8q_1_argbuf_r)
        readPointer_QTree_Boolma8q_1_argbuf_bufchan_d <= readPointer_QTree_Boolma8q_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolma8q_1_argbuf_bufchan_r = (! readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolma8q_1_argbuf_rwb_d = (readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Boolma8q_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolma8q_1_argbuf_rwb_r && readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolma8q_1_argbuf_rwb_r) && (! readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolma8q_1_argbuf_bufchan_buf <= readPointer_QTree_Boolma8q_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolw1sic_1_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_r = ((! readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolw1sic_1_1_argbuf_r)
        readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d <= readPointer_QTree_Boolw1sic_1_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_r = (! readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d = (readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf :
                                                         readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf <= {66'd0,
                                                             1'd0};
    else
      if ((readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_r && readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf <= {66'd0,
                                                               1'd0};
      else if (((! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_r) && (! readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_buf <= readPointer_QTree_Boolw1sic_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb,QTree_Bool) > [(lizzieLet1_1,QTree_Bool),
                                                                                  (lizzieLet1_2,QTree_Bool),
                                                                                  (lizzieLet1_3,QTree_Bool),
                                                                                  (lizzieLet1_4,QTree_Bool),
                                                                                  (lizzieLet1_5,QTree_Bool),
                                                                                  (lizzieLet1_6,QTree_Bool),
                                                                                  (lizzieLet1_7,QTree_Bool),
                                                                                  (lizzieLet1_8,QTree_Bool)] */
  logic [7:0] readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted;
  logic [7:0] readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_done;
  assign lizzieLet1_1_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet1_2_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet1_3_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet1_4_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet1_5_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet1_6_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet1_7_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet1_8_d = {readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted[7]))};
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_done = (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted | ({lizzieLet1_8_d[0],
                                                                                                                   lizzieLet1_7_d[0],
                                                                                                                   lizzieLet1_6_d[0],
                                                                                                                   lizzieLet1_5_d[0],
                                                                                                                   lizzieLet1_4_d[0],
                                                                                                                   lizzieLet1_3_d[0],
                                                                                                                   lizzieLet1_2_d[0],
                                                                                                                   lizzieLet1_1_d[0]} & {lizzieLet1_8_r,
                                                                                                                                         lizzieLet1_7_r,
                                                                                                                                         lizzieLet1_6_r,
                                                                                                                                         lizzieLet1_5_r,
                                                                                                                                         lizzieLet1_4_r,
                                                                                                                                         lizzieLet1_3_r,
                                                                                                                                         lizzieLet1_2_r,
                                                                                                                                         lizzieLet1_1_r}));
  assign readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_r = (& readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted <= 8'd0;
    else
      readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_r ? 8'd0 :
                                                             readPointer_QTree_Boolw1sic_1_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolw2sid_1_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolw2sid_1_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolw2sid_1_1_argbuf_r = ((! readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolw2sid_1_1_argbuf_r)
        readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d <= readPointer_QTree_Boolw2sid_1_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_r = (! readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_d = (readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf :
                                                         readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf <= {66'd0,
                                                             1'd0};
    else
      if ((readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_r && readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf <= {66'd0,
                                                               1'd0};
      else if (((! readPointer_QTree_Boolw2sid_1_1_argbuf_rwb_r) && (! readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_buf <= readPointer_QTree_Boolw2sid_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (sc_0_5_destruct,Pointer_CT$wmAdd_Bool) > (sc_0_5_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t sc_0_5_destruct_bufchan_d;
  logic sc_0_5_destruct_bufchan_r;
  assign sc_0_5_destruct_r = ((! sc_0_5_destruct_bufchan_d[0]) || sc_0_5_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_5_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_5_destruct_r)
        sc_0_5_destruct_bufchan_d <= sc_0_5_destruct_d;
  Pointer_CT$wmAdd_Bool_t sc_0_5_destruct_bufchan_buf;
  assign sc_0_5_destruct_bufchan_r = (! sc_0_5_destruct_bufchan_buf[0]);
  assign sc_0_5_1_argbuf_d = (sc_0_5_destruct_bufchan_buf[0] ? sc_0_5_destruct_bufchan_buf :
                              sc_0_5_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_5_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_5_1_argbuf_r && sc_0_5_destruct_bufchan_buf[0]))
        sc_0_5_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_5_1_argbuf_r) && (! sc_0_5_destruct_bufchan_buf[0])))
        sc_0_5_destruct_bufchan_buf <= sc_0_5_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (sc_0_9_destruct,Pointer_CTmain_mask_Bool) > (sc_0_9_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t sc_0_9_destruct_bufchan_d;
  logic sc_0_9_destruct_bufchan_r;
  assign sc_0_9_destruct_r = ((! sc_0_9_destruct_bufchan_d[0]) || sc_0_9_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_9_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_9_destruct_r)
        sc_0_9_destruct_bufchan_d <= sc_0_9_destruct_d;
  Pointer_CTmain_mask_Bool_t sc_0_9_destruct_bufchan_buf;
  assign sc_0_9_destruct_bufchan_r = (! sc_0_9_destruct_bufchan_buf[0]);
  assign sc_0_9_1_argbuf_d = (sc_0_9_destruct_bufchan_buf[0] ? sc_0_9_destruct_bufchan_buf :
                              sc_0_9_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_9_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_9_1_argbuf_r && sc_0_9_destruct_bufchan_buf[0]))
        sc_0_9_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_9_1_argbuf_r) && (! sc_0_9_destruct_bufchan_buf[0])))
        sc_0_9_destruct_bufchan_buf <= sc_0_9_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (scfarg_0_1_goMux_mux,Pointer_CTmain_mask_Bool) > (scfarg_0_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  Pointer_CTmain_mask_Bool_t scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (scfarg_0_goMux_mux,Pointer_CT$wmAdd_Bool) > (scfarg_0_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wmAdd_Bool_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8m_3_destruct,Pointer_QTree_Bool) > (t1a8m_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8m_3_destruct_bufchan_d;
  logic t1a8m_3_destruct_bufchan_r;
  assign t1a8m_3_destruct_r = ((! t1a8m_3_destruct_bufchan_d[0]) || t1a8m_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8m_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8m_3_destruct_r)
        t1a8m_3_destruct_bufchan_d <= t1a8m_3_destruct_d;
  Pointer_QTree_Bool_t t1a8m_3_destruct_bufchan_buf;
  assign t1a8m_3_destruct_bufchan_r = (! t1a8m_3_destruct_bufchan_buf[0]);
  assign t1a8m_3_1_argbuf_d = (t1a8m_3_destruct_bufchan_buf[0] ? t1a8m_3_destruct_bufchan_buf :
                               t1a8m_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8m_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8m_3_1_argbuf_r && t1a8m_3_destruct_bufchan_buf[0]))
        t1a8m_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8m_3_1_argbuf_r) && (! t1a8m_3_destruct_bufchan_buf[0])))
        t1a8m_3_destruct_bufchan_buf <= t1a8m_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t1a8x_3_destruct,Pointer_QTree_Bool) > (t1a8x_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t1a8x_3_destruct_bufchan_d;
  logic t1a8x_3_destruct_bufchan_r;
  assign t1a8x_3_destruct_r = ((! t1a8x_3_destruct_bufchan_d[0]) || t1a8x_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8x_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t1a8x_3_destruct_r)
        t1a8x_3_destruct_bufchan_d <= t1a8x_3_destruct_d;
  Pointer_QTree_Bool_t t1a8x_3_destruct_bufchan_buf;
  assign t1a8x_3_destruct_bufchan_r = (! t1a8x_3_destruct_bufchan_buf[0]);
  assign t1a8x_3_1_argbuf_d = (t1a8x_3_destruct_bufchan_buf[0] ? t1a8x_3_destruct_bufchan_buf :
                               t1a8x_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t1a8x_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t1a8x_3_1_argbuf_r && t1a8x_3_destruct_bufchan_buf[0]))
        t1a8x_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t1a8x_3_1_argbuf_r) && (! t1a8x_3_destruct_bufchan_buf[0])))
        t1a8x_3_destruct_bufchan_buf <= t1a8x_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8n_2_destruct,Pointer_QTree_Bool) > (t2a8n_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8n_2_destruct_bufchan_d;
  logic t2a8n_2_destruct_bufchan_r;
  assign t2a8n_2_destruct_r = ((! t2a8n_2_destruct_bufchan_d[0]) || t2a8n_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8n_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8n_2_destruct_r)
        t2a8n_2_destruct_bufchan_d <= t2a8n_2_destruct_d;
  Pointer_QTree_Bool_t t2a8n_2_destruct_bufchan_buf;
  assign t2a8n_2_destruct_bufchan_r = (! t2a8n_2_destruct_bufchan_buf[0]);
  assign t2a8n_2_1_argbuf_d = (t2a8n_2_destruct_bufchan_buf[0] ? t2a8n_2_destruct_bufchan_buf :
                               t2a8n_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8n_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8n_2_1_argbuf_r && t2a8n_2_destruct_bufchan_buf[0]))
        t2a8n_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8n_2_1_argbuf_r) && (! t2a8n_2_destruct_bufchan_buf[0])))
        t2a8n_2_destruct_bufchan_buf <= t2a8n_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t2a8y_2_destruct,Pointer_QTree_Bool) > (t2a8y_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t2a8y_2_destruct_bufchan_d;
  logic t2a8y_2_destruct_bufchan_r;
  assign t2a8y_2_destruct_r = ((! t2a8y_2_destruct_bufchan_d[0]) || t2a8y_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8y_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t2a8y_2_destruct_r)
        t2a8y_2_destruct_bufchan_d <= t2a8y_2_destruct_d;
  Pointer_QTree_Bool_t t2a8y_2_destruct_bufchan_buf;
  assign t2a8y_2_destruct_bufchan_r = (! t2a8y_2_destruct_bufchan_buf[0]);
  assign t2a8y_2_1_argbuf_d = (t2a8y_2_destruct_bufchan_buf[0] ? t2a8y_2_destruct_bufchan_buf :
                               t2a8y_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t2a8y_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t2a8y_2_1_argbuf_r && t2a8y_2_destruct_bufchan_buf[0]))
        t2a8y_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t2a8y_2_1_argbuf_r) && (! t2a8y_2_destruct_bufchan_buf[0])))
        t2a8y_2_destruct_bufchan_buf <= t2a8y_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8o_1_destruct,Pointer_QTree_Bool) > (t3a8o_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8o_1_destruct_bufchan_d;
  logic t3a8o_1_destruct_bufchan_r;
  assign t3a8o_1_destruct_r = ((! t3a8o_1_destruct_bufchan_d[0]) || t3a8o_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8o_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8o_1_destruct_r)
        t3a8o_1_destruct_bufchan_d <= t3a8o_1_destruct_d;
  Pointer_QTree_Bool_t t3a8o_1_destruct_bufchan_buf;
  assign t3a8o_1_destruct_bufchan_r = (! t3a8o_1_destruct_bufchan_buf[0]);
  assign t3a8o_1_1_argbuf_d = (t3a8o_1_destruct_bufchan_buf[0] ? t3a8o_1_destruct_bufchan_buf :
                               t3a8o_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8o_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8o_1_1_argbuf_r && t3a8o_1_destruct_bufchan_buf[0]))
        t3a8o_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8o_1_1_argbuf_r) && (! t3a8o_1_destruct_bufchan_buf[0])))
        t3a8o_1_destruct_bufchan_buf <= t3a8o_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t3a8z_1_destruct,Pointer_QTree_Bool) > (t3a8z_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t3a8z_1_destruct_bufchan_d;
  logic t3a8z_1_destruct_bufchan_r;
  assign t3a8z_1_destruct_r = ((! t3a8z_1_destruct_bufchan_d[0]) || t3a8z_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8z_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t3a8z_1_destruct_r)
        t3a8z_1_destruct_bufchan_d <= t3a8z_1_destruct_d;
  Pointer_QTree_Bool_t t3a8z_1_destruct_bufchan_buf;
  assign t3a8z_1_destruct_bufchan_r = (! t3a8z_1_destruct_bufchan_buf[0]);
  assign t3a8z_1_1_argbuf_d = (t3a8z_1_destruct_bufchan_buf[0] ? t3a8z_1_destruct_bufchan_buf :
                               t3a8z_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t3a8z_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t3a8z_1_1_argbuf_r && t3a8z_1_destruct_bufchan_buf[0]))
        t3a8z_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t3a8z_1_1_argbuf_r) && (! t3a8z_1_destruct_bufchan_buf[0])))
        t3a8z_1_destruct_bufchan_buf <= t3a8z_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8A_destruct,Pointer_QTree_Bool) > (t4a8A_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8A_destruct_bufchan_d;
  logic t4a8A_destruct_bufchan_r;
  assign t4a8A_destruct_r = ((! t4a8A_destruct_bufchan_d[0]) || t4a8A_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8A_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8A_destruct_r) t4a8A_destruct_bufchan_d <= t4a8A_destruct_d;
  Pointer_QTree_Bool_t t4a8A_destruct_bufchan_buf;
  assign t4a8A_destruct_bufchan_r = (! t4a8A_destruct_bufchan_buf[0]);
  assign t4a8A_1_argbuf_d = (t4a8A_destruct_bufchan_buf[0] ? t4a8A_destruct_bufchan_buf :
                             t4a8A_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8A_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8A_1_argbuf_r && t4a8A_destruct_bufchan_buf[0]))
        t4a8A_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8A_1_argbuf_r) && (! t4a8A_destruct_bufchan_buf[0])))
        t4a8A_destruct_bufchan_buf <= t4a8A_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (t4a8p_destruct,Pointer_QTree_Bool) > (t4a8p_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t t4a8p_destruct_bufchan_d;
  logic t4a8p_destruct_bufchan_r;
  assign t4a8p_destruct_r = ((! t4a8p_destruct_bufchan_d[0]) || t4a8p_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8p_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (t4a8p_destruct_r) t4a8p_destruct_bufchan_d <= t4a8p_destruct_d;
  Pointer_QTree_Bool_t t4a8p_destruct_bufchan_buf;
  assign t4a8p_destruct_bufchan_r = (! t4a8p_destruct_bufchan_buf[0]);
  assign t4a8p_1_argbuf_d = (t4a8p_destruct_bufchan_buf[0] ? t4a8p_destruct_bufchan_buf :
                             t4a8p_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) t4a8p_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((t4a8p_1_argbuf_r && t4a8p_destruct_bufchan_buf[0]))
        t4a8p_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! t4a8p_1_argbuf_r) && (! t4a8p_destruct_bufchan_buf[0])))
        t4a8p_destruct_bufchan_buf <= t4a8p_destruct_bufchan_d;
  
  /* buf (Ty MyBool) : (va8c_destruct,MyBool) > (va8c_1_argbuf,MyBool) */
  MyBool_t va8c_destruct_bufchan_d;
  logic va8c_destruct_bufchan_r;
  assign va8c_destruct_r = ((! va8c_destruct_bufchan_d[0]) || va8c_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8c_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (va8c_destruct_r) va8c_destruct_bufchan_d <= va8c_destruct_d;
  MyBool_t va8c_destruct_bufchan_buf;
  assign va8c_destruct_bufchan_r = (! va8c_destruct_bufchan_buf[0]);
  assign va8c_1_argbuf_d = (va8c_destruct_bufchan_buf[0] ? va8c_destruct_bufchan_buf :
                            va8c_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) va8c_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((va8c_1_argbuf_r && va8c_destruct_bufchan_buf[0]))
        va8c_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! va8c_1_argbuf_r) && (! va8c_destruct_bufchan_buf[0])))
        va8c_destruct_bufchan_buf <= va8c_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (w1sic_1_1,Pointer_QTree_Bool) > (w1sic_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t w1sic_1_1_bufchan_d;
  logic w1sic_1_1_bufchan_r;
  assign w1sic_1_1_r = ((! w1sic_1_1_bufchan_d[0]) || w1sic_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sic_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w1sic_1_1_r) w1sic_1_1_bufchan_d <= w1sic_1_1_d;
  Pointer_QTree_Bool_t w1sic_1_1_bufchan_buf;
  assign w1sic_1_1_bufchan_r = (! w1sic_1_1_bufchan_buf[0]);
  assign w1sic_1_1_argbuf_d = (w1sic_1_1_bufchan_buf[0] ? w1sic_1_1_bufchan_buf :
                               w1sic_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sic_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w1sic_1_1_argbuf_r && w1sic_1_1_bufchan_buf[0]))
        w1sic_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w1sic_1_1_argbuf_r) && (! w1sic_1_1_bufchan_buf[0])))
        w1sic_1_1_bufchan_buf <= w1sic_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (w1sic_1_goMux_mux,Pointer_QTree_Bool) > [(w1sic_1_1,Pointer_QTree_Bool),
                                                                         (w1sic_1_2,Pointer_QTree_Bool)] */
  logic [1:0] w1sic_1_goMux_mux_emitted;
  logic [1:0] w1sic_1_goMux_mux_done;
  assign w1sic_1_1_d = {w1sic_1_goMux_mux_d[16:1],
                        (w1sic_1_goMux_mux_d[0] && (! w1sic_1_goMux_mux_emitted[0]))};
  assign w1sic_1_2_d = {w1sic_1_goMux_mux_d[16:1],
                        (w1sic_1_goMux_mux_d[0] && (! w1sic_1_goMux_mux_emitted[1]))};
  assign w1sic_1_goMux_mux_done = (w1sic_1_goMux_mux_emitted | ({w1sic_1_2_d[0],
                                                                 w1sic_1_1_d[0]} & {w1sic_1_2_r,
                                                                                    w1sic_1_1_r}));
  assign w1sic_1_goMux_mux_r = (& w1sic_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w1sic_1_goMux_mux_emitted <= 2'd0;
    else
      w1sic_1_goMux_mux_emitted <= (w1sic_1_goMux_mux_r ? 2'd0 :
                                    w1sic_1_goMux_mux_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (w2sid_1_1,Pointer_QTree_Bool) > (w2sid_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t w2sid_1_1_bufchan_d;
  logic w2sid_1_1_bufchan_r;
  assign w2sid_1_1_r = ((! w2sid_1_1_bufchan_d[0]) || w2sid_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sid_1_1_bufchan_d <= {16'd0, 1'd0};
    else if (w2sid_1_1_r) w2sid_1_1_bufchan_d <= w2sid_1_1_d;
  Pointer_QTree_Bool_t w2sid_1_1_bufchan_buf;
  assign w2sid_1_1_bufchan_r = (! w2sid_1_1_bufchan_buf[0]);
  assign w2sid_1_1_argbuf_d = (w2sid_1_1_bufchan_buf[0] ? w2sid_1_1_bufchan_buf :
                               w2sid_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sid_1_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((w2sid_1_1_argbuf_r && w2sid_1_1_bufchan_buf[0]))
        w2sid_1_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! w2sid_1_1_argbuf_r) && (! w2sid_1_1_bufchan_buf[0])))
        w2sid_1_1_bufchan_buf <= w2sid_1_1_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (w2sid_1_goMux_mux,Pointer_QTree_Bool) > [(w2sid_1_1,Pointer_QTree_Bool),
                                                                         (w2sid_1_2,Pointer_QTree_Bool)] */
  logic [1:0] w2sid_1_goMux_mux_emitted;
  logic [1:0] w2sid_1_goMux_mux_done;
  assign w2sid_1_1_d = {w2sid_1_goMux_mux_d[16:1],
                        (w2sid_1_goMux_mux_d[0] && (! w2sid_1_goMux_mux_emitted[0]))};
  assign w2sid_1_2_d = {w2sid_1_goMux_mux_d[16:1],
                        (w2sid_1_goMux_mux_d[0] && (! w2sid_1_goMux_mux_emitted[1]))};
  assign w2sid_1_goMux_mux_done = (w2sid_1_goMux_mux_emitted | ({w2sid_1_2_d[0],
                                                                 w2sid_1_1_d[0]} & {w2sid_1_2_r,
                                                                                    w2sid_1_1_r}));
  assign w2sid_1_goMux_mux_r = (& w2sid_1_goMux_mux_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) w2sid_1_goMux_mux_emitted <= 2'd0;
    else
      w2sid_1_goMux_mux_emitted <= (w2sid_1_goMux_mux_r ? 2'd0 :
                                    w2sid_1_goMux_mux_done);
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet0_1_argbuf,Pointer_CT$wmAdd_Bool) > (writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_r = ((! writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet0_1_argbuf_r)
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d <= writeCT$wmAdd_BoollizzieLet0_1_argbuf_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_r = (! writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_d = (writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf :
                                                        writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_r && writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_r) && (! writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_buf <= writeCT$wmAdd_BoollizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) > (lizzieLet11_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_r = ((! writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_r)
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_BoollizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet20_1_argbuf,Pointer_CT$wmAdd_Bool) > (writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_r = ((! writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet20_1_argbuf_r)
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d <= writeCT$wmAdd_BoollizzieLet20_1_argbuf_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_r = (! writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_d = (writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf :
                                                         writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_r && writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_r) && (! writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_buf <= writeCT$wmAdd_BoollizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) > (sca2_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_r = ((! writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_r)
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_BoollizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet21_1_argbuf,Pointer_CT$wmAdd_Bool) > (writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_r = ((! writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet21_1_argbuf_r)
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d <= writeCT$wmAdd_BoollizzieLet21_1_argbuf_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_r = (! writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_d = (writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf :
                                                         writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_r && writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_r) && (! writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_buf <= writeCT$wmAdd_BoollizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) > (sca1_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_r = ((! writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_r)
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet22_1_argbuf,Pointer_CT$wmAdd_Bool) > (writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_r = ((! writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet22_1_argbuf_r)
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d <= writeCT$wmAdd_BoollizzieLet22_1_argbuf_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_r = (! writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_d = (writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf :
                                                         writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_r && writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_r) && (! writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_buf <= writeCT$wmAdd_BoollizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) > (sca0_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_r = ((! writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                               1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_r)
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                   1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_BoollizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf,Pointer_CT$wmAdd_Bool) > (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_r = ((! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_r)
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d <= writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_r = (! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf[0]);
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_d = (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf :
                                                          writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_r && writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_r) && (! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_buf <= writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wmAdd_Bool) : (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb,Pointer_CT$wmAdd_Bool) > (sca3_1_argbuf,Pointer_CT$wmAdd_Bool) */
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d;
  logic writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_r;
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_r = ((! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d[0]) || writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                1'd0};
    else
      if (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_r)
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d <= writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_d;
  Pointer_CT$wmAdd_Bool_t writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_r = (! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf :
                            writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_buf <= writeCT$wmAdd_BoollizzieLet8_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet16_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet16_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet16_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca3_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca3_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet18_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet18_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet18_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (lizzieLet4_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf :
                                    writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet25_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet25_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet25_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca2_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca2_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet26_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet26_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet26_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca1_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca1_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet27_1_argbuf,Pointer_CTmain_mask_Bool) > (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_r = ((! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet27_1_argbuf_r)
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d <= writeCTmain_mask_BoollizzieLet27_1_argbuf_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_r = (! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d = (writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf :
                                                            writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r && writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r) && (! writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_buf <= writeCTmain_mask_BoollizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_mask_Bool) : (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb,Pointer_CTmain_mask_Bool) > (sca0_1_1_argbuf,Pointer_CTmain_mask_Bool) */
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r = ((! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                  1'd0};
    else
      if (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_r)
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_d;
  Pointer_CTmain_mask_Bool_t writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_1_argbuf_d = (writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf :
                              writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                    1'd0};
    else
      if ((sca0_1_1_argbuf_r && writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                      1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCTmain_mask_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet10_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet10_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet10_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet12_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_argbuf_r = ((! writeQTree_BoollizzieLet12_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_argbuf_r)
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet12_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_d = (writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet12_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet12_1_argbuf_rwb_r && writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet12_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet12_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet12_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet12_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet12_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet0_1_1_argbuf_d = (writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet0_1_1_argbuf_r && writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet12_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_r = ((! writeQTree_BoollizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_r)
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_d = (writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet14_1_argbuf_rwb_r && writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet14_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet15_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_argbuf_r = ((! writeQTree_BoollizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_argbuf_r)
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet15_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_d = (writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet15_1_argbuf_rwb_r && writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet15_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet17_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet17_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet17_1_argbuf_r = ((! writeQTree_BoollizzieLet17_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet17_1_argbuf_r)
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet17_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet17_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_d = (writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet17_1_argbuf_rwb_r && writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet17_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet17_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet17_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet17_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet23_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet23_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet23_1_argbuf_r = ((! writeQTree_BoollizzieLet23_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet23_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet23_1_argbuf_r)
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet23_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet23_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_d = (writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet23_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet23_1_argbuf_rwb_r && writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet23_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet23_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet23_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet23_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet23_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet23_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet23_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_r = ((! writeQTree_BoollizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_r)
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_d = (writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet28_1_argbuf_rwb_r && writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet28_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_r = ((! writeQTree_BoollizzieLet3_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_r)
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_d = (writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet3_1_argbuf_rwb_r && writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet3_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet5_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_r = ((! writeQTree_BoollizzieLet4_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_r)
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_d = (writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet4_1_argbuf_rwb_r && writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet4_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet4_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet4_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet4_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_argbuf_d = (writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet6_1_argbuf_r && writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet6_1_argbuf_r) && (! writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet5_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_1_argbuf_r = ((! writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_1_argbuf_r)
        writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet5_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet5_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf :
                                                       writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet5_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet5_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet5_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet7_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet5_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet5_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet7_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_1_argbuf_r = ((! writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_1_argbuf_r)
        writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet7_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet7_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf :
                                                       writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet7_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet7_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet7_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet7_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet7_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_BoollizzieLet7_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet7_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet7_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf :
                                                       writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet9_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet9_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf :
                                  writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet9_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (wsib_2_2,MyDTBool_Bool_Bool) > (wsib_2_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t wsib_2_2_bufchan_d;
  logic wsib_2_2_bufchan_r;
  assign wsib_2_2_r = ((! wsib_2_2_bufchan_d[0]) || wsib_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_2_2_bufchan_d <= 1'd0;
    else if (wsib_2_2_r) wsib_2_2_bufchan_d <= wsib_2_2_d;
  MyDTBool_Bool_Bool_t wsib_2_2_bufchan_buf;
  assign wsib_2_2_bufchan_r = (! wsib_2_2_bufchan_buf[0]);
  assign wsib_2_2_argbuf_d = (wsib_2_2_bufchan_buf[0] ? wsib_2_2_bufchan_buf :
                              wsib_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_2_2_bufchan_buf <= 1'd0;
    else
      if ((wsib_2_2_argbuf_r && wsib_2_2_bufchan_buf[0]))
        wsib_2_2_bufchan_buf <= 1'd0;
      else if (((! wsib_2_2_argbuf_r) && (! wsib_2_2_bufchan_buf[0])))
        wsib_2_2_bufchan_buf <= wsib_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (wsib_2_destruct,MyDTBool_Bool_Bool) > [(wsib_2_1,MyDTBool_Bool_Bool),
                                                                       (wsib_2_2,MyDTBool_Bool_Bool)] */
  logic [1:0] wsib_2_destruct_emitted;
  logic [1:0] wsib_2_destruct_done;
  assign wsib_2_1_d = (wsib_2_destruct_d[0] && (! wsib_2_destruct_emitted[0]));
  assign wsib_2_2_d = (wsib_2_destruct_d[0] && (! wsib_2_destruct_emitted[1]));
  assign wsib_2_destruct_done = (wsib_2_destruct_emitted | ({wsib_2_2_d[0],
                                                             wsib_2_1_d[0]} & {wsib_2_2_r,
                                                                               wsib_2_1_r}));
  assign wsib_2_destruct_r = (& wsib_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_2_destruct_emitted <= 2'd0;
    else
      wsib_2_destruct_emitted <= (wsib_2_destruct_r ? 2'd0 :
                                  wsib_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (wsib_3_2,MyDTBool_Bool_Bool) > (wsib_3_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t wsib_3_2_bufchan_d;
  logic wsib_3_2_bufchan_r;
  assign wsib_3_2_r = ((! wsib_3_2_bufchan_d[0]) || wsib_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_3_2_bufchan_d <= 1'd0;
    else if (wsib_3_2_r) wsib_3_2_bufchan_d <= wsib_3_2_d;
  MyDTBool_Bool_Bool_t wsib_3_2_bufchan_buf;
  assign wsib_3_2_bufchan_r = (! wsib_3_2_bufchan_buf[0]);
  assign wsib_3_2_argbuf_d = (wsib_3_2_bufchan_buf[0] ? wsib_3_2_bufchan_buf :
                              wsib_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_3_2_bufchan_buf <= 1'd0;
    else
      if ((wsib_3_2_argbuf_r && wsib_3_2_bufchan_buf[0]))
        wsib_3_2_bufchan_buf <= 1'd0;
      else if (((! wsib_3_2_argbuf_r) && (! wsib_3_2_bufchan_buf[0])))
        wsib_3_2_bufchan_buf <= wsib_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (wsib_3_destruct,MyDTBool_Bool_Bool) > [(wsib_3_1,MyDTBool_Bool_Bool),
                                                                       (wsib_3_2,MyDTBool_Bool_Bool)] */
  logic [1:0] wsib_3_destruct_emitted;
  logic [1:0] wsib_3_destruct_done;
  assign wsib_3_1_d = (wsib_3_destruct_d[0] && (! wsib_3_destruct_emitted[0]));
  assign wsib_3_2_d = (wsib_3_destruct_d[0] && (! wsib_3_destruct_emitted[1]));
  assign wsib_3_destruct_done = (wsib_3_destruct_emitted | ({wsib_3_2_d[0],
                                                             wsib_3_1_d[0]} & {wsib_3_2_r,
                                                                               wsib_3_1_r}));
  assign wsib_3_destruct_r = (& wsib_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_3_destruct_emitted <= 2'd0;
    else
      wsib_3_destruct_emitted <= (wsib_3_destruct_r ? 2'd0 :
                                  wsib_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (wsib_4_destruct,MyDTBool_Bool_Bool) > (wsib_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t wsib_4_destruct_bufchan_d;
  logic wsib_4_destruct_bufchan_r;
  assign wsib_4_destruct_r = ((! wsib_4_destruct_bufchan_d[0]) || wsib_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_4_destruct_bufchan_d <= 1'd0;
    else
      if (wsib_4_destruct_r)
        wsib_4_destruct_bufchan_d <= wsib_4_destruct_d;
  MyDTBool_Bool_Bool_t wsib_4_destruct_bufchan_buf;
  assign wsib_4_destruct_bufchan_r = (! wsib_4_destruct_bufchan_buf[0]);
  assign wsib_4_1_argbuf_d = (wsib_4_destruct_bufchan_buf[0] ? wsib_4_destruct_bufchan_buf :
                              wsib_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wsib_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((wsib_4_1_argbuf_r && wsib_4_destruct_bufchan_buf[0]))
        wsib_4_destruct_bufchan_buf <= 1'd0;
      else if (((! wsib_4_1_argbuf_r) && (! wsib_4_destruct_bufchan_buf[0])))
        wsib_4_destruct_bufchan_buf <= wsib_4_destruct_bufchan_d;
endmodule