`timescale 1ns/1ns
import mMapKron_package::*;

module mMapKron(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Bool_src_d ,
  output logic \\QTree_Bool_src_r ,
  input QTree_Bool_t dummy_write_QTree_Bool_d,
  output logic dummy_write_QTree_Bool_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Bool_t m1adn_0_d,
  output logic m1adn_0_r,
  input Pointer_QTree_Bool_t m2ado_1_d,
  output logic m2ado_1_r,
  output \Word16#_t  forkHP1_QTree_Bool_snk_dout,
  input logic forkHP1_QTree_Bool_snk_rout,
  output Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_dout,
  input logic dummy_write_QTree_Bool_sink_rout,
  output Pointer_QTree_Nat_t \main_map'_Bool_Nat_resbuf_dout ,
  input logic \main_map'_Bool_Nat_resbuf_rout 
  );
  /* --define=INPUTS=((__05CQTree_Bool_src, 0, 1, Go), (dummy_write_QTree_Bool, 66, 73786976294838206464, QTree_Bool), (sourceGo, 0, 1, Go), (m1adn_0, 16, 65536, Pointer_QTree_Bool), (m2ado_1, 16, 65536, Pointer_QTree_Bool)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Bool_snk, 16, 65536, Word16__023), (dummy_write_QTree_Bool_sink, 16, 65536, Pointer_QTree_Bool), (main_map__027_Bool_Nat_resbuf, 16, 65536, Pointer_QTree_Nat)) */
  /* TYPE_START
Nat 16 1 (0,[0]) (1,[16p])
CTmain_map__027_Bool_Nat 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p]) (3,[16p,16p,16p,0,0,16p]) (4,[16p,16p,16p,16p])
QTree_Nat 16 2 (0,[0]) (1,[16p]) (2,[16p,16p,16p,16p]) (3,[0])
QTree_Bool 16 2 (0,[0]) (1,[1]) (2,[16p,16p,16p,16p]) (3,[0])
CTmap__027__027_map__027__027_Bool_Bool_Bool 16 3 (0,[0]) (1,[16p,0,0,1,16p,16p,16p]) (2,[16p,16p,0,0,1,16p,16p]) (3,[16p,16p,16p,0,0,1,16p]) (4,[16p,16p,16p,16p])
CTkron_kron_Bool_Bool_Bool 16 3 (0,[0]) (1,[16p,0,0,16p,16p,16p,16p]) (2,[16p,16p,0,0,16p,16p,16p]) (3,[16p,16p,16p,0,0,16p,16p]) (4,[16p,16p,16p,16p])
TupGo___MyDTNat_Bool___Pointer_Nat 16 0 (0,[0,0,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool 16 0 (0,[0,0,0,16p,16p,16p])
TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map__027_Bool_Nat 16 0 (0,[0,0,0,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap__027__027_map__027__027_Bool_Bool_Bool 16 0 (0,[0,0,0,1,16p,16p])
TupGo___Pointer_Nat___Pointer_Nat 16 0 (0,[0,16p,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool 16 0 (0,[0,0,0,16p,16p])
TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool 16 0 (0,[0,0,0,16p])
TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool 16 0 (0,[0,0,0,1,16p])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go_5_d;
  logic go_5_r;
  Go_t go_6_d;
  logic go_6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  Go_t go__11_d;
  logic go__11_r;
  Go_t go__12_d;
  logic go__12_r;
  Go_t go__13_d;
  logic go__13_r;
  Go_t go__14_d;
  logic go__14_r;
  Go_t go__15_d;
  logic go__15_r;
  Go_t go__16_d;
  logic go__16_r;
  \Word16#_t  initHP_Nat_d;
  logic initHP_Nat_r;
  \Word16#_t  incrHP_Nat_d;
  logic incrHP_Nat_r;
  Go_t incrHP_mergeNat_d;
  logic incrHP_mergeNat_r;
  Go_t incrHP_Nat1_d;
  logic incrHP_Nat1_r;
  Go_t incrHP_Nat2_d;
  logic incrHP_Nat2_r;
  \Word16#_t  addHP_Nat_d;
  logic addHP_Nat_r;
  \Word16#_t  mergeHP_Nat_d;
  logic mergeHP_Nat_r;
  Go_t incrHP_mergeNat_buf_d;
  logic incrHP_mergeNat_buf_r;
  \Word16#_t  mergeHP_Nat_buf_d;
  logic mergeHP_Nat_buf_r;
  \Word16#_t  forkHP1_Nat_d;
  logic forkHP1_Nat_r;
  \Word16#_t  forkHP1_Na2_d;
  logic forkHP1_Na2_r;
  \Word16#_t  forkHP1_Na3_d;
  logic forkHP1_Na3_r;
  C2_t memMergeChoice_Nat_d;
  logic memMergeChoice_Nat_r;
  MemIn_Nat_t memMergeIn_Nat_d;
  logic memMergeIn_Nat_r;
  MemOut_Nat_t memOut_Nat_d;
  logic memOut_Nat_r;
  MemOut_Nat_t memReadOut_Nat_d;
  logic memReadOut_Nat_r;
  MemOut_Nat_t memWriteOut_Nat_d;
  logic memWriteOut_Nat_r;
  MemIn_Nat_t memMergeIn_Nat_dbuf_d;
  logic memMergeIn_Nat_dbuf_r;
  MemIn_Nat_t memMergeIn_Nat_rbuf_d;
  logic memMergeIn_Nat_rbuf_r;
  MemOut_Nat_t memOut_Nat_dbuf_d;
  logic memOut_Nat_dbuf_r;
  MemOut_Nat_t memOut_Nat_rbuf_d;
  logic memOut_Nat_rbuf_r;
  C2_t readMerge_choice_Nat_d;
  logic readMerge_choice_Nat_r;
  Pointer_Nat_t readMerge_data_Nat_d;
  logic readMerge_data_Nat_r;
  Nat_t readPointer_Natxadg_1_argbuf_d;
  logic readPointer_Natxadg_1_argbuf_r;
  Nat_t readPointer_Natyadh_1_argbuf_d;
  logic readPointer_Natyadh_1_argbuf_r;
  \Word16#_t  destructReadIn_Nat_d;
  logic destructReadIn_Nat_r;
  MemIn_Nat_t dconReadIn_Nat_d;
  logic dconReadIn_Nat_r;
  Nat_t destructReadOut_Nat_d;
  logic destructReadOut_Nat_r;
  C4_t writeMerge_choice_Nat_d;
  logic writeMerge_choice_Nat_r;
  Nat_t writeMerge_data_Nat_d;
  logic writeMerge_data_Nat_r;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_d;
  logic writeNatlizzieLet0_1_argbuf_r;
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_d;
  logic writeNatlizzieLet1_1_argbuf_r;
  Pointer_Nat_t writeNatlizzieLet39_1_argbuf_d;
  logic writeNatlizzieLet39_1_argbuf_r;
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_d;
  logic writeNatlizzieLet40_1_argbuf_r;
  MemIn_Nat_t dconWriteIn_Nat_d;
  logic dconWriteIn_Nat_r;
  Pointer_Nat_t dconPtr_Nat_d;
  logic dconPtr_Nat_r;
  Pointer_Nat_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  Pointer_Nat_t demuxWriteResult_Nat_d;
  logic demuxWriteResult_Nat_r;
  \Word16#_t  \initHP_CTmain_map'_Bool_Nat_d ;
  logic \initHP_CTmain_map'_Bool_Nat_r ;
  \Word16#_t  \incrHP_CTmain_map'_Bool_Nat_d ;
  logic \incrHP_CTmain_map'_Bool_Nat_r ;
  Go_t \incrHP_mergeCTmain_map'_Bool_Nat_d ;
  logic \incrHP_mergeCTmain_map'_Bool_Nat_r ;
  Go_t \incrHP_CTmain_map'_Bool_Nat1_d ;
  logic \incrHP_CTmain_map'_Bool_Nat1_r ;
  Go_t \incrHP_CTmain_map'_Bool_Nat2_d ;
  logic \incrHP_CTmain_map'_Bool_Nat2_r ;
  \Word16#_t  \addHP_CTmain_map'_Bool_Nat_d ;
  logic \addHP_CTmain_map'_Bool_Nat_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Bool_Nat_d ;
  logic \mergeHP_CTmain_map'_Bool_Nat_r ;
  Go_t \incrHP_mergeCTmain_map'_Bool_Nat_buf_d ;
  logic \incrHP_mergeCTmain_map'_Bool_Nat_buf_r ;
  \Word16#_t  \mergeHP_CTmain_map'_Bool_Nat_buf_d ;
  logic \mergeHP_CTmain_map'_Bool_Nat_buf_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Bool_Nat_d ;
  logic \forkHP1_CTmain_map'_Bool_Nat_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Bool_Na2_d ;
  logic \forkHP1_CTmain_map'_Bool_Na2_r ;
  \Word16#_t  \forkHP1_CTmain_map'_Bool_Na3_d ;
  logic \forkHP1_CTmain_map'_Bool_Na3_r ;
  C2_t \memMergeChoice_CTmain_map'_Bool_Nat_d ;
  logic \memMergeChoice_CTmain_map'_Bool_Nat_r ;
  \MemIn_CTmain_map'_Bool_Nat_t  \memMergeIn_CTmain_map'_Bool_Nat_d ;
  logic \memMergeIn_CTmain_map'_Bool_Nat_r ;
  \MemOut_CTmain_map'_Bool_Nat_t  \memOut_CTmain_map'_Bool_Nat_d ;
  logic \memOut_CTmain_map'_Bool_Nat_r ;
  \MemOut_CTmain_map'_Bool_Nat_t  \memReadOut_CTmain_map'_Bool_Nat_d ;
  logic \memReadOut_CTmain_map'_Bool_Nat_r ;
  \MemOut_CTmain_map'_Bool_Nat_t  \memWriteOut_CTmain_map'_Bool_Nat_d ;
  logic \memWriteOut_CTmain_map'_Bool_Nat_r ;
  \MemIn_CTmain_map'_Bool_Nat_t  \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d ;
  logic \memMergeIn_CTmain_map'_Bool_Nat_dbuf_r ;
  \MemIn_CTmain_map'_Bool_Nat_t  \memMergeIn_CTmain_map'_Bool_Nat_rbuf_d ;
  logic \memMergeIn_CTmain_map'_Bool_Nat_rbuf_r ;
  \MemOut_CTmain_map'_Bool_Nat_t  \memOut_CTmain_map'_Bool_Nat_dbuf_d ;
  logic \memOut_CTmain_map'_Bool_Nat_dbuf_r ;
  \MemOut_CTmain_map'_Bool_Nat_t  \memOut_CTmain_map'_Bool_Nat_rbuf_d ;
  logic \memOut_CTmain_map'_Bool_Nat_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmain_map'_Bool_Nat_d ;
  logic \destructReadIn_CTmain_map'_Bool_Nat_r ;
  \MemIn_CTmain_map'_Bool_Nat_t  \dconReadIn_CTmain_map'_Bool_Nat_d ;
  logic \dconReadIn_CTmain_map'_Bool_Nat_r ;
  \CTmain_map'_Bool_Nat_t  \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmain_map'_Bool_Nat_d ;
  logic \writeMerge_choice_CTmain_map'_Bool_Nat_r ;
  \CTmain_map'_Bool_Nat_t  \writeMerge_data_CTmain_map'_Bool_Nat_d ;
  logic \writeMerge_data_CTmain_map'_Bool_Nat_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_r ;
  \MemIn_CTmain_map'_Bool_Nat_t  \dconWriteIn_CTmain_map'_Bool_Nat_d ;
  logic \dconWriteIn_CTmain_map'_Bool_Nat_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \dconPtr_CTmain_map'_Bool_Nat_d ;
  logic \dconPtr_CTmain_map'_Bool_Nat_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  \Pointer_CTmain_map'_Bool_Nat_t  \demuxWriteResult_CTmain_map'_Bool_Nat_d ;
  logic \demuxWriteResult_CTmain_map'_Bool_Nat_r ;
  \Word16#_t  initHP_QTree_Nat_d;
  logic initHP_QTree_Nat_r;
  \Word16#_t  incrHP_QTree_Nat_d;
  logic incrHP_QTree_Nat_r;
  Go_t incrHP_mergeQTree_Nat_d;
  logic incrHP_mergeQTree_Nat_r;
  Go_t incrHP_QTree_Nat1_d;
  logic incrHP_QTree_Nat1_r;
  Go_t incrHP_QTree_Nat2_d;
  logic incrHP_QTree_Nat2_r;
  \Word16#_t  addHP_QTree_Nat_d;
  logic addHP_QTree_Nat_r;
  \Word16#_t  mergeHP_QTree_Nat_d;
  logic mergeHP_QTree_Nat_r;
  Go_t incrHP_mergeQTree_Nat_buf_d;
  logic incrHP_mergeQTree_Nat_buf_r;
  \Word16#_t  mergeHP_QTree_Nat_buf_d;
  logic mergeHP_QTree_Nat_buf_r;
  \Word16#_t  forkHP1_QTree_Nat_d;
  logic forkHP1_QTree_Nat_r;
  \Word16#_t  forkHP1_QTree_Na2_d;
  logic forkHP1_QTree_Na2_r;
  \Word16#_t  forkHP1_QTree_Na3_d;
  logic forkHP1_QTree_Na3_r;
  MemOut_QTree_Nat_t memWriteOut_QTree_Nat_d;
  logic memWriteOut_QTree_Nat_r;
  C5_t writeMerge_choice_QTree_Nat_d;
  logic writeMerge_choice_QTree_Nat_r;
  QTree_Nat_t writeMerge_data_QTree_Nat_d;
  logic writeMerge_data_QTree_Nat_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_d;
  logic writeQTree_NatlizzieLet11_1_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_d;
  logic writeQTree_NatlizzieLet33_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_d;
  logic writeQTree_NatlizzieLet7_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_d;
  logic writeQTree_NatlizzieLet8_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_d;
  logic writeQTree_NatlizzieLet9_1_argbuf_r;
  MemIn_QTree_Nat_t dconWriteIn_QTree_Nat_d;
  logic dconWriteIn_QTree_Nat_r;
  Pointer_QTree_Nat_t dconPtr_QTree_Nat_d;
  logic dconPtr_QTree_Nat_r;
  Pointer_QTree_Nat_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Pointer_QTree_Nat_t demuxWriteResult_QTree_Nat_d;
  logic demuxWriteResult_QTree_Nat_r;
  \Word16#_t  initHP_QTree_Bool_d;
  logic initHP_QTree_Bool_r;
  \Word16#_t  incrHP_QTree_Bool_d;
  logic incrHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_d;
  logic incrHP_mergeQTree_Bool_r;
  Go_t incrHP_QTree_Bool1_d;
  logic incrHP_QTree_Bool1_r;
  Go_t incrHP_QTree_Bool2_d;
  logic incrHP_QTree_Bool2_r;
  \Word16#_t  addHP_QTree_Bool_d;
  logic addHP_QTree_Bool_r;
  \Word16#_t  mergeHP_QTree_Bool_d;
  logic mergeHP_QTree_Bool_r;
  Go_t incrHP_mergeQTree_Bool_buf_d;
  logic incrHP_mergeQTree_Bool_buf_r;
  \Word16#_t  mergeHP_QTree_Bool_buf_d;
  logic mergeHP_QTree_Bool_buf_r;
  Go_t go_1_dummy_write_QTree_Bool_d;
  logic go_1_dummy_write_QTree_Bool_r;
  Go_t go_2_dummy_write_QTree_Bool_d;
  logic go_2_dummy_write_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_d;
  logic forkHP1_QTree_Bool_r;
  \Word16#_t  forkHP1_QTree_Bool_snk_d;
  logic forkHP1_QTree_Bool_snk_r;
  \Word16#_t  forkHP1_QTree_Boo3_d;
  logic forkHP1_QTree_Boo3_r;
  \Word16#_t  forkHP1_QTree_Boo4_d;
  logic forkHP1_QTree_Boo4_r;
  C2_t memMergeChoice_QTree_Bool_d;
  logic memMergeChoice_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_d;
  logic memMergeIn_QTree_Bool_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_d;
  logic memOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memReadOut_QTree_Bool_d;
  logic memReadOut_QTree_Bool_r;
  MemOut_QTree_Bool_t memWriteOut_QTree_Bool_d;
  logic memWriteOut_QTree_Bool_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_dbuf_d;
  logic memMergeIn_QTree_Bool_dbuf_r;
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_rbuf_d;
  logic memMergeIn_QTree_Bool_rbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_dbuf_d;
  logic memOut_QTree_Bool_dbuf_r;
  MemOut_QTree_Bool_t memOut_QTree_Bool_rbuf_d;
  logic memOut_QTree_Bool_rbuf_r;
  C3_t readMerge_choice_QTree_Bool_d;
  logic readMerge_choice_QTree_Bool_r;
  Pointer_QTree_Bool_t readMerge_data_QTree_Bool_d;
  logic readMerge_data_QTree_Bool_r;
  QTree_Bool_t readPointer_QTree_Boolm1ad9_1_argbuf_d;
  logic readPointer_QTree_Boolm1ad9_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_BoolmacS_1_argbuf_d;
  logic readPointer_QTree_BoolmacS_1_argbuf_r;
  QTree_Bool_t readPointer_QTree_Boolmad1_1_argbuf_d;
  logic readPointer_QTree_Boolmad1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Bool_d;
  logic destructReadIn_QTree_Bool_r;
  MemIn_QTree_Bool_t dconReadIn_QTree_Bool_d;
  logic dconReadIn_QTree_Bool_r;
  QTree_Bool_t destructReadOut_QTree_Bool_d;
  logic destructReadOut_QTree_Bool_r;
  C9_t writeMerge_choice_QTree_Bool_d;
  logic writeMerge_choice_QTree_Bool_r;
  QTree_Bool_t writeMerge_data_QTree_Bool_d;
  logic writeMerge_data_QTree_Bool_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_r;
  Pointer_QTree_Bool_t dummy_write_QTree_Bool_sink_d;
  logic dummy_write_QTree_Bool_sink_r;
  MemIn_QTree_Bool_t dconWriteIn_QTree_Bool_d;
  logic dconWriteIn_QTree_Bool_r;
  Pointer_QTree_Bool_t dconPtr_QTree_Bool_d;
  logic dconPtr_QTree_Bool_r;
  Pointer_QTree_Bool_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Pointer_QTree_Bool_t demuxWriteResult_QTree_Bool_d;
  logic demuxWriteResult_QTree_Bool_r;
  \Word16#_t  \initHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \initHP_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \incrHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_CTmap''_map''_Bool_Bool_Bool1_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool1_r ;
  Go_t \incrHP_CTmap''_map''_Bool_Bool_Bool2_d ;
  logic \incrHP_CTmap''_map''_Bool_Bool_Bool2_r ;
  \Word16#_t  \addHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \addHP_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_r ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ;
  \Word16#_t  \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d ;
  logic \forkHP1_CTmap''_map''_Bool_Bool_Boo3_r ;
  C2_t \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memReadOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memReadOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memWriteOut_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \memWriteOut_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r ;
  \Word16#_t  \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \destructReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r ;
  C5_t \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_r ;
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \dconPtr_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \dconPtr_CTmap''_map''_Bool_Bool_Bool_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d ;
  logic \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ;
  \Word16#_t  initHP_CTkron_kron_Bool_Bool_Bool_d;
  logic initHP_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  incrHP_CTkron_kron_Bool_Bool_Bool_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_CTkron_kron_Bool_Bool_Bool1_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool1_r;
  Go_t incrHP_CTkron_kron_Bool_Bool_Bool2_d;
  logic incrHP_CTkron_kron_Bool_Bool_Bool2_r;
  \Word16#_t  addHP_CTkron_kron_Bool_Bool_Bool_d;
  logic addHP_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_r;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Bool_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Bool_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Boo2_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Boo2_r;
  \Word16#_t  forkHP1_CTkron_kron_Bool_Bool_Boo3_d;
  logic forkHP1_CTkron_kron_Bool_Bool_Boo3_r;
  C2_t memMergeChoice_CTkron_kron_Bool_Bool_Bool_d;
  logic memMergeChoice_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memReadOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memReadOut_CTkron_kron_Bool_Bool_Bool_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memWriteOut_CTkron_kron_Bool_Bool_Bool_d;
  logic memWriteOut_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  logic memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r;
  \Word16#_t  destructReadIn_CTkron_kron_Bool_Bool_Bool_d;
  logic destructReadIn_CTkron_kron_Bool_Bool_Bool_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t dconReadIn_CTkron_kron_Bool_Bool_Bool_d;
  logic dconReadIn_CTkron_kron_Bool_Bool_Bool_r;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d;
  logic writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r;
  CTkron_kron_Bool_Bool_Bool_t writeMerge_data_CTkron_kron_Bool_Bool_Bool_d;
  logic writeMerge_data_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_r;
  MemIn_CTkron_kron_Bool_Bool_Bool_t dconWriteIn_CTkron_kron_Bool_Bool_Bool_d;
  logic dconWriteIn_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t dconPtr_CTkron_kron_Bool_Bool_Bool_d;
  logic dconPtr_CTkron_kron_Bool_Bool_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  Pointer_CTkron_kron_Bool_Bool_Bool_t demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d;
  logic demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r;
  Go_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r;
  MyDTBool_Bool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r;
  MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r;
  MyDTBool_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTBool_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTBool_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t es_0_2_1_d;
  logic es_0_2_1_r;
  MyBool_t es_0_2_2_d;
  logic es_0_2_2_r;
  MyBool_t es_0_2_3_d;
  logic es_0_2_3_r;
  Go_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r;
  MyDTBool_Bool_Bool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r;
  MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_r;
  MyDTBool_Bool_Bool_t arg0_4_1_d;
  logic arg0_4_1_r;
  MyDTBool_Bool_Bool_t arg0_4_2_d;
  logic arg0_4_2_r;
  MyDTBool_Bool_Bool_t arg0_4_3_d;
  logic arg0_4_3_r;
  MyDTBool_Bool_Bool_t arg0_4_4_d;
  logic arg0_4_4_r;
  MyBool_t xacw_1_1_d;
  logic xacw_1_1_r;
  MyBool_t xacw_1_2_d;
  logic xacw_1_2_r;
  Go_t applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d;
  logic applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_r;
  MyDTBool_Nat_t applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d;
  logic applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_r;
  MyBool_t applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d;
  logic applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_r;
  MyDTBool_Nat_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTBool_Nat_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTBool_Nat_t arg0_2_3_d;
  logic arg0_2_3_r;
  Pointer_Nat_t xacw_1_d;
  logic xacw_1_r;
  Pointer_Nat_t xacw_2_d;
  logic xacw_2_r;
  Go_t applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d;
  logic applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_r;
  MyDTNat_Bool_t applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d;
  logic applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_r;
  Pointer_Nat_t applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d;
  logic applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_r;
  MyDTNat_Bool_t arg0_6_1_d;
  logic arg0_6_1_r;
  MyDTNat_Bool_t arg0_6_2_d;
  logic arg0_6_2_r;
  MyDTNat_Bool_t arg0_6_3_d;
  logic arg0_6_3_r;
  MyBool_t es_0_1_1_d;
  logic es_0_1_1_r;
  MyBool_t es_0_1_2_d;
  logic es_0_1_2_r;
  MyBool_t es_0_1_3_d;
  logic es_0_1_3_r;
  MyBool_t arg0_1Dcon_main1_d;
  logic arg0_1Dcon_main1_r;
  MyBool_t arg0_1Dcon_main1_1_d;
  logic arg0_1Dcon_main1_1_r;
  MyBool_t arg0_1Dcon_main1_2_d;
  logic arg0_1Dcon_main1_2_r;
  Go_t arg0_1Dcon_main1_1MyFalse_d;
  logic arg0_1Dcon_main1_1MyFalse_r;
  Go_t arg0_1Dcon_main1_1MyTrue_d;
  logic arg0_1Dcon_main1_1MyTrue_r;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTrue_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTrue_r;
  MyBool_t applyfnBool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_5_resbuf_r;
  MyBool_t arg0_1Dcon_main1_1MyTrue_1MyFalse_d;
  logic arg0_1Dcon_main1_1MyTrue_1MyFalse_r;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r;
  Go_t arg0_2Dcon_main1_d;
  logic arg0_2Dcon_main1_r;
  MyBool_t arg0_2_1Dcon_to_nat_d;
  logic arg0_2_1Dcon_to_nat_r;
  MyBool_t arg0_2_1Dcon_to_nat_1_d;
  logic arg0_2_1Dcon_to_nat_1_r;
  MyBool_t arg0_2_1Dcon_to_nat_2_d;
  logic arg0_2_1Dcon_to_nat_2_r;
  Go_t arg0_2_1Dcon_to_nat_1MyFalse_d;
  logic arg0_2_1Dcon_to_nat_1MyFalse_r;
  Go_t arg0_2_1Dcon_to_nat_1MyTrue_d;
  logic arg0_2_1Dcon_to_nat_1MyTrue_r;
  Nat_t arg0_2_1Dcon_to_nat_1MyFalse_1Zero_d;
  logic arg0_2_1Dcon_to_nat_1MyFalse_1Zero_r;
  Nat_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_d;
  logic arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_r;
  TupGo_t to_nat1TupGo_1_d;
  logic to_nat1TupGo_1_r;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d;
  logic writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_r;
  Go_t arg0_2_2Dcon_to_nat_d;
  logic arg0_2_2Dcon_to_nat_r;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_d;
  logic writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_r;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r;
  MyBool_t \arg0_4_1Dcon_&&_d ;
  logic \arg0_4_1Dcon_&&_r ;
  MyBool_t \arg0_4_2Dcon_&&_d ;
  logic \arg0_4_2Dcon_&&_r ;
  MyBool_t \arg0_4_2Dcon_&&_1_d ;
  logic \arg0_4_2Dcon_&&_1_r ;
  MyBool_t \arg0_4_2Dcon_&&_2_d ;
  logic \arg0_4_2Dcon_&&_2_r ;
  MyBool_t \arg0_4_2Dcon_&&_3_d ;
  logic \arg0_4_2Dcon_&&_3_r ;
  MyBool_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  MyBool_t \arg0_4_2Dcon_&&_1MyTrue_d ;
  logic \arg0_4_2Dcon_&&_1MyTrue_r ;
  Go_t \arg0_4_2Dcon_&&_2MyFalse_d ;
  logic \arg0_4_2Dcon_&&_2MyFalse_r ;
  Go_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  MyBool_t \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_d ;
  logic \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_r ;
  MyBool_t applyfnBool_Bool_Bool_5_resbuf_d;
  logic applyfnBool_Bool_Bool_5_resbuf_r;
  MyBool_t \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d ;
  logic \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_r ;
  Go_t \arg0_4_3Dcon_&&_d ;
  logic \arg0_4_3Dcon_&&_r ;
  MyBool_t \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_d ;
  logic \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_r ;
  Pointer_Nat_t arg0_6_1Dcon_is_z_nut_d;
  logic arg0_6_1Dcon_is_z_nut_r;
  Pointer_Nat_t arg0_6_1Dcon_is_z_nut_1_argbuf_d;
  logic arg0_6_1Dcon_is_z_nut_1_argbuf_r;
  Go_t arg0_6_2Dcon_is_z_nut_d;
  logic arg0_6_2Dcon_is_z_nut_r;
  Go_t arg0_6_2Dcon_is_z_nut_1_d;
  logic arg0_6_2Dcon_is_z_nut_1_r;
  Go_t arg0_6_2Dcon_is_z_nut_2_d;
  logic arg0_6_2Dcon_is_z_nut_2_r;
  Nat_t arg0_6_2Dcon_is_z_nut_1Zero_d;
  logic arg0_6_2Dcon_is_z_nut_1Zero_r;
  Nat_t lizzieLet1_1_argbuf_d;
  logic lizzieLet1_1_argbuf_r;
  Go_t arg0_6_2Dcon_is_z_nut_2_argbuf_d;
  logic arg0_6_2Dcon_is_z_nut_2_argbuf_r;
  TupGo___Pointer_Nat___Pointer_Nat_t eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d;
  logic eqNatTupGo___Pointer_Nat___Pointer_Nat_1_r;
  MyBool_t eqNat_1_mux_d;
  logic eqNat_1_mux_r;
  Go_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_r;
  MyDTBool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_r;
  MyDTBool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r;
  Go_t call_kron_kron_Bool_Bool_Bool_initBufi_d;
  logic call_kron_kron_Bool_Bool_Bool_initBufi_r;
  C5_t go_6_goMux_choice_d;
  logic go_6_goMux_choice_r;
  Go_t go_6_goMux_data_d;
  logic go_6_goMux_data_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork1_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork1_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork2_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork2_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork3_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork3_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork4_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork4_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork5_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork5_r;
  Go_t call_kron_kron_Bool_Bool_Bool_unlockFork6_d;
  logic call_kron_kron_Bool_Bool_Bool_unlockFork6_r;
  Go_t call_kron_kron_Bool_Bool_Bool_initBuf_d;
  logic call_kron_kron_Bool_Bool_Bool_initBuf_r;
  Go_t call_kron_kron_Bool_Bool_Bool_goMux1_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux1_r;
  MyDTBool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux2_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux2_r;
  MyDTBool_Bool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux3_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux3_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_Bool_goMux4_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux4_r;
  Pointer_QTree_Bool_t call_kron_kron_Bool_Bool_Bool_goMux5_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux5_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_Bool_goMux6_d;
  logic call_kron_kron_Bool_Bool_Bool_goMux6_r;
  Go_t \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_r ;
  MyDTNat_Bool_t \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_r ;
  MyDTBool_Nat_t \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_r ;
  Pointer_QTree_Bool_t \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_r ;
  Go_t \call_main_map'_Bool_Nat_initBufi_d ;
  logic \call_main_map'_Bool_Nat_initBufi_r ;
  C5_t go_7_goMux_choice_d;
  logic go_7_goMux_choice_r;
  Go_t go_7_goMux_data_d;
  logic go_7_goMux_data_r;
  Go_t \call_main_map'_Bool_Nat_unlockFork1_d ;
  logic \call_main_map'_Bool_Nat_unlockFork1_r ;
  Go_t \call_main_map'_Bool_Nat_unlockFork2_d ;
  logic \call_main_map'_Bool_Nat_unlockFork2_r ;
  Go_t \call_main_map'_Bool_Nat_unlockFork3_d ;
  logic \call_main_map'_Bool_Nat_unlockFork3_r ;
  Go_t \call_main_map'_Bool_Nat_unlockFork4_d ;
  logic \call_main_map'_Bool_Nat_unlockFork4_r ;
  Go_t \call_main_map'_Bool_Nat_unlockFork5_d ;
  logic \call_main_map'_Bool_Nat_unlockFork5_r ;
  Go_t \call_main_map'_Bool_Nat_initBuf_d ;
  logic \call_main_map'_Bool_Nat_initBuf_r ;
  Go_t \call_main_map'_Bool_Nat_goMux1_d ;
  logic \call_main_map'_Bool_Nat_goMux1_r ;
  MyDTNat_Bool_t \call_main_map'_Bool_Nat_goMux2_d ;
  logic \call_main_map'_Bool_Nat_goMux2_r ;
  MyDTBool_Nat_t \call_main_map'_Bool_Nat_goMux3_d ;
  logic \call_main_map'_Bool_Nat_goMux3_r ;
  Pointer_QTree_Bool_t \call_main_map'_Bool_Nat_goMux4_d ;
  logic \call_main_map'_Bool_Nat_goMux4_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  \call_main_map'_Bool_Nat_goMux5_d ;
  logic \call_main_map'_Bool_Nat_goMux5_r ;
  Go_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_r ;
  MyDTBool_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_r ;
  MyDTBool_Bool_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_r ;
  MyBool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_r ;
  Pointer_QTree_Bool_t \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_initBufi_d ;
  logic \call_map''_map''_Bool_Bool_Bool_initBufi_r ;
  C5_t go_8_goMux_choice_d;
  logic go_8_goMux_choice_r;
  Go_t go_8_goMux_data_d;
  logic go_8_goMux_data_r;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork1_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork1_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork2_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork3_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork3_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork4_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork4_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork5_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork5_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_unlockFork6_d ;
  logic \call_map''_map''_Bool_Bool_Bool_unlockFork6_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_initBuf_d ;
  logic \call_map''_map''_Bool_Bool_Bool_initBuf_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_goMux1_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux1_r ;
  MyDTBool_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux2_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux2_r ;
  MyDTBool_Bool_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux3_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux3_r ;
  MyBool_t \call_map''_map''_Bool_Bool_Bool_goMux4_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux4_r ;
  Pointer_QTree_Bool_t \call_map''_map''_Bool_Bool_Bool_goMux5_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux5_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_Bool_goMux6_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goMux6_r ;
  Go_t eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d;
  logic eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_r;
  Pointer_Nat_t eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d;
  logic eqNatTupGo___Pointer_Nat___Pointer_Natxadg_r;
  Pointer_Nat_t eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d;
  logic eqNatTupGo___Pointer_Nat___Pointer_Natyadh_r;
  MyBool_t applyfnNat_Bool_5_resbuf_d;
  logic applyfnNat_Bool_5_resbuf_r;
  Go_t eqNat_initBufi_d;
  logic eqNat_initBufi_r;
  C2_t go_9_goMux_choice_d;
  logic go_9_goMux_choice_r;
  Go_t go_9_goMux_data_d;
  logic go_9_goMux_data_r;
  Go_t eqNat_unlockFork1_d;
  logic eqNat_unlockFork1_r;
  Go_t eqNat_unlockFork2_d;
  logic eqNat_unlockFork2_r;
  Go_t eqNat_unlockFork3_d;
  logic eqNat_unlockFork3_r;
  Go_t eqNat_initBuf_d;
  logic eqNat_initBuf_r;
  Go_t eqNat_goMux1_d;
  logic eqNat_goMux1_r;
  Pointer_Nat_t eqNat_goMux2_d;
  logic eqNat_goMux2_r;
  Pointer_Nat_t eqNat_goMux3_d;
  logic eqNat_goMux3_r;
  Go_t es_0_1_1MyFalse_d;
  logic es_0_1_1MyFalse_r;
  Go_t es_0_1_1MyTrue_d;
  logic es_0_1_1MyTrue_r;
  Go_t es_0_1_1MyFalse_1_argbuf_d;
  logic es_0_1_1MyFalse_1_argbuf_r;
  Go_t es_0_1_1MyTrue_1_d;
  logic es_0_1_1MyTrue_1_r;
  Go_t es_0_1_1MyTrue_2_d;
  logic es_0_1_1MyTrue_2_r;
  QTree_Nat_t es_0_1_1MyTrue_1QNone_Nat_d;
  logic es_0_1_1MyTrue_1QNone_Nat_r;
  QTree_Nat_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t es_0_1_1MyTrue_2_argbuf_d;
  logic es_0_1_1MyTrue_2_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyFalse_d;
  logic es_0_1_2MyFalse_r;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyTrue_d;
  logic es_0_1_2MyTrue_r;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyFalse_1_argbuf_d;
  logic es_0_1_2MyFalse_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyTrue_1_argbuf_d;
  logic es_0_1_2MyTrue_1_argbuf_r;
  Pointer_Nat_t es_0_1_3MyFalse_d;
  logic es_0_1_3MyFalse_r;
  Pointer_Nat_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  QTree_Nat_t es_0_1_3MyFalse_1QVal_Nat_d;
  logic es_0_1_3MyFalse_1QVal_Nat_r;
  QTree_Nat_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Go_t es_0_2_1MyFalse_d;
  logic es_0_2_1MyFalse_r;
  Go_t es_0_2_1MyTrue_d;
  logic es_0_2_1MyTrue_r;
  Go_t es_0_2_1MyFalse_1_argbuf_d;
  logic es_0_2_1MyFalse_1_argbuf_r;
  Go_t es_0_2_1MyTrue_1_d;
  logic es_0_2_1MyTrue_1_r;
  Go_t es_0_2_1MyTrue_2_d;
  logic es_0_2_1MyTrue_2_r;
  QTree_Bool_t es_0_2_1MyTrue_1QNone_Bool_d;
  logic es_0_2_1MyTrue_1QNone_Bool_r;
  QTree_Bool_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Go_t es_0_2_1MyTrue_2_argbuf_d;
  logic es_0_2_1MyTrue_2_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyFalse_d;
  logic es_0_2_2MyFalse_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyTrue_d;
  logic es_0_2_2MyTrue_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyFalse_1_argbuf_d;
  logic es_0_2_2MyFalse_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyTrue_1_argbuf_d;
  logic es_0_2_2MyTrue_1_argbuf_r;
  MyBool_t es_0_2_3MyFalse_d;
  logic es_0_2_3MyFalse_r;
  MyBool_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  QTree_Bool_t es_0_2_3MyFalse_1QVal_Bool_d;
  logic es_0_2_3MyFalse_1QVal_Bool_r;
  QTree_Bool_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  MyDTBool_Nat_t gacR_2_2_argbuf_d;
  logic gacR_2_2_argbuf_r;
  MyDTBool_Nat_t gacR_2_1_d;
  logic gacR_2_1_r;
  MyDTBool_Nat_t gacR_2_2_d;
  logic gacR_2_2_r;
  MyDTBool_Nat_t gacR_3_2_argbuf_d;
  logic gacR_3_2_argbuf_r;
  MyDTBool_Nat_t gacR_3_1_d;
  logic gacR_3_1_r;
  MyDTBool_Nat_t gacR_3_2_d;
  logic gacR_3_2_r;
  MyDTBool_Nat_t gacR_4_1_argbuf_d;
  logic gacR_4_1_argbuf_r;
  MyDTBool_Bool_Bool_t gacZ_2_2_argbuf_d;
  logic gacZ_2_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacZ_2_1_d;
  logic gacZ_2_1_r;
  MyDTBool_Bool_Bool_t gacZ_2_2_d;
  logic gacZ_2_2_r;
  MyDTBool_Bool_Bool_t gacZ_3_2_argbuf_d;
  logic gacZ_3_2_argbuf_r;
  MyDTBool_Bool_Bool_t gacZ_3_1_d;
  logic gacZ_3_1_r;
  MyDTBool_Bool_Bool_t gacZ_3_2_d;
  logic gacZ_3_2_r;
  MyDTBool_Bool_Bool_t gacZ_4_1_argbuf_d;
  logic gacZ_4_1_argbuf_r;
  MyDTBool_Bool_Bool_t gad8_2_2_argbuf_d;
  logic gad8_2_2_argbuf_r;
  MyDTBool_Bool_Bool_t gad8_2_1_d;
  logic gad8_2_1_r;
  MyDTBool_Bool_Bool_t gad8_2_2_d;
  logic gad8_2_2_r;
  MyDTBool_Bool_Bool_t gad8_3_2_argbuf_d;
  logic gad8_3_2_argbuf_r;
  MyDTBool_Bool_Bool_t gad8_3_1_d;
  logic gad8_3_1_r;
  MyDTBool_Bool_Bool_t gad8_3_2_d;
  logic gad8_3_2_r;
  MyDTBool_Bool_Bool_t gad8_4_1_argbuf_d;
  logic gad8_4_1_argbuf_r;
  MyDTBool_Nat_t go_1Dcon_to_nat_d;
  logic go_1Dcon_to_nat_r;
  CTkron_kron_Bool_Bool_Bool_t go_10_1Lkron_kron_Bool_Bool_Boolsbos_d;
  logic go_10_1Lkron_kron_Bool_Bool_Boolsbos_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  Go_t go_10_2_argbuf_d;
  logic go_10_2_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_t call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d;
  logic call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r;
  \CTmain_map'_Bool_Nat_t  \go_11_1Lmain_map'_Bool_Natsbos_d ;
  logic \go_11_1Lmain_map'_Bool_Natsbos_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  Go_t go_11_2_argbuf_d;
  logic go_11_2_argbuf_r;
  \TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_t  \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d ;
  logic \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_d ;
  logic \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet23_1_argbuf_d;
  logic lizzieLet23_1_argbuf_r;
  Go_t go_12_2_argbuf_d;
  logic go_12_2_argbuf_r;
  \TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_t  \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d ;
  logic \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r ;
  C4_t go_13_goMux_choice_1_d;
  logic go_13_goMux_choice_1_r;
  C4_t go_13_goMux_choice_2_d;
  logic go_13_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C5_t go_14_goMux_choice_1_d;
  logic go_14_goMux_choice_1_r;
  C5_t go_14_goMux_choice_2_d;
  logic go_14_goMux_choice_2_r;
  Pointer_QTree_Nat_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTmain_map'_Bool_Nat_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C5_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C5_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  Pointer_QTree_Bool_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  Nat_t lizzieLet39_1_argbuf_d;
  logic lizzieLet39_1_argbuf_r;
  MyDTBool_Nat_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  MyDTNat_Bool_t go_2Dcon_is_z_nut_d;
  logic go_2Dcon_is_z_nut_r;
  MyDTNat_Bool_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  MyDTBool_Bool_Bool_t \go_3Dcon_&&_d ;
  logic \go_3Dcon_&&_r ;
  MyDTBool_Bool_Bool_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  MyDTBool_Bool_t go_4Dcon_main1_d;
  logic go_4Dcon_main1_r;
  MyDTBool_Bool_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t go_5_argbuf_d;
  logic go_5_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r;
  Go_t go_6_argbuf_d;
  logic go_6_argbuf_r;
  TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_r ;
  C5_t go_6_goMux_choice_1_d;
  logic go_6_goMux_choice_1_r;
  C5_t go_6_goMux_choice_2_d;
  logic go_6_goMux_choice_2_r;
  C5_t go_6_goMux_choice_3_d;
  logic go_6_goMux_choice_3_r;
  C5_t go_6_goMux_choice_4_d;
  logic go_6_goMux_choice_4_r;
  C5_t go_6_goMux_choice_5_d;
  logic go_6_goMux_choice_5_r;
  MyDTBool_Bool_t isZad7_goMux_mux_d;
  logic isZad7_goMux_mux_r;
  MyDTBool_Bool_Bool_t gad8_goMux_mux_d;
  logic gad8_goMux_mux_r;
  Pointer_QTree_Bool_t m1ad9_goMux_mux_d;
  logic m1ad9_goMux_mux_r;
  Pointer_QTree_Bool_t m2ada_goMux_mux_d;
  logic m2ada_goMux_mux_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_7_goMux_choice_1_d;
  logic go_7_goMux_choice_1_r;
  C5_t go_7_goMux_choice_2_d;
  logic go_7_goMux_choice_2_r;
  C5_t go_7_goMux_choice_3_d;
  logic go_7_goMux_choice_3_r;
  C5_t go_7_goMux_choice_4_d;
  logic go_7_goMux_choice_4_r;
  MyDTNat_Bool_t isZacQ_goMux_mux_d;
  logic isZacQ_goMux_mux_r;
  MyDTBool_Nat_t gacR_goMux_mux_d;
  logic gacR_goMux_mux_r;
  Pointer_QTree_Bool_t macS_goMux_mux_d;
  logic macS_goMux_mux_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_8_goMux_choice_1_d;
  logic go_8_goMux_choice_1_r;
  C5_t go_8_goMux_choice_2_d;
  logic go_8_goMux_choice_2_r;
  C5_t go_8_goMux_choice_3_d;
  logic go_8_goMux_choice_3_r;
  C5_t go_8_goMux_choice_4_d;
  logic go_8_goMux_choice_4_r;
  C5_t go_8_goMux_choice_5_d;
  logic go_8_goMux_choice_5_r;
  MyDTBool_Bool_t isZacY_goMux_mux_d;
  logic isZacY_goMux_mux_r;
  MyDTBool_Bool_Bool_t gacZ_goMux_mux_d;
  logic gacZ_goMux_mux_r;
  MyBool_t \v'ad0_goMux_mux_d ;
  logic \v'ad0_goMux_mux_r ;
  Pointer_QTree_Bool_t mad1_goMux_mux_d;
  logic mad1_goMux_mux_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  C2_t go_9_goMux_choice_1_d;
  logic go_9_goMux_choice_1_r;
  C2_t go_9_goMux_choice_2_d;
  logic go_9_goMux_choice_2_r;
  Pointer_Nat_t xadg_goMux_mux_d;
  logic xadg_goMux_mux_r;
  Pointer_Nat_t yadh_goMux_mux_d;
  logic yadh_goMux_mux_r;
  MyDTNat_Bool_t isZacQ_2_2_argbuf_d;
  logic isZacQ_2_2_argbuf_r;
  MyDTNat_Bool_t isZacQ_2_1_d;
  logic isZacQ_2_1_r;
  MyDTNat_Bool_t isZacQ_2_2_d;
  logic isZacQ_2_2_r;
  MyDTNat_Bool_t isZacQ_3_2_argbuf_d;
  logic isZacQ_3_2_argbuf_r;
  MyDTNat_Bool_t isZacQ_3_1_d;
  logic isZacQ_3_1_r;
  MyDTNat_Bool_t isZacQ_3_2_d;
  logic isZacQ_3_2_r;
  MyDTNat_Bool_t isZacQ_4_1_argbuf_d;
  logic isZacQ_4_1_argbuf_r;
  MyDTBool_Bool_t isZacY_2_2_argbuf_d;
  logic isZacY_2_2_argbuf_r;
  MyDTBool_Bool_t isZacY_2_1_d;
  logic isZacY_2_1_r;
  MyDTBool_Bool_t isZacY_2_2_d;
  logic isZacY_2_2_r;
  MyDTBool_Bool_t isZacY_3_2_argbuf_d;
  logic isZacY_3_2_argbuf_r;
  MyDTBool_Bool_t isZacY_3_1_d;
  logic isZacY_3_1_r;
  MyDTBool_Bool_t isZacY_3_2_d;
  logic isZacY_3_2_r;
  MyDTBool_Bool_t isZacY_4_1_argbuf_d;
  logic isZacY_4_1_argbuf_r;
  MyDTBool_Bool_t isZad7_2_2_argbuf_d;
  logic isZad7_2_2_argbuf_r;
  MyDTBool_Bool_t isZad7_2_1_d;
  logic isZad7_2_1_r;
  MyDTBool_Bool_t isZad7_2_2_d;
  logic isZad7_2_2_r;
  MyDTBool_Bool_t isZad7_3_2_argbuf_d;
  logic isZad7_3_2_argbuf_r;
  MyDTBool_Bool_t isZad7_3_1_d;
  logic isZad7_3_1_r;
  MyDTBool_Bool_t isZad7_3_2_d;
  logic isZad7_3_2_r;
  MyDTBool_Bool_t isZad7_4_1_argbuf_d;
  logic isZad7_4_1_argbuf_r;
  Go_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_r;
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_r;
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_r;
  MyDTBool_Bool_Bool_t gad8_1_1_argbuf_d;
  logic gad8_1_1_argbuf_r;
  Go_t go_10_1_d;
  logic go_10_1_r;
  Go_t go_10_2_d;
  logic go_10_2_r;
  MyDTBool_Bool_t isZad7_1_1_argbuf_d;
  logic isZad7_1_1_argbuf_r;
  Pointer_QTree_Bool_t m1ad9_1_1_argbuf_d;
  logic m1ad9_1_1_argbuf_r;
  Pointer_QTree_Bool_t m2ada_1_1_argbuf_d;
  logic m2ada_1_1_argbuf_r;
  Pointer_QTree_Bool_t es_2_1_argbuf_d;
  logic es_2_1_argbuf_r;
  Nat_t lizzieLet40_1_argbuf_d;
  logic lizzieLet40_1_argbuf_r;
  Pointer_QTree_Bool_t q1ad3_destruct_d;
  logic q1ad3_destruct_r;
  Pointer_QTree_Bool_t q2ad4_destruct_d;
  logic q2ad4_destruct_r;
  Pointer_QTree_Bool_t q3ad5_destruct_d;
  logic q3ad5_destruct_r;
  Pointer_QTree_Bool_t q4ad6_destruct_d;
  logic q4ad6_destruct_r;
  MyBool_t vad2_destruct_d;
  logic vad2_destruct_r;
  QTree_Bool_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  QTree_Bool_t lizzieLet12_1_1QVal_Bool_d;
  logic lizzieLet12_1_1QVal_Bool_r;
  QTree_Bool_t lizzieLet12_1_1QNode_Bool_d;
  logic lizzieLet12_1_1QNode_Bool_r;
  QTree_Bool_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTBool_Bool_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QVal_Bool_d;
  logic lizzieLet12_1_3QVal_Bool_r;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_d;
  logic lizzieLet12_1_3QNode_Bool_r;
  MyDTBool_Bool_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_1_d;
  logic lizzieLet12_1_3QNode_Bool_1_r;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_2_d;
  logic lizzieLet12_1_3QNode_Bool_2_r;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_2_argbuf_d;
  logic lizzieLet12_1_3QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QVal_Bool_1_argbuf_d;
  logic lizzieLet12_1_3QVal_Bool_1_argbuf_r;
  Go_t lizzieLet12_1_4QNone_Bool_d;
  logic lizzieLet12_1_4QNone_Bool_r;
  Go_t lizzieLet12_1_4QVal_Bool_d;
  logic lizzieLet12_1_4QVal_Bool_r;
  Go_t lizzieLet12_1_4QNode_Bool_d;
  logic lizzieLet12_1_4QNode_Bool_r;
  Go_t lizzieLet12_1_4QError_Bool_d;
  logic lizzieLet12_1_4QError_Bool_r;
  Go_t lizzieLet12_1_4QError_Bool_1_d;
  logic lizzieLet12_1_4QError_Bool_1_r;
  Go_t lizzieLet12_1_4QError_Bool_2_d;
  logic lizzieLet12_1_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet12_1_4QError_Bool_1QError_Bool_d;
  logic lizzieLet12_1_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t lizzieLet12_1_4QError_Bool_2_argbuf_d;
  logic lizzieLet12_1_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet12_1_4QNode_Bool_1_argbuf_d;
  logic lizzieLet12_1_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet12_1_4QNone_Bool_1_d;
  logic lizzieLet12_1_4QNone_Bool_1_r;
  Go_t lizzieLet12_1_4QNone_Bool_2_d;
  logic lizzieLet12_1_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet12_1_4QNone_Bool_1QNone_Bool_d;
  logic lizzieLet12_1_4QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet13_1_1_argbuf_d;
  logic lizzieLet13_1_1_argbuf_r;
  Go_t lizzieLet12_1_4QNone_Bool_2_argbuf_d;
  logic lizzieLet12_1_4QNone_Bool_2_argbuf_r;
  C5_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t lizzieLet12_1_4QVal_Bool_1_d;
  logic lizzieLet12_1_4QVal_Bool_1_r;
  Go_t lizzieLet12_1_4QVal_Bool_2_d;
  logic lizzieLet12_1_4QVal_Bool_2_r;
  Go_t lizzieLet12_1_4QVal_Bool_3_d;
  logic lizzieLet12_1_4QVal_Bool_3_r;
  Go_t lizzieLet12_1_4QVal_Bool_1_argbuf_d;
  logic lizzieLet12_1_4QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_t applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d;
  logic applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r;
  Go_t lizzieLet12_1_4QVal_Bool_2_argbuf_d;
  logic lizzieLet12_1_4QVal_Bool_2_argbuf_r;
  TupGo___MyDTBool_Bool___MyBool_t applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d;
  logic applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r;
  MyDTBool_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  MyDTBool_Bool_t lizzieLet12_1_5QVal_Bool_d;
  logic lizzieLet12_1_5QVal_Bool_r;
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_d;
  logic lizzieLet12_1_5QNode_Bool_r;
  MyDTBool_Bool_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_1_d;
  logic lizzieLet12_1_5QNode_Bool_1_r;
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_2_d;
  logic lizzieLet12_1_5QNode_Bool_2_r;
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_2_argbuf_d;
  logic lizzieLet12_1_5QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_t lizzieLet12_1_5QVal_Bool_1_argbuf_d;
  logic lizzieLet12_1_5QVal_Bool_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QNone_Bool_d;
  logic lizzieLet12_1_6QNone_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QVal_Bool_d;
  logic lizzieLet12_1_6QVal_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QNode_Bool_d;
  logic lizzieLet12_1_6QNode_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QError_Bool_d;
  logic lizzieLet12_1_6QError_Bool_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QError_Bool_1_argbuf_d;
  logic lizzieLet12_1_6QError_Bool_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QNone_Bool_1_argbuf_d;
  logic lizzieLet12_1_6QNone_Bool_1_argbuf_r;
  MyBool_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  MyBool_t lizzieLet12_1_7QVal_Bool_d;
  logic lizzieLet12_1_7QVal_Bool_r;
  MyBool_t lizzieLet12_1_7QNode_Bool_d;
  logic lizzieLet12_1_7QNode_Bool_r;
  MyBool_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  MyBool_t lizzieLet12_1_7QNode_Bool_1_d;
  logic lizzieLet12_1_7QNode_Bool_1_r;
  MyBool_t lizzieLet12_1_7QNode_Bool_2_d;
  logic lizzieLet12_1_7QNode_Bool_2_r;
  MyBool_t lizzieLet12_1_7QNode_Bool_2_argbuf_d;
  logic lizzieLet12_1_7QNode_Bool_2_argbuf_r;
  MyBool_t lizzieLet12_1_7QVal_Bool_1_argbuf_d;
  logic lizzieLet12_1_7QVal_Bool_1_argbuf_r;
  Pointer_Nat_t x1adj_destruct_d;
  logic x1adj_destruct_r;
  Nat_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  Nat_t lizzieLet18_1Succ_d;
  logic lizzieLet18_1Succ_r;
  Go_t lizzieLet18_3Zero_d;
  logic lizzieLet18_3Zero_r;
  Go_t lizzieLet18_3Succ_d;
  logic lizzieLet18_3Succ_r;
  Nat_t lizzieLet18_4Zero_d;
  logic lizzieLet18_4Zero_r;
  Nat_t lizzieLet18_4Succ_d;
  logic lizzieLet18_4Succ_r;
  Nat_t lizzieLet18_4Succ_1_d;
  logic lizzieLet18_4Succ_1_r;
  Nat_t lizzieLet18_4Succ_2_d;
  logic lizzieLet18_4Succ_2_r;
  Nat_t lizzieLet18_4Succ_3_d;
  logic lizzieLet18_4Succ_3_r;
  Nat_t lizzieLet18_4Succ_4_d;
  logic lizzieLet18_4Succ_4_r;
  Pointer_Nat_t y1adk_destruct_d;
  logic y1adk_destruct_r;
  Nat_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  Nat_t lizzieLet18_4Succ_1Succ_d;
  logic lizzieLet18_4Succ_1Succ_r;
  Go_t lizzieLet18_4Succ_3Zero_d;
  logic lizzieLet18_4Succ_3Zero_r;
  Go_t lizzieLet18_4Succ_3Succ_d;
  logic lizzieLet18_4Succ_3Succ_r;
  Go_t lizzieLet18_4Succ_3Succ_1_argbuf_d;
  logic lizzieLet18_4Succ_3Succ_1_argbuf_r;
  MyBool_t lizzieLet18_4Succ_3Zero_1MyFalse_d;
  logic lizzieLet18_4Succ_3Zero_1MyFalse_r;
  Pointer_Nat_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  Pointer_Nat_t lizzieLet18_4Succ_4Succ_d;
  logic lizzieLet18_4Succ_4Succ_r;
  Pointer_Nat_t lizzieLet18_4Succ_4Succ_1_argbuf_d;
  logic lizzieLet18_4Succ_4Succ_1_argbuf_r;
  Go_t lizzieLet18_4Zero_1Zero_d;
  logic lizzieLet18_4Zero_1Zero_r;
  Go_t lizzieLet18_4Zero_1Succ_d;
  logic lizzieLet18_4Zero_1Succ_r;
  MyBool_t lizzieLet18_4Zero_1Succ_1MyFalse_d;
  logic lizzieLet18_4Zero_1Succ_1MyFalse_r;
  MyBool_t lizzieLet18_4Zero_1Zero_1MyTrue_d;
  logic lizzieLet18_4Zero_1Zero_1MyTrue_r;
  MyBool_t lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d;
  logic lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_r;
  MyBool_t lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d;
  logic lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_r;
  MyBool_t lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_d;
  logic lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_r;
  MyBool_t lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d;
  logic lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_r;
  Go_t eqNat_goConst_d;
  logic eqNat_goConst_r;
  Pointer_QTree_Bool_t es_1_2_destruct_d;
  logic es_1_2_destruct_r;
  Pointer_QTree_Bool_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Bool_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  Pointer_QTree_Bool_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Bool_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  MyDTBool_Bool_t isZad7_4_destruct_d;
  logic isZad7_4_destruct_r;
  MyDTBool_Bool_Bool_t gad8_4_destruct_d;
  logic gad8_4_destruct_r;
  Pointer_QTree_Bool_t q1adc_3_destruct_d;
  logic q1adc_3_destruct_r;
  Pointer_QTree_Bool_t m2ada_4_destruct_d;
  logic m2ada_4_destruct_r;
  Pointer_QTree_Bool_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  MyDTBool_Bool_t isZad7_3_destruct_d;
  logic isZad7_3_destruct_r;
  MyDTBool_Bool_Bool_t gad8_3_destruct_d;
  logic gad8_3_destruct_r;
  Pointer_QTree_Bool_t q1adc_2_destruct_d;
  logic q1adc_2_destruct_r;
  Pointer_QTree_Bool_t m2ada_3_destruct_d;
  logic m2ada_3_destruct_r;
  Pointer_QTree_Bool_t q2add_2_destruct_d;
  logic q2add_2_destruct_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  MyDTBool_Bool_t isZad7_2_destruct_d;
  logic isZad7_2_destruct_r;
  MyDTBool_Bool_Bool_t gad8_2_destruct_d;
  logic gad8_2_destruct_r;
  Pointer_QTree_Bool_t q1adc_1_destruct_d;
  logic q1adc_1_destruct_r;
  Pointer_QTree_Bool_t m2ada_2_destruct_d;
  logic m2ada_2_destruct_r;
  Pointer_QTree_Bool_t q2add_1_destruct_d;
  logic q2add_1_destruct_r;
  Pointer_QTree_Bool_t q3ade_1_destruct_d;
  logic q3ade_1_destruct_r;
  CTkron_kron_Bool_Bool_Bool_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_r;
  Go_t _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d;
  logic lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_r;
  QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r;
  QTree_Bool_t lizzieLet28_1_argbuf_d;
  logic lizzieLet28_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d;
  logic lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Bool_t lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d;
  logic lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r;
  Go_t call_kron_kron_Bool_Bool_Bool_goConst_d;
  logic call_kron_kron_Bool_Bool_Bool_goConst_r;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_d;
  logic kron_kron_Bool_Bool_Bool_resbuf_r;
  Pointer_QTree_Nat_t es_2_3_destruct_d;
  logic es_2_3_destruct_r;
  Pointer_QTree_Nat_t es_3_5_destruct_d;
  logic es_3_5_destruct_r;
  Pointer_QTree_Nat_t es_4_3_destruct_d;
  logic es_4_3_destruct_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Nat_t es_3_4_destruct_d;
  logic es_3_4_destruct_r;
  Pointer_QTree_Nat_t es_4_2_destruct_d;
  logic es_4_2_destruct_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  MyDTNat_Bool_t isZacQ_4_destruct_d;
  logic isZacQ_4_destruct_r;
  MyDTBool_Nat_t gacR_4_destruct_d;
  logic gacR_4_destruct_r;
  Pointer_QTree_Bool_t q1acU_3_destruct_d;
  logic q1acU_3_destruct_r;
  Pointer_QTree_Nat_t es_4_1_destruct_d;
  logic es_4_1_destruct_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  MyDTNat_Bool_t isZacQ_3_destruct_d;
  logic isZacQ_3_destruct_r;
  MyDTBool_Nat_t gacR_3_destruct_d;
  logic gacR_3_destruct_r;
  Pointer_QTree_Bool_t q1acU_2_destruct_d;
  logic q1acU_2_destruct_r;
  Pointer_QTree_Bool_t q2acV_2_destruct_d;
  logic q2acV_2_destruct_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  MyDTNat_Bool_t isZacQ_2_destruct_d;
  logic isZacQ_2_destruct_r;
  MyDTBool_Nat_t gacR_2_destruct_d;
  logic gacR_2_destruct_r;
  Pointer_QTree_Bool_t q1acU_1_destruct_d;
  logic q1acU_1_destruct_r;
  Pointer_QTree_Bool_t q2acV_1_destruct_d;
  logic q2acV_1_destruct_r;
  Pointer_QTree_Bool_t q3acW_1_destruct_d;
  logic q3acW_1_destruct_r;
  \CTmain_map'_Bool_Nat_t  _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_1Lcall_main_map'_Bool_Nat3_d ;
  logic \lizzieLet29_1Lcall_main_map'_Bool_Nat3_r ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_1Lcall_main_map'_Bool_Nat2_d ;
  logic \lizzieLet29_1Lcall_main_map'_Bool_Nat2_r ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_1Lcall_main_map'_Bool_Nat1_d ;
  logic \lizzieLet29_1Lcall_main_map'_Bool_Nat1_r ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_1Lcall_main_map'_Bool_Nat0_d ;
  logic \lizzieLet29_1Lcall_main_map'_Bool_Nat0_r ;
  Go_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat3_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat3_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat2_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat2_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat1_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat1_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat0_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat0_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_r ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lmain_map'_Bool_Natsbos_d ;
  logic \lizzieLet29_4Lmain_map'_Bool_Natsbos_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat3_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat3_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat2_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat2_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat1_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat1_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat0_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat0_r ;
  QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_r ;
  QTree_Nat_t lizzieLet33_1_argbuf_d;
  logic lizzieLet33_1_argbuf_r;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  Pointer_QTree_Nat_t \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_r ;
  Go_t \call_main_map'_Bool_Nat_goConst_d ;
  logic \call_main_map'_Bool_Nat_goConst_r ;
  Pointer_QTree_Nat_t \main_map'_Bool_Nat_resbuf_d ;
  logic \main_map'_Bool_Nat_resbuf_r ;
  Pointer_QTree_Bool_t q1adc_destruct_d;
  logic q1adc_destruct_r;
  Pointer_QTree_Bool_t q2add_destruct_d;
  logic q2add_destruct_r;
  Pointer_QTree_Bool_t q3ade_destruct_d;
  logic q3ade_destruct_r;
  Pointer_QTree_Bool_t q4adf_destruct_d;
  logic q4adf_destruct_r;
  MyBool_t vadb_destruct_d;
  logic vadb_destruct_r;
  QTree_Bool_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  QTree_Bool_t lizzieLet2_1QVal_Bool_d;
  logic lizzieLet2_1QVal_Bool_r;
  QTree_Bool_t lizzieLet2_1QNode_Bool_d;
  logic lizzieLet2_1QNode_Bool_r;
  QTree_Bool_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  MyDTBool_Bool_Bool_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet2_3QVal_Bool_d;
  logic lizzieLet2_3QVal_Bool_r;
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_d;
  logic lizzieLet2_3QNode_Bool_r;
  MyDTBool_Bool_Bool_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_1_d;
  logic lizzieLet2_3QNode_Bool_1_r;
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_2_d;
  logic lizzieLet2_3QNode_Bool_2_r;
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_2_argbuf_d;
  logic lizzieLet2_3QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_Bool_t lizzieLet2_3QVal_Bool_1_argbuf_d;
  logic lizzieLet2_3QVal_Bool_1_argbuf_r;
  Go_t lizzieLet2_4QNone_Bool_d;
  logic lizzieLet2_4QNone_Bool_r;
  Go_t lizzieLet2_4QVal_Bool_d;
  logic lizzieLet2_4QVal_Bool_r;
  Go_t lizzieLet2_4QNode_Bool_d;
  logic lizzieLet2_4QNode_Bool_r;
  Go_t lizzieLet2_4QError_Bool_d;
  logic lizzieLet2_4QError_Bool_r;
  Go_t lizzieLet2_4QError_Bool_1_d;
  logic lizzieLet2_4QError_Bool_1_r;
  Go_t lizzieLet2_4QError_Bool_2_d;
  logic lizzieLet2_4QError_Bool_2_r;
  QTree_Bool_t lizzieLet2_4QError_Bool_1QError_Bool_d;
  logic lizzieLet2_4QError_Bool_1QError_Bool_r;
  QTree_Bool_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Go_t lizzieLet2_4QError_Bool_2_argbuf_d;
  logic lizzieLet2_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet2_4QNode_Bool_1_argbuf_d;
  logic lizzieLet2_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet2_4QNone_Bool_1_d;
  logic lizzieLet2_4QNone_Bool_1_r;
  Go_t lizzieLet2_4QNone_Bool_2_d;
  logic lizzieLet2_4QNone_Bool_2_r;
  QTree_Bool_t lizzieLet2_4QNone_Bool_1QNone_Bool_d;
  logic lizzieLet2_4QNone_Bool_1QNone_Bool_r;
  QTree_Bool_t lizzieLet3_1_argbuf_d;
  logic lizzieLet3_1_argbuf_r;
  Go_t lizzieLet2_4QNone_Bool_2_argbuf_d;
  logic lizzieLet2_4QNone_Bool_2_argbuf_r;
  C4_t go_13_goMux_choice_d;
  logic go_13_goMux_choice_r;
  Go_t go_13_goMux_data_d;
  logic go_13_goMux_data_r;
  Go_t lizzieLet2_4QVal_Bool_1_d;
  logic lizzieLet2_4QVal_Bool_1_r;
  Go_t lizzieLet2_4QVal_Bool_2_d;
  logic lizzieLet2_4QVal_Bool_2_r;
  Go_t lizzieLet2_4QVal_Bool_1_argbuf_d;
  logic lizzieLet2_4QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r ;
  Go_t lizzieLet2_4QVal_Bool_2_argbuf_d;
  logic lizzieLet2_4QVal_Bool_2_argbuf_r;
  MyDTBool_Bool_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  MyDTBool_Bool_t lizzieLet2_5QVal_Bool_d;
  logic lizzieLet2_5QVal_Bool_r;
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_d;
  logic lizzieLet2_5QNode_Bool_r;
  MyDTBool_Bool_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_1_d;
  logic lizzieLet2_5QNode_Bool_1_r;
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_2_d;
  logic lizzieLet2_5QNode_Bool_2_r;
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_2_argbuf_d;
  logic lizzieLet2_5QNode_Bool_2_argbuf_r;
  MyDTBool_Bool_t lizzieLet2_5QVal_Bool_1_argbuf_d;
  logic lizzieLet2_5QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet2_6QVal_Bool_d;
  logic lizzieLet2_6QVal_Bool_r;
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_d;
  logic lizzieLet2_6QNode_Bool_r;
  Pointer_QTree_Bool_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_1_d;
  logic lizzieLet2_6QNode_Bool_1_r;
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_2_d;
  logic lizzieLet2_6QNode_Bool_2_r;
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_2_argbuf_d;
  logic lizzieLet2_6QNode_Bool_2_argbuf_r;
  Pointer_QTree_Bool_t lizzieLet2_6QVal_Bool_1_argbuf_d;
  logic lizzieLet2_6QVal_Bool_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNone_Bool_d;
  logic lizzieLet2_7QNone_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QVal_Bool_d;
  logic lizzieLet2_7QVal_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNode_Bool_d;
  logic lizzieLet2_7QNode_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QError_Bool_d;
  logic lizzieLet2_7QError_Bool_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QError_Bool_1_argbuf_d;
  logic lizzieLet2_7QError_Bool_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  logic lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet4_1_argbuf_d;
  logic lizzieLet4_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNone_Bool_1_argbuf_d;
  logic lizzieLet2_7QNone_Bool_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QVal_Bool_1_argbuf_d;
  logic lizzieLet2_7QVal_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t es_2_4_destruct_d;
  logic es_2_4_destruct_r;
  Pointer_QTree_Bool_t es_3_7_destruct_d;
  logic es_3_7_destruct_r;
  Pointer_QTree_Bool_t es_4_6_destruct_d;
  logic es_4_6_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Bool_t es_3_6_destruct_d;
  logic es_3_6_destruct_r;
  Pointer_QTree_Bool_t es_4_5_destruct_d;
  logic es_4_5_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  MyDTBool_Bool_t isZacY_4_destruct_d;
  logic isZacY_4_destruct_r;
  MyDTBool_Bool_Bool_t gacZ_4_destruct_d;
  logic gacZ_4_destruct_r;
  MyBool_t \v'ad0_4_destruct_d ;
  logic \v'ad0_4_destruct_r ;
  Pointer_QTree_Bool_t q1ad3_3_destruct_d;
  logic q1ad3_3_destruct_r;
  Pointer_QTree_Bool_t es_4_4_destruct_d;
  logic es_4_4_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  MyDTBool_Bool_t isZacY_3_destruct_d;
  logic isZacY_3_destruct_r;
  MyDTBool_Bool_Bool_t gacZ_3_destruct_d;
  logic gacZ_3_destruct_r;
  MyBool_t \v'ad0_3_destruct_d ;
  logic \v'ad0_3_destruct_r ;
  Pointer_QTree_Bool_t q1ad3_2_destruct_d;
  logic q1ad3_2_destruct_r;
  Pointer_QTree_Bool_t q2ad4_2_destruct_d;
  logic q2ad4_2_destruct_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  MyDTBool_Bool_t isZacY_2_destruct_d;
  logic isZacY_2_destruct_r;
  MyDTBool_Bool_Bool_t gacZ_2_destruct_d;
  logic gacZ_2_destruct_r;
  MyBool_t \v'ad0_2_destruct_d ;
  logic \v'ad0_2_destruct_r ;
  Pointer_QTree_Bool_t q1ad3_1_destruct_d;
  logic q1ad3_1_destruct_r;
  Pointer_QTree_Bool_t q2ad4_1_destruct_d;
  logic q2ad4_1_destruct_r;
  Pointer_QTree_Bool_t q3ad5_1_destruct_d;
  logic q3ad5_1_destruct_r;
  \CTmap''_map''_Bool_Bool_Bool_t  _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_r ;
  Go_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d ;
  logic \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_r ;
  QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_r ;
  QTree_Bool_t lizzieLet38_1_argbuf_d;
  logic lizzieLet38_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet37_1_argbuf_d;
  logic lizzieLet37_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet36_1_argbuf_d;
  logic lizzieLet36_1_argbuf_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet35_1_argbuf_d;
  logic lizzieLet35_1_argbuf_r;
  Pointer_QTree_Bool_t \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r ;
  Go_t \call_map''_map''_Bool_Bool_Bool_goConst_d ;
  logic \call_map''_map''_Bool_Bool_Bool_goConst_r ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_d ;
  logic \map''_map''_Bool_Bool_Bool_resbuf_r ;
  Pointer_QTree_Bool_t q1acU_destruct_d;
  logic q1acU_destruct_r;
  Pointer_QTree_Bool_t q2acV_destruct_d;
  logic q2acV_destruct_r;
  Pointer_QTree_Bool_t q3acW_destruct_d;
  logic q3acW_destruct_r;
  Pointer_QTree_Bool_t q4acX_destruct_d;
  logic q4acX_destruct_r;
  MyBool_t vacT_destruct_d;
  logic vacT_destruct_r;
  QTree_Bool_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  QTree_Bool_t lizzieLet6_1QVal_Bool_d;
  logic lizzieLet6_1QVal_Bool_r;
  QTree_Bool_t lizzieLet6_1QNode_Bool_d;
  logic lizzieLet6_1QNode_Bool_r;
  QTree_Bool_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  MyDTBool_Nat_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTBool_Nat_t lizzieLet6_3QVal_Bool_d;
  logic lizzieLet6_3QVal_Bool_r;
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_d;
  logic lizzieLet6_3QNode_Bool_r;
  MyDTBool_Nat_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_1_d;
  logic lizzieLet6_3QNode_Bool_1_r;
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_2_d;
  logic lizzieLet6_3QNode_Bool_2_r;
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_2_argbuf_d;
  logic lizzieLet6_3QNode_Bool_2_argbuf_r;
  MyDTBool_Nat_t lizzieLet6_3QVal_Bool_1_argbuf_d;
  logic lizzieLet6_3QVal_Bool_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Bool_d;
  logic lizzieLet6_4QNone_Bool_r;
  Go_t lizzieLet6_4QVal_Bool_d;
  logic lizzieLet6_4QVal_Bool_r;
  Go_t lizzieLet6_4QNode_Bool_d;
  logic lizzieLet6_4QNode_Bool_r;
  Go_t lizzieLet6_4QError_Bool_d;
  logic lizzieLet6_4QError_Bool_r;
  Go_t lizzieLet6_4QError_Bool_1_d;
  logic lizzieLet6_4QError_Bool_1_r;
  Go_t lizzieLet6_4QError_Bool_2_d;
  logic lizzieLet6_4QError_Bool_2_r;
  QTree_Nat_t lizzieLet6_4QError_Bool_1QError_Nat_d;
  logic lizzieLet6_4QError_Bool_1QError_Nat_r;
  QTree_Nat_t lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet6_4QError_Bool_2_argbuf_d;
  logic lizzieLet6_4QError_Bool_2_argbuf_r;
  Go_t lizzieLet6_4QNode_Bool_1_argbuf_d;
  logic lizzieLet6_4QNode_Bool_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Bool_1_d;
  logic lizzieLet6_4QNone_Bool_1_r;
  Go_t lizzieLet6_4QNone_Bool_2_d;
  logic lizzieLet6_4QNone_Bool_2_r;
  QTree_Nat_t lizzieLet6_4QNone_Bool_1QNone_Nat_d;
  logic lizzieLet6_4QNone_Bool_1QNone_Nat_r;
  QTree_Nat_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Bool_2_argbuf_d;
  logic lizzieLet6_4QNone_Bool_2_argbuf_r;
  C5_t go_14_goMux_choice_d;
  logic go_14_goMux_choice_r;
  Go_t go_14_goMux_data_d;
  logic go_14_goMux_data_r;
  Go_t lizzieLet6_4QVal_Bool_1_d;
  logic lizzieLet6_4QVal_Bool_1_r;
  Go_t lizzieLet6_4QVal_Bool_2_d;
  logic lizzieLet6_4QVal_Bool_2_r;
  Go_t lizzieLet6_4QVal_Bool_3_d;
  logic lizzieLet6_4QVal_Bool_3_r;
  Go_t lizzieLet6_4QVal_Bool_1_argbuf_d;
  logic lizzieLet6_4QVal_Bool_1_argbuf_r;
  TupGo___MyDTBool_Nat___MyBool_t applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d;
  logic applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_r;
  Go_t lizzieLet6_4QVal_Bool_2_argbuf_d;
  logic lizzieLet6_4QVal_Bool_2_argbuf_r;
  TupGo___MyDTNat_Bool___Pointer_Nat_t applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d;
  logic applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_r;
  MyDTNat_Bool_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  MyDTNat_Bool_t lizzieLet6_5QVal_Bool_d;
  logic lizzieLet6_5QVal_Bool_r;
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_d;
  logic lizzieLet6_5QNode_Bool_r;
  MyDTNat_Bool_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_1_d;
  logic lizzieLet6_5QNode_Bool_1_r;
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_2_d;
  logic lizzieLet6_5QNode_Bool_2_r;
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_2_argbuf_d;
  logic lizzieLet6_5QNode_Bool_2_argbuf_r;
  MyDTNat_Bool_t lizzieLet6_5QVal_Bool_1_argbuf_d;
  logic lizzieLet6_5QVal_Bool_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QNone_Bool_d;
  logic lizzieLet6_6QNone_Bool_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QVal_Bool_d;
  logic lizzieLet6_6QVal_Bool_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QNode_Bool_d;
  logic lizzieLet6_6QNode_Bool_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QError_Bool_d;
  logic lizzieLet6_6QError_Bool_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QError_Bool_1_argbuf_d;
  logic lizzieLet6_6QError_Bool_1_argbuf_r;
  \CTmain_map'_Bool_Nat_t  \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_d ;
  logic \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QNone_Bool_1_argbuf_d;
  logic lizzieLet6_6QNone_Bool_1_argbuf_r;
  Pointer_QTree_Bool_t m1ad9_1_argbuf_d;
  logic m1ad9_1_argbuf_r;
  Pointer_QTree_Bool_t m2ada_2_2_argbuf_d;
  logic m2ada_2_2_argbuf_r;
  Pointer_QTree_Bool_t m2ada_2_1_d;
  logic m2ada_2_1_r;
  Pointer_QTree_Bool_t m2ada_2_2_d;
  logic m2ada_2_2_r;
  Pointer_QTree_Bool_t m2ada_3_2_argbuf_d;
  logic m2ada_3_2_argbuf_r;
  Pointer_QTree_Bool_t m2ada_3_1_d;
  logic m2ada_3_1_r;
  Pointer_QTree_Bool_t m2ada_3_2_d;
  logic m2ada_3_2_r;
  Pointer_QTree_Bool_t m2ada_4_1_argbuf_d;
  logic m2ada_4_1_argbuf_r;
  Pointer_QTree_Bool_t macS_1_argbuf_d;
  logic macS_1_argbuf_r;
  Pointer_QTree_Bool_t mad1_1_argbuf_d;
  logic mad1_1_argbuf_r;
  Go_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_r ;
  MyDTNat_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_r ;
  MyDTBool_Nat_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_r ;
  Pointer_QTree_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_r ;
  MyDTBool_Nat_t gacR_1_1_argbuf_d;
  logic gacR_1_1_argbuf_r;
  Go_t go_11_1_d;
  logic go_11_1_r;
  Go_t go_11_2_d;
  logic go_11_2_r;
  MyDTNat_Bool_t isZacQ_1_1_argbuf_d;
  logic isZacQ_1_1_argbuf_r;
  Pointer_QTree_Bool_t macS_1_1_argbuf_d;
  logic macS_1_1_argbuf_r;
  Go_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_r ;
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_r ;
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_r ;
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_r ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_r ;
  MyDTBool_Bool_Bool_t gacZ_1_1_argbuf_d;
  logic gacZ_1_1_argbuf_r;
  Go_t go_12_1_d;
  logic go_12_1_r;
  Go_t go_12_2_d;
  logic go_12_2_r;
  MyDTBool_Bool_t isZacY_1_1_argbuf_d;
  logic isZacY_1_1_argbuf_r;
  Pointer_QTree_Bool_t mad1_1_1_argbuf_d;
  logic mad1_1_1_argbuf_r;
  MyBool_t \v'ad0_1_1_argbuf_d ;
  logic \v'ad0_1_1_argbuf_r ;
  Pointer_QTree_Bool_t lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Pointer_QTree_Bool_t q1acU_3_1_argbuf_d;
  logic q1acU_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1ad3_3_1_argbuf_d;
  logic q1ad3_3_1_argbuf_r;
  Pointer_QTree_Bool_t q1adc_3_1_argbuf_d;
  logic q1adc_3_1_argbuf_r;
  Pointer_QTree_Bool_t q2acV_2_1_argbuf_d;
  logic q2acV_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2ad4_2_1_argbuf_d;
  logic q2ad4_2_1_argbuf_r;
  Pointer_QTree_Bool_t q2add_2_1_argbuf_d;
  logic q2add_2_1_argbuf_r;
  Pointer_QTree_Bool_t q3acW_1_1_argbuf_d;
  logic q3acW_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3ad5_1_1_argbuf_d;
  logic q3ad5_1_1_argbuf_r;
  Pointer_QTree_Bool_t q3ade_1_1_argbuf_d;
  logic q3ade_1_1_argbuf_r;
  Pointer_QTree_Bool_t q4acX_1_argbuf_d;
  logic q4acX_1_argbuf_r;
  Pointer_QTree_Bool_t q4ad6_1_argbuf_d;
  logic q4ad6_1_argbuf_r;
  Pointer_QTree_Bool_t q4adf_1_argbuf_d;
  logic q4adf_1_argbuf_r;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_1_d;
  logic lizzieLet24_1_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_2_d;
  logic lizzieLet24_2_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_3_d;
  logic lizzieLet24_3_r;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4_d;
  logic lizzieLet24_4_r;
  \CTmain_map'_Bool_Nat_t  \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_r ;
  \CTmain_map'_Bool_Nat_t  lizzieLet29_1_d;
  logic lizzieLet29_1_r;
  \CTmain_map'_Bool_Nat_t  lizzieLet29_2_d;
  logic lizzieLet29_2_r;
  \CTmain_map'_Bool_Nat_t  lizzieLet29_3_d;
  logic lizzieLet29_3_r;
  \CTmain_map'_Bool_Nat_t  lizzieLet29_4_d;
  logic lizzieLet29_4_r;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r ;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet34_1_d;
  logic lizzieLet34_1_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet34_2_d;
  logic lizzieLet34_2_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet34_3_d;
  logic lizzieLet34_3_r;
  \CTmap''_map''_Bool_Bool_Bool_t  lizzieLet34_4_d;
  logic lizzieLet34_4_r;
  Nat_t readPointer_Natxadg_1_argbuf_rwb_d;
  logic readPointer_Natxadg_1_argbuf_rwb_r;
  Nat_t lizzieLet18_1_d;
  logic lizzieLet18_1_r;
  Nat_t lizzieLet18_2_d;
  logic lizzieLet18_2_r;
  Nat_t lizzieLet18_3_d;
  logic lizzieLet18_3_r;
  Nat_t lizzieLet18_4_d;
  logic lizzieLet18_4_r;
  Nat_t readPointer_Natyadh_1_argbuf_rwb_d;
  logic readPointer_Natyadh_1_argbuf_rwb_r;
  QTree_Bool_t readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolm1ad9_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet2_1_d;
  logic lizzieLet2_1_r;
  QTree_Bool_t lizzieLet2_2_d;
  logic lizzieLet2_2_r;
  QTree_Bool_t lizzieLet2_3_d;
  logic lizzieLet2_3_r;
  QTree_Bool_t lizzieLet2_4_d;
  logic lizzieLet2_4_r;
  QTree_Bool_t lizzieLet2_5_d;
  logic lizzieLet2_5_r;
  QTree_Bool_t lizzieLet2_6_d;
  logic lizzieLet2_6_r;
  QTree_Bool_t lizzieLet2_7_d;
  logic lizzieLet2_7_r;
  QTree_Bool_t readPointer_QTree_BoolmacS_1_argbuf_rwb_d;
  logic readPointer_QTree_BoolmacS_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Bool_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Bool_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Bool_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Bool_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Bool_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Bool_t readPointer_QTree_Boolmad1_1_argbuf_rwb_d;
  logic readPointer_QTree_Boolmad1_1_argbuf_rwb_r;
  QTree_Bool_t lizzieLet12_1_1_d;
  logic lizzieLet12_1_1_r;
  QTree_Bool_t lizzieLet12_1_2_d;
  logic lizzieLet12_1_2_r;
  QTree_Bool_t lizzieLet12_1_3_d;
  logic lizzieLet12_1_3_r;
  QTree_Bool_t lizzieLet12_1_4_d;
  logic lizzieLet12_1_4_r;
  QTree_Bool_t lizzieLet12_1_5_d;
  logic lizzieLet12_1_5_r;
  QTree_Bool_t lizzieLet12_1_6_d;
  logic lizzieLet12_1_6_r;
  QTree_Bool_t lizzieLet12_1_7_d;
  logic lizzieLet12_1_7_r;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Go_t to_nat1TupGogo_16_d;
  logic to_nat1TupGogo_16_r;
  Nat_t go_16_1Zero_d;
  logic go_16_1Zero_r;
  MyBool_t \v'ad0_2_2_argbuf_d ;
  logic \v'ad0_2_2_argbuf_r ;
  MyBool_t \v'ad0_2_1_d ;
  logic \v'ad0_2_1_r ;
  MyBool_t \v'ad0_2_2_d ;
  logic \v'ad0_2_2_r ;
  MyBool_t \v'ad0_3_2_argbuf_d ;
  logic \v'ad0_3_2_argbuf_r ;
  MyBool_t \v'ad0_3_1_d ;
  logic \v'ad0_3_1_r ;
  MyBool_t \v'ad0_3_2_d ;
  logic \v'ad0_3_2_r ;
  MyBool_t \v'ad0_4_1_argbuf_d ;
  logic \v'ad0_4_1_argbuf_r ;
  MyBool_t vacT_1_argbuf_d;
  logic vacT_1_argbuf_r;
  MyBool_t vad2_1_argbuf_d;
  logic vad2_1_argbuf_r;
  MyBool_t vadb_1_argbuf_d;
  logic vadb_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet14_1_1_argbuf_d;
  logic lizzieLet14_1_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_r;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_r ;
  \Pointer_CTmain_map'_Bool_Nat_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_r ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_rwb_d;
  logic writeNatlizzieLet0_1_argbuf_rwb_r;
  Pointer_Nat_t applyfnBool_Nat_5_resbuf_d;
  logic applyfnBool_Nat_5_resbuf_r;
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_rwb_d;
  logic writeNatlizzieLet1_1_argbuf_rwb_r;
  Pointer_Nat_t es_1_1_1_argbuf_d;
  logic es_1_1_1_argbuf_r;
  Pointer_Nat_t writeNatlizzieLet39_1_argbuf_rwb_d;
  logic writeNatlizzieLet39_1_argbuf_rwb_r;
  Nat_t lizzieLet0_1_1Succ_d;
  logic lizzieLet0_1_1Succ_r;
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_rwb_d;
  logic writeNatlizzieLet40_1_argbuf_rwb_r;
  Pointer_Nat_t to_nat1_resbuf_d;
  logic to_nat1_resbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_r;
  Pointer_QTree_Bool_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_rwb_d;
  logic writeQTree_NatlizzieLet11_1_1_argbuf_rwb_r;
  Pointer_QTree_Nat_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_rwb_d;
  logic writeQTree_NatlizzieLet33_1_argbuf_rwb_r;
  Pointer_QTree_Nat_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_NatlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Nat_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_rwb_d;
  logic writeQTree_NatlizzieLet8_1_argbuf_rwb_r;
  Pointer_QTree_Nat_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_NatlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Nat_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_Nat_t xacw_1_argbuf_d;
  logic xacw_1_argbuf_r;
  MyBool_t xacw_1_1_argbuf_d;
  logic xacw_1_1_argbuf_r;
  Pointer_Nat_t xadg_1_argbuf_d;
  logic xadg_1_argbuf_r;
  Pointer_Nat_t y1adk_1_argbuf_d;
  logic y1adk_1_argbuf_r;
  Pointer_Nat_t yadh_1_argbuf_d;
  logic yadh_1_argbuf_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go_5,Go),
                                (go_6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go),
                                (go__11,Go),
                                (go__12,Go),
                                (go__13,Go),
                                (go__14,Go),
                                (go__15,Go),
                                (go__16,Go)] */
  logic [15:0] sourceGo_emitted;
  logic [15:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign go__11_d = (sourceGo_d[0] && (! sourceGo_emitted[10]));
  assign go__12_d = (sourceGo_d[0] && (! sourceGo_emitted[11]));
  assign go__13_d = (sourceGo_d[0] && (! sourceGo_emitted[12]));
  assign go__14_d = (sourceGo_d[0] && (! sourceGo_emitted[13]));
  assign go__15_d = (sourceGo_d[0] && (! sourceGo_emitted[14]));
  assign go__16_d = (sourceGo_d[0] && (! sourceGo_emitted[15]));
  assign sourceGo_done = (sourceGo_emitted | ({go__16_d[0],
                                               go__15_d[0],
                                               go__14_d[0],
                                               go__13_d[0],
                                               go__12_d[0],
                                               go__11_d[0],
                                               go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go_6_d[0],
                                               go_5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__16_r,
                                                             go__15_r,
                                                             go__14_r,
                                                             go__13_r,
                                                             go__12_r,
                                                             go__11_r,
                                                             go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go_6_r,
                                                             go_5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 16'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 16'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,Lit 0) : (go__7,Go) > (initHP_Nat,Word16#) */
  assign initHP_Nat_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_Nat_r;
  
  /* const (Ty Word16#,Lit 1) : (incrHP_Nat1,Go) > (incrHP_Nat,Word16#) */
  assign incrHP_Nat_d = {16'd1, incrHP_Nat1_d[0]};
  assign incrHP_Nat1_r = incrHP_Nat_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_Nat2,Go)] > (incrHP_mergeNat,Go) */
  logic [1:0] incrHP_mergeNat_selected;
  logic [1:0] incrHP_mergeNat_select;
  always_comb
    begin
      incrHP_mergeNat_selected = 2'd0;
      if ((| incrHP_mergeNat_select))
        incrHP_mergeNat_selected = incrHP_mergeNat_select;
      else
        if (go__8_d[0]) incrHP_mergeNat_selected[0] = 1'd1;
        else if (incrHP_Nat2_d[0]) incrHP_mergeNat_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeNat_select <= 2'd0;
    else
      incrHP_mergeNat_select <= (incrHP_mergeNat_r ? 2'd0 :
                                 incrHP_mergeNat_selected);
  always_comb
    if (incrHP_mergeNat_selected[0]) incrHP_mergeNat_d = go__8_d;
    else if (incrHP_mergeNat_selected[1])
      incrHP_mergeNat_d = incrHP_Nat2_d;
    else incrHP_mergeNat_d = 1'd0;
  assign {incrHP_Nat2_r,
          go__8_r} = (incrHP_mergeNat_r ? incrHP_mergeNat_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeNat_buf,Go) > [(incrHP_Nat1,Go),
                                           (incrHP_Nat2,Go)] */
  logic [1:0] incrHP_mergeNat_buf_emitted;
  logic [1:0] incrHP_mergeNat_buf_done;
  assign incrHP_Nat1_d = (incrHP_mergeNat_buf_d[0] && (! incrHP_mergeNat_buf_emitted[0]));
  assign incrHP_Nat2_d = (incrHP_mergeNat_buf_d[0] && (! incrHP_mergeNat_buf_emitted[1]));
  assign incrHP_mergeNat_buf_done = (incrHP_mergeNat_buf_emitted | ({incrHP_Nat2_d[0],
                                                                     incrHP_Nat1_d[0]} & {incrHP_Nat2_r,
                                                                                          incrHP_Nat1_r}));
  assign incrHP_mergeNat_buf_r = (& incrHP_mergeNat_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeNat_buf_emitted <= 2'd0;
    else
      incrHP_mergeNat_buf_emitted <= (incrHP_mergeNat_buf_r ? 2'd0 :
                                      incrHP_mergeNat_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_Nat,Word16#) (forkHP1_Nat,Word16#) > (addHP_Nat,Word16#) */
  assign addHP_Nat_d = {(incrHP_Nat_d[16:1] + forkHP1_Nat_d[16:1]),
                        (incrHP_Nat_d[0] && forkHP1_Nat_d[0])};
  assign {incrHP_Nat_r,
          forkHP1_Nat_r} = {2 {(addHP_Nat_r && addHP_Nat_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_Nat,Word16#),
                      (addHP_Nat,Word16#)] > (mergeHP_Nat,Word16#) */
  logic [1:0] mergeHP_Nat_selected;
  logic [1:0] mergeHP_Nat_select;
  always_comb
    begin
      mergeHP_Nat_selected = 2'd0;
      if ((| mergeHP_Nat_select))
        mergeHP_Nat_selected = mergeHP_Nat_select;
      else
        if (initHP_Nat_d[0]) mergeHP_Nat_selected[0] = 1'd1;
        else if (addHP_Nat_d[0]) mergeHP_Nat_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_Nat_select <= 2'd0;
    else
      mergeHP_Nat_select <= (mergeHP_Nat_r ? 2'd0 :
                             mergeHP_Nat_selected);
  always_comb
    if (mergeHP_Nat_selected[0]) mergeHP_Nat_d = initHP_Nat_d;
    else if (mergeHP_Nat_selected[1]) mergeHP_Nat_d = addHP_Nat_d;
    else mergeHP_Nat_d = {16'd0, 1'd0};
  assign {addHP_Nat_r,
          initHP_Nat_r} = (mergeHP_Nat_r ? mergeHP_Nat_selected :
                           2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeNat,Go) > (incrHP_mergeNat_buf,Go) */
  Go_t incrHP_mergeNat_bufchan_d;
  logic incrHP_mergeNat_bufchan_r;
  assign incrHP_mergeNat_r = ((! incrHP_mergeNat_bufchan_d[0]) || incrHP_mergeNat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeNat_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeNat_r)
        incrHP_mergeNat_bufchan_d <= incrHP_mergeNat_d;
  Go_t incrHP_mergeNat_bufchan_buf;
  assign incrHP_mergeNat_bufchan_r = (! incrHP_mergeNat_bufchan_buf[0]);
  assign incrHP_mergeNat_buf_d = (incrHP_mergeNat_bufchan_buf[0] ? incrHP_mergeNat_bufchan_buf :
                                  incrHP_mergeNat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeNat_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeNat_buf_r && incrHP_mergeNat_bufchan_buf[0]))
        incrHP_mergeNat_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeNat_buf_r) && (! incrHP_mergeNat_bufchan_buf[0])))
        incrHP_mergeNat_bufchan_buf <= incrHP_mergeNat_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_Nat,Word16#) > (mergeHP_Nat_buf,Word16#) */
  \Word16#_t  mergeHP_Nat_bufchan_d;
  logic mergeHP_Nat_bufchan_r;
  assign mergeHP_Nat_r = ((! mergeHP_Nat_bufchan_d[0]) || mergeHP_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_Nat_bufchan_d <= {16'd0, 1'd0};
    else if (mergeHP_Nat_r) mergeHP_Nat_bufchan_d <= mergeHP_Nat_d;
  \Word16#_t  mergeHP_Nat_bufchan_buf;
  assign mergeHP_Nat_bufchan_r = (! mergeHP_Nat_bufchan_buf[0]);
  assign mergeHP_Nat_buf_d = (mergeHP_Nat_bufchan_buf[0] ? mergeHP_Nat_bufchan_buf :
                              mergeHP_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_Nat_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_Nat_buf_r && mergeHP_Nat_bufchan_buf[0]))
        mergeHP_Nat_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_Nat_buf_r) && (! mergeHP_Nat_bufchan_buf[0])))
        mergeHP_Nat_bufchan_buf <= mergeHP_Nat_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_Nat_buf,Word16#) > [(forkHP1_Nat,Word16#),
                                                 (forkHP1_Na2,Word16#),
                                                 (forkHP1_Na3,Word16#)] */
  logic [2:0] mergeHP_Nat_buf_emitted;
  logic [2:0] mergeHP_Nat_buf_done;
  assign forkHP1_Nat_d = {mergeHP_Nat_buf_d[16:1],
                          (mergeHP_Nat_buf_d[0] && (! mergeHP_Nat_buf_emitted[0]))};
  assign forkHP1_Na2_d = {mergeHP_Nat_buf_d[16:1],
                          (mergeHP_Nat_buf_d[0] && (! mergeHP_Nat_buf_emitted[1]))};
  assign forkHP1_Na3_d = {mergeHP_Nat_buf_d[16:1],
                          (mergeHP_Nat_buf_d[0] && (! mergeHP_Nat_buf_emitted[2]))};
  assign mergeHP_Nat_buf_done = (mergeHP_Nat_buf_emitted | ({forkHP1_Na3_d[0],
                                                             forkHP1_Na2_d[0],
                                                             forkHP1_Nat_d[0]} & {forkHP1_Na3_r,
                                                                                  forkHP1_Na2_r,
                                                                                  forkHP1_Nat_r}));
  assign mergeHP_Nat_buf_r = (& mergeHP_Nat_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_Nat_buf_emitted <= 3'd0;
    else
      mergeHP_Nat_buf_emitted <= (mergeHP_Nat_buf_r ? 3'd0 :
                                  mergeHP_Nat_buf_done);
  
  /* mergectrl (Ty C2,Ty MemIn_Nat) : [(dconReadIn_Nat,MemIn_Nat),
                                  (dconWriteIn_Nat,MemIn_Nat)] > (memMergeChoice_Nat,C2) (memMergeIn_Nat,MemIn_Nat) */
  logic [1:0] dconReadIn_Nat_select_d;
  assign dconReadIn_Nat_select_d = ((| dconReadIn_Nat_select_q) ? dconReadIn_Nat_select_q :
                                    (dconReadIn_Nat_d[0] ? 2'd1 :
                                     (dconWriteIn_Nat_d[0] ? 2'd2 :
                                      2'd0)));
  logic [1:0] dconReadIn_Nat_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_Nat_select_q <= 2'd0;
    else
      dconReadIn_Nat_select_q <= (dconReadIn_Nat_done ? 2'd0 :
                                  dconReadIn_Nat_select_d);
  logic [1:0] dconReadIn_Nat_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_Nat_emit_q <= 2'd0;
    else
      dconReadIn_Nat_emit_q <= (dconReadIn_Nat_done ? 2'd0 :
                                dconReadIn_Nat_emit_d);
  logic [1:0] dconReadIn_Nat_emit_d;
  assign dconReadIn_Nat_emit_d = (dconReadIn_Nat_emit_q | ({memMergeChoice_Nat_d[0],
                                                            memMergeIn_Nat_d[0]} & {memMergeChoice_Nat_r,
                                                                                    memMergeIn_Nat_r}));
  logic dconReadIn_Nat_done;
  assign dconReadIn_Nat_done = (& dconReadIn_Nat_emit_d);
  assign {dconWriteIn_Nat_r,
          dconReadIn_Nat_r} = (dconReadIn_Nat_done ? dconReadIn_Nat_select_d :
                               2'd0);
  assign memMergeIn_Nat_d = ((dconReadIn_Nat_select_d[0] && (! dconReadIn_Nat_emit_q[0])) ? dconReadIn_Nat_d :
                             ((dconReadIn_Nat_select_d[1] && (! dconReadIn_Nat_emit_q[0])) ? dconWriteIn_Nat_d :
                              {34'd0, 1'd0}));
  assign memMergeChoice_Nat_d = ((dconReadIn_Nat_select_d[0] && (! dconReadIn_Nat_emit_q[1])) ? C1_2_dc(1'd1) :
                                 ((dconReadIn_Nat_select_d[1] && (! dconReadIn_Nat_emit_q[1])) ? C2_2_dc(1'd1) :
                                  {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_Nat,
      Ty MemOut_Nat) : (memMergeIn_Nat_dbuf,MemIn_Nat) > (memOut_Nat,MemOut_Nat) */
  logic [16:0] memMergeIn_Nat_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_Nat_dbuf_address;
  logic [16:0] memMergeIn_Nat_dbuf_din;
  logic [16:0] memOut_Nat_q;
  logic memOut_Nat_valid;
  logic memMergeIn_Nat_dbuf_we;
  logic memOut_Nat_we;
  assign memMergeIn_Nat_dbuf_din = memMergeIn_Nat_dbuf_d[34:18];
  assign memMergeIn_Nat_dbuf_address = memMergeIn_Nat_dbuf_d[17:2];
  assign memMergeIn_Nat_dbuf_we = (memMergeIn_Nat_dbuf_d[1:1] && memMergeIn_Nat_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_Nat_we <= 1'd0;
        memOut_Nat_valid <= 1'd0;
      end
    else
      begin
        memOut_Nat_we <= memMergeIn_Nat_dbuf_we;
        memOut_Nat_valid <= memMergeIn_Nat_dbuf_d[0];
        if (memMergeIn_Nat_dbuf_we)
          begin
            memMergeIn_Nat_dbuf_mem[memMergeIn_Nat_dbuf_address] <= memMergeIn_Nat_dbuf_din;
            memOut_Nat_q <= memMergeIn_Nat_dbuf_din;
          end
        else
          memOut_Nat_q <= memMergeIn_Nat_dbuf_mem[memMergeIn_Nat_dbuf_address];
      end
  assign memOut_Nat_d = {memOut_Nat_q,
                         memOut_Nat_we,
                         memOut_Nat_valid};
  assign memMergeIn_Nat_dbuf_r = ((! memOut_Nat_valid) || memOut_Nat_r);
  logic [31:0] profiling_MemIn_Nat_read;
  logic [31:0] profiling_MemIn_Nat_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_Nat_write <= 0;
        profiling_MemIn_Nat_read <= 0;
      end
    else
      if ((memMergeIn_Nat_dbuf_we == 1'd1))
        profiling_MemIn_Nat_write <= (profiling_MemIn_Nat_write + 1);
      else
        if ((memOut_Nat_valid == 1'd1))
          profiling_MemIn_Nat_read <= (profiling_MemIn_Nat_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_Nat) : (memMergeChoice_Nat,C2) (memOut_Nat_dbuf,MemOut_Nat) > [(memReadOut_Nat,MemOut_Nat),
                                                                                (memWriteOut_Nat,MemOut_Nat)] */
  logic [1:0] memOut_Nat_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_Nat_d[0] && memOut_Nat_dbuf_d[0]))
      unique case (memMergeChoice_Nat_d[1:1])
        1'd0: memOut_Nat_dbuf_onehotd = 2'd1;
        1'd1: memOut_Nat_dbuf_onehotd = 2'd2;
        default: memOut_Nat_dbuf_onehotd = 2'd0;
      endcase
    else memOut_Nat_dbuf_onehotd = 2'd0;
  assign memReadOut_Nat_d = {memOut_Nat_dbuf_d[18:1],
                             memOut_Nat_dbuf_onehotd[0]};
  assign memWriteOut_Nat_d = {memOut_Nat_dbuf_d[18:1],
                              memOut_Nat_dbuf_onehotd[1]};
  assign memOut_Nat_dbuf_r = (| (memOut_Nat_dbuf_onehotd & {memWriteOut_Nat_r,
                                                            memReadOut_Nat_r}));
  assign memMergeChoice_Nat_r = memOut_Nat_dbuf_r;
  
  /* dbuf (Ty MemIn_Nat) : (memMergeIn_Nat_rbuf,MemIn_Nat) > (memMergeIn_Nat_dbuf,MemIn_Nat) */
  assign memMergeIn_Nat_rbuf_r = ((! memMergeIn_Nat_dbuf_d[0]) || memMergeIn_Nat_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_Nat_dbuf_d <= {34'd0, 1'd0};
    else
      if (memMergeIn_Nat_rbuf_r)
        memMergeIn_Nat_dbuf_d <= memMergeIn_Nat_rbuf_d;
  
  /* rbuf (Ty MemIn_Nat) : (memMergeIn_Nat,MemIn_Nat) > (memMergeIn_Nat_rbuf,MemIn_Nat) */
  MemIn_Nat_t memMergeIn_Nat_buf;
  assign memMergeIn_Nat_r = (! memMergeIn_Nat_buf[0]);
  assign memMergeIn_Nat_rbuf_d = (memMergeIn_Nat_buf[0] ? memMergeIn_Nat_buf :
                                  memMergeIn_Nat_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_Nat_buf <= {34'd0, 1'd0};
    else
      if ((memMergeIn_Nat_rbuf_r && memMergeIn_Nat_buf[0]))
        memMergeIn_Nat_buf <= {34'd0, 1'd0};
      else if (((! memMergeIn_Nat_rbuf_r) && (! memMergeIn_Nat_buf[0])))
        memMergeIn_Nat_buf <= memMergeIn_Nat_d;
  
  /* dbuf (Ty MemOut_Nat) : (memOut_Nat_rbuf,MemOut_Nat) > (memOut_Nat_dbuf,MemOut_Nat) */
  assign memOut_Nat_rbuf_r = ((! memOut_Nat_dbuf_d[0]) || memOut_Nat_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_Nat_dbuf_d <= {18'd0, 1'd0};
    else if (memOut_Nat_rbuf_r) memOut_Nat_dbuf_d <= memOut_Nat_rbuf_d;
  
  /* rbuf (Ty MemOut_Nat) : (memOut_Nat,MemOut_Nat) > (memOut_Nat_rbuf,MemOut_Nat) */
  MemOut_Nat_t memOut_Nat_buf;
  assign memOut_Nat_r = (! memOut_Nat_buf[0]);
  assign memOut_Nat_rbuf_d = (memOut_Nat_buf[0] ? memOut_Nat_buf :
                              memOut_Nat_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_Nat_buf <= {18'd0, 1'd0};
    else
      if ((memOut_Nat_rbuf_r && memOut_Nat_buf[0]))
        memOut_Nat_buf <= {18'd0, 1'd0};
      else if (((! memOut_Nat_rbuf_r) && (! memOut_Nat_buf[0])))
        memOut_Nat_buf <= memOut_Nat_d;
  
  /* mergectrl (Ty C2,Ty Pointer_Nat) : [(xadg_1_argbuf,Pointer_Nat),
                                    (yadh_1_argbuf,Pointer_Nat)] > (readMerge_choice_Nat,C2) (readMerge_data_Nat,Pointer_Nat) */
  logic [1:0] xadg_1_argbuf_select_d;
  assign xadg_1_argbuf_select_d = ((| xadg_1_argbuf_select_q) ? xadg_1_argbuf_select_q :
                                   (xadg_1_argbuf_d[0] ? 2'd1 :
                                    (yadh_1_argbuf_d[0] ? 2'd2 :
                                     2'd0)));
  logic [1:0] xadg_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xadg_1_argbuf_select_q <= 2'd0;
    else
      xadg_1_argbuf_select_q <= (xadg_1_argbuf_done ? 2'd0 :
                                 xadg_1_argbuf_select_d);
  logic [1:0] xadg_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xadg_1_argbuf_emit_q <= 2'd0;
    else
      xadg_1_argbuf_emit_q <= (xadg_1_argbuf_done ? 2'd0 :
                               xadg_1_argbuf_emit_d);
  logic [1:0] xadg_1_argbuf_emit_d;
  assign xadg_1_argbuf_emit_d = (xadg_1_argbuf_emit_q | ({readMerge_choice_Nat_d[0],
                                                          readMerge_data_Nat_d[0]} & {readMerge_choice_Nat_r,
                                                                                      readMerge_data_Nat_r}));
  logic xadg_1_argbuf_done;
  assign xadg_1_argbuf_done = (& xadg_1_argbuf_emit_d);
  assign {yadh_1_argbuf_r,
          xadg_1_argbuf_r} = (xadg_1_argbuf_done ? xadg_1_argbuf_select_d :
                              2'd0);
  assign readMerge_data_Nat_d = ((xadg_1_argbuf_select_d[0] && (! xadg_1_argbuf_emit_q[0])) ? xadg_1_argbuf_d :
                                 ((xadg_1_argbuf_select_d[1] && (! xadg_1_argbuf_emit_q[0])) ? yadh_1_argbuf_d :
                                  {16'd0, 1'd0}));
  assign readMerge_choice_Nat_d = ((xadg_1_argbuf_select_d[0] && (! xadg_1_argbuf_emit_q[1])) ? C1_2_dc(1'd1) :
                                   ((xadg_1_argbuf_select_d[1] && (! xadg_1_argbuf_emit_q[1])) ? C2_2_dc(1'd1) :
                                    {1'd0, 1'd0}));
  
  /* demux (Ty C2,
       Ty Nat) : (readMerge_choice_Nat,C2) (destructReadOut_Nat,Nat) > [(readPointer_Natxadg_1_argbuf,Nat),
                                                                        (readPointer_Natyadh_1_argbuf,Nat)] */
  logic [1:0] destructReadOut_Nat_onehotd;
  always_comb
    if ((readMerge_choice_Nat_d[0] && destructReadOut_Nat_d[0]))
      unique case (readMerge_choice_Nat_d[1:1])
        1'd0: destructReadOut_Nat_onehotd = 2'd1;
        1'd1: destructReadOut_Nat_onehotd = 2'd2;
        default: destructReadOut_Nat_onehotd = 2'd0;
      endcase
    else destructReadOut_Nat_onehotd = 2'd0;
  assign readPointer_Natxadg_1_argbuf_d = {destructReadOut_Nat_d[17:1],
                                           destructReadOut_Nat_onehotd[0]};
  assign readPointer_Natyadh_1_argbuf_d = {destructReadOut_Nat_d[17:1],
                                           destructReadOut_Nat_onehotd[1]};
  assign destructReadOut_Nat_r = (| (destructReadOut_Nat_onehotd & {readPointer_Natyadh_1_argbuf_r,
                                                                    readPointer_Natxadg_1_argbuf_r}));
  assign readMerge_choice_Nat_r = destructReadOut_Nat_r;
  
  /* destruct (Ty Pointer_Nat,
          Dcon Pointer_Nat) : (readMerge_data_Nat,Pointer_Nat) > [(destructReadIn_Nat,Word16#)] */
  assign destructReadIn_Nat_d = {readMerge_data_Nat_d[16:1],
                                 readMerge_data_Nat_d[0]};
  assign readMerge_data_Nat_r = destructReadIn_Nat_r;
  
  /* dcon (Ty MemIn_Nat,
      Dcon ReadIn_Nat) : [(destructReadIn_Nat,Word16#)] > (dconReadIn_Nat,MemIn_Nat) */
  assign dconReadIn_Nat_d = ReadIn_Nat_dc((& {destructReadIn_Nat_d[0]}), destructReadIn_Nat_d);
  assign {destructReadIn_Nat_r} = {1 {(dconReadIn_Nat_r && dconReadIn_Nat_d[0])}};
  
  /* destruct (Ty MemOut_Nat,
          Dcon ReadOut_Nat) : (memReadOut_Nat,MemOut_Nat) > [(destructReadOut_Nat,Nat)] */
  assign destructReadOut_Nat_d = {memReadOut_Nat_d[18:2],
                                  memReadOut_Nat_d[0]};
  assign memReadOut_Nat_r = destructReadOut_Nat_r;
  
  /* mergectrl (Ty C4,Ty Nat) : [(lizzieLet0_1_argbuf,Nat),
                            (lizzieLet1_1_argbuf,Nat),
                            (lizzieLet39_1_argbuf,Nat),
                            (lizzieLet40_1_argbuf,Nat)] > (writeMerge_choice_Nat,C4) (writeMerge_data_Nat,Nat) */
  logic [3:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 4'd1 :
                                          (lizzieLet1_1_argbuf_d[0] ? 4'd2 :
                                           (lizzieLet39_1_argbuf_d[0] ? 4'd4 :
                                            (lizzieLet40_1_argbuf_d[0] ? 4'd8 :
                                             4'd0)))));
  logic [3:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 4'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 4'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_Nat_d[0],
                                                                      writeMerge_data_Nat_d[0]} & {writeMerge_choice_Nat_r,
                                                                                                   writeMerge_data_Nat_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet40_1_argbuf_r,
          lizzieLet39_1_argbuf_r,
          lizzieLet1_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    4'd0);
  assign writeMerge_data_Nat_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                  ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet1_1_argbuf_d :
                                   ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet39_1_argbuf_d :
                                    ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet40_1_argbuf_d :
                                     {17'd0, 1'd0}))));
  assign writeMerge_choice_Nat_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                    ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                     ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                      ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                       {2'd0, 1'd0}))));
  
  /* demux (Ty C4,
       Ty Pointer_Nat) : (writeMerge_choice_Nat,C4) (demuxWriteResult_Nat,Pointer_Nat) > [(writeNatlizzieLet0_1_argbuf,Pointer_Nat),
                                                                                          (writeNatlizzieLet1_1_argbuf,Pointer_Nat),
                                                                                          (writeNatlizzieLet39_1_argbuf,Pointer_Nat),
                                                                                          (writeNatlizzieLet40_1_argbuf,Pointer_Nat)] */
  logic [3:0] demuxWriteResult_Nat_onehotd;
  always_comb
    if ((writeMerge_choice_Nat_d[0] && demuxWriteResult_Nat_d[0]))
      unique case (writeMerge_choice_Nat_d[2:1])
        2'd0: demuxWriteResult_Nat_onehotd = 4'd1;
        2'd1: demuxWriteResult_Nat_onehotd = 4'd2;
        2'd2: demuxWriteResult_Nat_onehotd = 4'd4;
        2'd3: demuxWriteResult_Nat_onehotd = 4'd8;
        default: demuxWriteResult_Nat_onehotd = 4'd0;
      endcase
    else demuxWriteResult_Nat_onehotd = 4'd0;
  assign writeNatlizzieLet0_1_argbuf_d = {demuxWriteResult_Nat_d[16:1],
                                          demuxWriteResult_Nat_onehotd[0]};
  assign writeNatlizzieLet1_1_argbuf_d = {demuxWriteResult_Nat_d[16:1],
                                          demuxWriteResult_Nat_onehotd[1]};
  assign writeNatlizzieLet39_1_argbuf_d = {demuxWriteResult_Nat_d[16:1],
                                           demuxWriteResult_Nat_onehotd[2]};
  assign writeNatlizzieLet40_1_argbuf_d = {demuxWriteResult_Nat_d[16:1],
                                           demuxWriteResult_Nat_onehotd[3]};
  assign demuxWriteResult_Nat_r = (| (demuxWriteResult_Nat_onehotd & {writeNatlizzieLet40_1_argbuf_r,
                                                                      writeNatlizzieLet39_1_argbuf_r,
                                                                      writeNatlizzieLet1_1_argbuf_r,
                                                                      writeNatlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_Nat_r = demuxWriteResult_Nat_r;
  
  /* dcon (Ty MemIn_Nat,Dcon WriteIn_Nat) : [(forkHP1_Na2,Word16#),
                                        (writeMerge_data_Nat,Nat)] > (dconWriteIn_Nat,MemIn_Nat) */
  assign dconWriteIn_Nat_d = WriteIn_Nat_dc((& {forkHP1_Na2_d[0],
                                                writeMerge_data_Nat_d[0]}), forkHP1_Na2_d, writeMerge_data_Nat_d);
  assign {forkHP1_Na2_r,
          writeMerge_data_Nat_r} = {2 {(dconWriteIn_Nat_r && dconWriteIn_Nat_d[0])}};
  
  /* dcon (Ty Pointer_Nat,
      Dcon Pointer_Nat) : [(forkHP1_Na3,Word16#)] > (dconPtr_Nat,Pointer_Nat) */
  assign dconPtr_Nat_d = Pointer_Nat_dc((& {forkHP1_Na3_d[0]}), forkHP1_Na3_d);
  assign {forkHP1_Na3_r} = {1 {(dconPtr_Nat_r && dconPtr_Nat_d[0])}};
  
  /* demux (Ty MemOut_Nat,
       Ty Pointer_Nat) : (memWriteOut_Nat,MemOut_Nat) (dconPtr_Nat,Pointer_Nat) > [(_40,Pointer_Nat),
                                                                                   (demuxWriteResult_Nat,Pointer_Nat)] */
  logic [1:0] dconPtr_Nat_onehotd;
  always_comb
    if ((memWriteOut_Nat_d[0] && dconPtr_Nat_d[0]))
      unique case (memWriteOut_Nat_d[1:1])
        1'd0: dconPtr_Nat_onehotd = 2'd1;
        1'd1: dconPtr_Nat_onehotd = 2'd2;
        default: dconPtr_Nat_onehotd = 2'd0;
      endcase
    else dconPtr_Nat_onehotd = 2'd0;
  assign _40_d = {dconPtr_Nat_d[16:1], dconPtr_Nat_onehotd[0]};
  assign demuxWriteResult_Nat_d = {dconPtr_Nat_d[16:1],
                                   dconPtr_Nat_onehotd[1]};
  assign dconPtr_Nat_r = (| (dconPtr_Nat_onehotd & {demuxWriteResult_Nat_r,
                                                    _40_r}));
  assign memWriteOut_Nat_r = dconPtr_Nat_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTmain_map'_Bool_Nat,Word16#) */
  assign \initHP_CTmain_map'_Bool_Nat_d  = {16'd0, go__9_d[0]};
  assign go__9_r = \initHP_CTmain_map'_Bool_Nat_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmain_map'_Bool_Nat1,Go) > (incrHP_CTmain_map'_Bool_Nat,Word16#) */
  assign \incrHP_CTmain_map'_Bool_Nat_d  = {16'd1,
                                            \incrHP_CTmain_map'_Bool_Nat1_d [0]};
  assign \incrHP_CTmain_map'_Bool_Nat1_r  = \incrHP_CTmain_map'_Bool_Nat_r ;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTmain_map'_Bool_Nat2,Go)] > (incrHP_mergeCTmain_map'_Bool_Nat,Go) */
  logic [1:0] \incrHP_mergeCTmain_map'_Bool_Nat_selected ;
  logic [1:0] \incrHP_mergeCTmain_map'_Bool_Nat_select ;
  always_comb
    begin
      \incrHP_mergeCTmain_map'_Bool_Nat_selected  = 2'd0;
      if ((| \incrHP_mergeCTmain_map'_Bool_Nat_select ))
        \incrHP_mergeCTmain_map'_Bool_Nat_selected  = \incrHP_mergeCTmain_map'_Bool_Nat_select ;
      else
        if (go__10_d[0])
          \incrHP_mergeCTmain_map'_Bool_Nat_selected [0] = 1'd1;
        else if (\incrHP_CTmain_map'_Bool_Nat2_d [0])
          \incrHP_mergeCTmain_map'_Bool_Nat_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Bool_Nat_select  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Bool_Nat_select  <= (\incrHP_mergeCTmain_map'_Bool_Nat_r  ? 2'd0 :
                                                    \incrHP_mergeCTmain_map'_Bool_Nat_selected );
  always_comb
    if (\incrHP_mergeCTmain_map'_Bool_Nat_selected [0])
      \incrHP_mergeCTmain_map'_Bool_Nat_d  = go__10_d;
    else if (\incrHP_mergeCTmain_map'_Bool_Nat_selected [1])
      \incrHP_mergeCTmain_map'_Bool_Nat_d  = \incrHP_CTmain_map'_Bool_Nat2_d ;
    else \incrHP_mergeCTmain_map'_Bool_Nat_d  = 1'd0;
  assign {\incrHP_CTmain_map'_Bool_Nat2_r ,
          go__10_r} = (\incrHP_mergeCTmain_map'_Bool_Nat_r  ? \incrHP_mergeCTmain_map'_Bool_Nat_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmain_map'_Bool_Nat_buf,Go) > [(incrHP_CTmain_map'_Bool_Nat1,Go),
                                                            (incrHP_CTmain_map'_Bool_Nat2,Go)] */
  logic [1:0] \incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmain_map'_Bool_Nat_buf_done ;
  assign \incrHP_CTmain_map'_Bool_Nat1_d  = (\incrHP_mergeCTmain_map'_Bool_Nat_buf_d [0] && (! \incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted [0]));
  assign \incrHP_CTmain_map'_Bool_Nat2_d  = (\incrHP_mergeCTmain_map'_Bool_Nat_buf_d [0] && (! \incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted [1]));
  assign \incrHP_mergeCTmain_map'_Bool_Nat_buf_done  = (\incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted  | ({\incrHP_CTmain_map'_Bool_Nat2_d [0],
                                                                                                           \incrHP_CTmain_map'_Bool_Nat1_d [0]} & {\incrHP_CTmain_map'_Bool_Nat2_r ,
                                                                                                                                                   \incrHP_CTmain_map'_Bool_Nat1_r }));
  assign \incrHP_mergeCTmain_map'_Bool_Nat_buf_r  = (& \incrHP_mergeCTmain_map'_Bool_Nat_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmain_map'_Bool_Nat_buf_emitted  <= (\incrHP_mergeCTmain_map'_Bool_Nat_buf_r  ? 2'd0 :
                                                         \incrHP_mergeCTmain_map'_Bool_Nat_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmain_map'_Bool_Nat,Word16#) (forkHP1_CTmain_map'_Bool_Nat,Word16#) > (addHP_CTmain_map'_Bool_Nat,Word16#) */
  assign \addHP_CTmain_map'_Bool_Nat_d  = {(\incrHP_CTmain_map'_Bool_Nat_d [16:1] + \forkHP1_CTmain_map'_Bool_Nat_d [16:1]),
                                           (\incrHP_CTmain_map'_Bool_Nat_d [0] && \forkHP1_CTmain_map'_Bool_Nat_d [0])};
  assign {\incrHP_CTmain_map'_Bool_Nat_r ,
          \forkHP1_CTmain_map'_Bool_Nat_r } = {2 {(\addHP_CTmain_map'_Bool_Nat_r  && \addHP_CTmain_map'_Bool_Nat_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmain_map'_Bool_Nat,Word16#),
                      (addHP_CTmain_map'_Bool_Nat,Word16#)] > (mergeHP_CTmain_map'_Bool_Nat,Word16#) */
  logic [1:0] \mergeHP_CTmain_map'_Bool_Nat_selected ;
  logic [1:0] \mergeHP_CTmain_map'_Bool_Nat_select ;
  always_comb
    begin
      \mergeHP_CTmain_map'_Bool_Nat_selected  = 2'd0;
      if ((| \mergeHP_CTmain_map'_Bool_Nat_select ))
        \mergeHP_CTmain_map'_Bool_Nat_selected  = \mergeHP_CTmain_map'_Bool_Nat_select ;
      else
        if (\initHP_CTmain_map'_Bool_Nat_d [0])
          \mergeHP_CTmain_map'_Bool_Nat_selected [0] = 1'd1;
        else if (\addHP_CTmain_map'_Bool_Nat_d [0])
          \mergeHP_CTmain_map'_Bool_Nat_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \mergeHP_CTmain_map'_Bool_Nat_select  <= 2'd0;
    else
      \mergeHP_CTmain_map'_Bool_Nat_select  <= (\mergeHP_CTmain_map'_Bool_Nat_r  ? 2'd0 :
                                                \mergeHP_CTmain_map'_Bool_Nat_selected );
  always_comb
    if (\mergeHP_CTmain_map'_Bool_Nat_selected [0])
      \mergeHP_CTmain_map'_Bool_Nat_d  = \initHP_CTmain_map'_Bool_Nat_d ;
    else if (\mergeHP_CTmain_map'_Bool_Nat_selected [1])
      \mergeHP_CTmain_map'_Bool_Nat_d  = \addHP_CTmain_map'_Bool_Nat_d ;
    else \mergeHP_CTmain_map'_Bool_Nat_d  = {16'd0, 1'd0};
  assign {\addHP_CTmain_map'_Bool_Nat_r ,
          \initHP_CTmain_map'_Bool_Nat_r } = (\mergeHP_CTmain_map'_Bool_Nat_r  ? \mergeHP_CTmain_map'_Bool_Nat_selected  :
                                              2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmain_map'_Bool_Nat,Go) > (incrHP_mergeCTmain_map'_Bool_Nat_buf,Go) */
  Go_t \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d ;
  logic \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_r ;
  assign \incrHP_mergeCTmain_map'_Bool_Nat_r  = ((! \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d [0]) || \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmain_map'_Bool_Nat_r )
        \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d  <= \incrHP_mergeCTmain_map'_Bool_Nat_d ;
  Go_t \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf ;
  assign \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_r  = (! \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf [0]);
  assign \incrHP_mergeCTmain_map'_Bool_Nat_buf_d  = (\incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf [0] ? \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf  :
                                                     \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmain_map'_Bool_Nat_buf_r  && \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf [0]))
        \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmain_map'_Bool_Nat_buf_r ) && (! \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf [0])))
        \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_buf  <= \incrHP_mergeCTmain_map'_Bool_Nat_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmain_map'_Bool_Nat,Word16#) > (mergeHP_CTmain_map'_Bool_Nat_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmain_map'_Bool_Nat_bufchan_d ;
  logic \mergeHP_CTmain_map'_Bool_Nat_bufchan_r ;
  assign \mergeHP_CTmain_map'_Bool_Nat_r  = ((! \mergeHP_CTmain_map'_Bool_Nat_bufchan_d [0]) || \mergeHP_CTmain_map'_Bool_Nat_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Bool_Nat_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmain_map'_Bool_Nat_r )
        \mergeHP_CTmain_map'_Bool_Nat_bufchan_d  <= \mergeHP_CTmain_map'_Bool_Nat_d ;
  \Word16#_t  \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf ;
  assign \mergeHP_CTmain_map'_Bool_Nat_bufchan_r  = (! \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf [0]);
  assign \mergeHP_CTmain_map'_Bool_Nat_buf_d  = (\mergeHP_CTmain_map'_Bool_Nat_bufchan_buf [0] ? \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf  :
                                                 \mergeHP_CTmain_map'_Bool_Nat_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTmain_map'_Bool_Nat_buf_r  && \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf [0]))
        \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTmain_map'_Bool_Nat_buf_r ) && (! \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf [0])))
        \mergeHP_CTmain_map'_Bool_Nat_bufchan_buf  <= \mergeHP_CTmain_map'_Bool_Nat_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmain_map'_Bool_Nat_buf,Word16#) > [(forkHP1_CTmain_map'_Bool_Nat,Word16#),
                                                                  (forkHP1_CTmain_map'_Bool_Na2,Word16#),
                                                                  (forkHP1_CTmain_map'_Bool_Na3,Word16#)] */
  logic [2:0] \mergeHP_CTmain_map'_Bool_Nat_buf_emitted ;
  logic [2:0] \mergeHP_CTmain_map'_Bool_Nat_buf_done ;
  assign \forkHP1_CTmain_map'_Bool_Nat_d  = {\mergeHP_CTmain_map'_Bool_Nat_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Bool_Nat_buf_d [0] && (! \mergeHP_CTmain_map'_Bool_Nat_buf_emitted [0]))};
  assign \forkHP1_CTmain_map'_Bool_Na2_d  = {\mergeHP_CTmain_map'_Bool_Nat_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Bool_Nat_buf_d [0] && (! \mergeHP_CTmain_map'_Bool_Nat_buf_emitted [1]))};
  assign \forkHP1_CTmain_map'_Bool_Na3_d  = {\mergeHP_CTmain_map'_Bool_Nat_buf_d [16:1],
                                             (\mergeHP_CTmain_map'_Bool_Nat_buf_d [0] && (! \mergeHP_CTmain_map'_Bool_Nat_buf_emitted [2]))};
  assign \mergeHP_CTmain_map'_Bool_Nat_buf_done  = (\mergeHP_CTmain_map'_Bool_Nat_buf_emitted  | ({\forkHP1_CTmain_map'_Bool_Na3_d [0],
                                                                                                   \forkHP1_CTmain_map'_Bool_Na2_d [0],
                                                                                                   \forkHP1_CTmain_map'_Bool_Nat_d [0]} & {\forkHP1_CTmain_map'_Bool_Na3_r ,
                                                                                                                                           \forkHP1_CTmain_map'_Bool_Na2_r ,
                                                                                                                                           \forkHP1_CTmain_map'_Bool_Nat_r }));
  assign \mergeHP_CTmain_map'_Bool_Nat_buf_r  = (& \mergeHP_CTmain_map'_Bool_Nat_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmain_map'_Bool_Nat_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmain_map'_Bool_Nat_buf_emitted  <= (\mergeHP_CTmain_map'_Bool_Nat_buf_r  ? 3'd0 :
                                                     \mergeHP_CTmain_map'_Bool_Nat_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmain_map'_Bool_Nat) : [(dconReadIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat),
                                             (dconWriteIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat)] > (memMergeChoice_CTmain_map'_Bool_Nat,C2) (memMergeIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat) */
  logic [1:0] \dconReadIn_CTmain_map'_Bool_Nat_select_d ;
  assign \dconReadIn_CTmain_map'_Bool_Nat_select_d  = ((| \dconReadIn_CTmain_map'_Bool_Nat_select_q ) ? \dconReadIn_CTmain_map'_Bool_Nat_select_q  :
                                                       (\dconReadIn_CTmain_map'_Bool_Nat_d [0] ? 2'd1 :
                                                        (\dconWriteIn_CTmain_map'_Bool_Nat_d [0] ? 2'd2 :
                                                         2'd0)));
  logic [1:0] \dconReadIn_CTmain_map'_Bool_Nat_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Bool_Nat_select_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Bool_Nat_select_q  <= (\dconReadIn_CTmain_map'_Bool_Nat_done  ? 2'd0 :
                                                     \dconReadIn_CTmain_map'_Bool_Nat_select_d );
  logic [1:0] \dconReadIn_CTmain_map'_Bool_Nat_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmain_map'_Bool_Nat_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmain_map'_Bool_Nat_emit_q  <= (\dconReadIn_CTmain_map'_Bool_Nat_done  ? 2'd0 :
                                                   \dconReadIn_CTmain_map'_Bool_Nat_emit_d );
  logic [1:0] \dconReadIn_CTmain_map'_Bool_Nat_emit_d ;
  assign \dconReadIn_CTmain_map'_Bool_Nat_emit_d  = (\dconReadIn_CTmain_map'_Bool_Nat_emit_q  | ({\memMergeChoice_CTmain_map'_Bool_Nat_d [0],
                                                                                                  \memMergeIn_CTmain_map'_Bool_Nat_d [0]} & {\memMergeChoice_CTmain_map'_Bool_Nat_r ,
                                                                                                                                             \memMergeIn_CTmain_map'_Bool_Nat_r }));
  logic \dconReadIn_CTmain_map'_Bool_Nat_done ;
  assign \dconReadIn_CTmain_map'_Bool_Nat_done  = (& \dconReadIn_CTmain_map'_Bool_Nat_emit_d );
  assign {\dconWriteIn_CTmain_map'_Bool_Nat_r ,
          \dconReadIn_CTmain_map'_Bool_Nat_r } = (\dconReadIn_CTmain_map'_Bool_Nat_done  ? \dconReadIn_CTmain_map'_Bool_Nat_select_d  :
                                                  2'd0);
  assign \memMergeIn_CTmain_map'_Bool_Nat_d  = ((\dconReadIn_CTmain_map'_Bool_Nat_select_d [0] && (! \dconReadIn_CTmain_map'_Bool_Nat_emit_q [0])) ? \dconReadIn_CTmain_map'_Bool_Nat_d  :
                                                ((\dconReadIn_CTmain_map'_Bool_Nat_select_d [1] && (! \dconReadIn_CTmain_map'_Bool_Nat_emit_q [0])) ? \dconWriteIn_CTmain_map'_Bool_Nat_d  :
                                                 {84'd0, 1'd0}));
  assign \memMergeChoice_CTmain_map'_Bool_Nat_d  = ((\dconReadIn_CTmain_map'_Bool_Nat_select_d [0] && (! \dconReadIn_CTmain_map'_Bool_Nat_emit_q [1])) ? C1_2_dc(1'd1) :
                                                    ((\dconReadIn_CTmain_map'_Bool_Nat_select_d [1] && (! \dconReadIn_CTmain_map'_Bool_Nat_emit_q [1])) ? C2_2_dc(1'd1) :
                                                     {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmain_map'_Bool_Nat,
      Ty MemOut_CTmain_map'_Bool_Nat) : (memMergeIn_CTmain_map'_Bool_Nat_dbuf,MemIn_CTmain_map'_Bool_Nat) > (memOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat) */
  logic [66:0] \memMergeIn_CTmain_map'_Bool_Nat_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmain_map'_Bool_Nat_dbuf_address ;
  logic [66:0] \memMergeIn_CTmain_map'_Bool_Nat_dbuf_din ;
  logic [66:0] \memOut_CTmain_map'_Bool_Nat_q ;
  logic \memOut_CTmain_map'_Bool_Nat_valid ;
  logic \memMergeIn_CTmain_map'_Bool_Nat_dbuf_we ;
  logic \memOut_CTmain_map'_Bool_Nat_we ;
  assign \memMergeIn_CTmain_map'_Bool_Nat_dbuf_din  = \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [84:18];
  assign \memMergeIn_CTmain_map'_Bool_Nat_dbuf_address  = \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [17:2];
  assign \memMergeIn_CTmain_map'_Bool_Nat_dbuf_we  = (\memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [1:1] && \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmain_map'_Bool_Nat_we  <= 1'd0;
        \memOut_CTmain_map'_Bool_Nat_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmain_map'_Bool_Nat_we  <= \memMergeIn_CTmain_map'_Bool_Nat_dbuf_we ;
        \memOut_CTmain_map'_Bool_Nat_valid  <= \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [0];
        if (\memMergeIn_CTmain_map'_Bool_Nat_dbuf_we )
          begin
            \memMergeIn_CTmain_map'_Bool_Nat_dbuf_mem [\memMergeIn_CTmain_map'_Bool_Nat_dbuf_address ] <= \memMergeIn_CTmain_map'_Bool_Nat_dbuf_din ;
            \memOut_CTmain_map'_Bool_Nat_q  <= \memMergeIn_CTmain_map'_Bool_Nat_dbuf_din ;
          end
        else
          \memOut_CTmain_map'_Bool_Nat_q  <= \memMergeIn_CTmain_map'_Bool_Nat_dbuf_mem [\memMergeIn_CTmain_map'_Bool_Nat_dbuf_address ];
      end
  assign \memOut_CTmain_map'_Bool_Nat_d  = {\memOut_CTmain_map'_Bool_Nat_q ,
                                            \memOut_CTmain_map'_Bool_Nat_we ,
                                            \memOut_CTmain_map'_Bool_Nat_valid };
  assign \memMergeIn_CTmain_map'_Bool_Nat_dbuf_r  = ((! \memOut_CTmain_map'_Bool_Nat_valid ) || \memOut_CTmain_map'_Bool_Nat_r );
  logic [31:0] \profiling_MemIn_CTmain_map'_Bool_Nat_read ;
  logic [31:0] \profiling_MemIn_CTmain_map'_Bool_Nat_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTmain_map'_Bool_Nat_write  <= 0;
        \profiling_MemIn_CTmain_map'_Bool_Nat_read  <= 0;
      end
    else
      if ((\memMergeIn_CTmain_map'_Bool_Nat_dbuf_we  == 1'd1))
        \profiling_MemIn_CTmain_map'_Bool_Nat_write  <= (\profiling_MemIn_CTmain_map'_Bool_Nat_write  + 1);
      else
        if ((\memOut_CTmain_map'_Bool_Nat_valid  == 1'd1))
          \profiling_MemIn_CTmain_map'_Bool_Nat_read  <= (\profiling_MemIn_CTmain_map'_Bool_Nat_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmain_map'_Bool_Nat) : (memMergeChoice_CTmain_map'_Bool_Nat,C2) (memOut_CTmain_map'_Bool_Nat_dbuf,MemOut_CTmain_map'_Bool_Nat) > [(memReadOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat),
                                                                                                                                                    (memWriteOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat)] */
  logic [1:0] \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmain_map'_Bool_Nat_d [0] && \memOut_CTmain_map'_Bool_Nat_dbuf_d [0]))
      unique case (\memMergeChoice_CTmain_map'_Bool_Nat_d [1:1])
        1'd0: \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmain_map'_Bool_Nat_d  = {\memOut_CTmain_map'_Bool_Nat_dbuf_d [68:1],
                                                \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd [0]};
  assign \memWriteOut_CTmain_map'_Bool_Nat_d  = {\memOut_CTmain_map'_Bool_Nat_dbuf_d [68:1],
                                                 \memOut_CTmain_map'_Bool_Nat_dbuf_onehotd [1]};
  assign \memOut_CTmain_map'_Bool_Nat_dbuf_r  = (| (\memOut_CTmain_map'_Bool_Nat_dbuf_onehotd  & {\memWriteOut_CTmain_map'_Bool_Nat_r ,
                                                                                                  \memReadOut_CTmain_map'_Bool_Nat_r }));
  assign \memMergeChoice_CTmain_map'_Bool_Nat_r  = \memOut_CTmain_map'_Bool_Nat_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmain_map'_Bool_Nat) : (memMergeIn_CTmain_map'_Bool_Nat_rbuf,MemIn_CTmain_map'_Bool_Nat) > (memMergeIn_CTmain_map'_Bool_Nat_dbuf,MemIn_CTmain_map'_Bool_Nat) */
  assign \memMergeIn_CTmain_map'_Bool_Nat_rbuf_r  = ((! \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d [0]) || \memMergeIn_CTmain_map'_Bool_Nat_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d  <= {84'd0, 1'd0};
    else
      if (\memMergeIn_CTmain_map'_Bool_Nat_rbuf_r )
        \memMergeIn_CTmain_map'_Bool_Nat_dbuf_d  <= \memMergeIn_CTmain_map'_Bool_Nat_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmain_map'_Bool_Nat) : (memMergeIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat) > (memMergeIn_CTmain_map'_Bool_Nat_rbuf,MemIn_CTmain_map'_Bool_Nat) */
  \MemIn_CTmain_map'_Bool_Nat_t  \memMergeIn_CTmain_map'_Bool_Nat_buf ;
  assign \memMergeIn_CTmain_map'_Bool_Nat_r  = (! \memMergeIn_CTmain_map'_Bool_Nat_buf [0]);
  assign \memMergeIn_CTmain_map'_Bool_Nat_rbuf_d  = (\memMergeIn_CTmain_map'_Bool_Nat_buf [0] ? \memMergeIn_CTmain_map'_Bool_Nat_buf  :
                                                     \memMergeIn_CTmain_map'_Bool_Nat_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmain_map'_Bool_Nat_buf  <= {84'd0, 1'd0};
    else
      if ((\memMergeIn_CTmain_map'_Bool_Nat_rbuf_r  && \memMergeIn_CTmain_map'_Bool_Nat_buf [0]))
        \memMergeIn_CTmain_map'_Bool_Nat_buf  <= {84'd0, 1'd0};
      else if (((! \memMergeIn_CTmain_map'_Bool_Nat_rbuf_r ) && (! \memMergeIn_CTmain_map'_Bool_Nat_buf [0])))
        \memMergeIn_CTmain_map'_Bool_Nat_buf  <= \memMergeIn_CTmain_map'_Bool_Nat_d ;
  
  /* dbuf (Ty MemOut_CTmain_map'_Bool_Nat) : (memOut_CTmain_map'_Bool_Nat_rbuf,MemOut_CTmain_map'_Bool_Nat) > (memOut_CTmain_map'_Bool_Nat_dbuf,MemOut_CTmain_map'_Bool_Nat) */
  assign \memOut_CTmain_map'_Bool_Nat_rbuf_r  = ((! \memOut_CTmain_map'_Bool_Nat_dbuf_d [0]) || \memOut_CTmain_map'_Bool_Nat_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Bool_Nat_dbuf_d  <= {68'd0, 1'd0};
    else
      if (\memOut_CTmain_map'_Bool_Nat_rbuf_r )
        \memOut_CTmain_map'_Bool_Nat_dbuf_d  <= \memOut_CTmain_map'_Bool_Nat_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmain_map'_Bool_Nat) : (memOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat) > (memOut_CTmain_map'_Bool_Nat_rbuf,MemOut_CTmain_map'_Bool_Nat) */
  \MemOut_CTmain_map'_Bool_Nat_t  \memOut_CTmain_map'_Bool_Nat_buf ;
  assign \memOut_CTmain_map'_Bool_Nat_r  = (! \memOut_CTmain_map'_Bool_Nat_buf [0]);
  assign \memOut_CTmain_map'_Bool_Nat_rbuf_d  = (\memOut_CTmain_map'_Bool_Nat_buf [0] ? \memOut_CTmain_map'_Bool_Nat_buf  :
                                                 \memOut_CTmain_map'_Bool_Nat_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmain_map'_Bool_Nat_buf  <= {68'd0, 1'd0};
    else
      if ((\memOut_CTmain_map'_Bool_Nat_rbuf_r  && \memOut_CTmain_map'_Bool_Nat_buf [0]))
        \memOut_CTmain_map'_Bool_Nat_buf  <= {68'd0, 1'd0};
      else if (((! \memOut_CTmain_map'_Bool_Nat_rbuf_r ) && (! \memOut_CTmain_map'_Bool_Nat_buf [0])))
        \memOut_CTmain_map'_Bool_Nat_buf  <= \memOut_CTmain_map'_Bool_Nat_d ;
  
  /* destruct (Ty Pointer_CTmain_map'_Bool_Nat,
          Dcon Pointer_CTmain_map'_Bool_Nat) : (scfarg_0_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > [(destructReadIn_CTmain_map'_Bool_Nat,Word16#)] */
  assign \destructReadIn_CTmain_map'_Bool_Nat_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                    scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTmain_map'_Bool_Nat_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Bool_Nat,
      Dcon ReadIn_CTmain_map'_Bool_Nat) : [(destructReadIn_CTmain_map'_Bool_Nat,Word16#)] > (dconReadIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat) */
  assign \dconReadIn_CTmain_map'_Bool_Nat_d  = \ReadIn_CTmain_map'_Bool_Nat_dc ((& {\destructReadIn_CTmain_map'_Bool_Nat_d [0]}), \destructReadIn_CTmain_map'_Bool_Nat_d );
  assign {\destructReadIn_CTmain_map'_Bool_Nat_r } = {1 {(\dconReadIn_CTmain_map'_Bool_Nat_r  && \dconReadIn_CTmain_map'_Bool_Nat_d [0])}};
  
  /* destruct (Ty MemOut_CTmain_map'_Bool_Nat,
          Dcon ReadOut_CTmain_map'_Bool_Nat) : (memReadOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat) > [(readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf,CTmain_map'_Bool_Nat)] */
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_d  = {\memReadOut_CTmain_map'_Bool_Nat_d [68:2],
                                                                    \memReadOut_CTmain_map'_Bool_Nat_d [0]};
  assign \memReadOut_CTmain_map'_Bool_Nat_r  = \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmain_map'_Bool_Nat) : [(lizzieLet10_1_argbuf,CTmain_map'_Bool_Nat),
                                       (lizzieLet22_1_argbuf,CTmain_map'_Bool_Nat),
                                       (lizzieLet30_1_argbuf,CTmain_map'_Bool_Nat),
                                       (lizzieLet31_1_argbuf,CTmain_map'_Bool_Nat),
                                       (lizzieLet32_1_argbuf,CTmain_map'_Bool_Nat)] > (writeMerge_choice_CTmain_map'_Bool_Nat,C5) (writeMerge_data_CTmain_map'_Bool_Nat,CTmain_map'_Bool_Nat) */
  logic [4:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet22_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet30_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet31_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet32_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 5'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({\writeMerge_choice_CTmain_map'_Bool_Nat_d [0],
                                                                        \writeMerge_data_CTmain_map'_Bool_Nat_d [0]} & {\writeMerge_choice_CTmain_map'_Bool_Nat_r ,
                                                                                                                        \writeMerge_data_CTmain_map'_Bool_Nat_r }));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {lizzieLet32_1_argbuf_r,
          lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmain_map'_Bool_Nat_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                                     ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                                      ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                                       ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                        ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                                         {67'd0, 1'd0})))));
  assign \writeMerge_choice_CTmain_map'_Bool_Nat_d  = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                       ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                        ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                         ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                          ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                           {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmain_map'_Bool_Nat) : (writeMerge_choice_CTmain_map'_Bool_Nat,C5) (demuxWriteResult_CTmain_map'_Bool_Nat,Pointer_CTmain_map'_Bool_Nat) > [(writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                                                              (writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                                                              (writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                                                              (writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                                                              (writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf,Pointer_CTmain_map'_Bool_Nat)] */
  logic [4:0] \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmain_map'_Bool_Nat_d [0] && \demuxWriteResult_CTmain_map'_Bool_Nat_d [0]))
      unique case (\writeMerge_choice_CTmain_map'_Bool_Nat_d [3:1])
        3'd0: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd16;
        default: \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  = 5'd0;
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Bool_Nat_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd [0]};
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Bool_Nat_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd [1]};
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Bool_Nat_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd [2]};
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Bool_Nat_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd [3]};
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_d  = {\demuxWriteResult_CTmain_map'_Bool_Nat_d [16:1],
                                                              \demuxWriteResult_CTmain_map'_Bool_Nat_onehotd [4]};
  assign \demuxWriteResult_CTmain_map'_Bool_Nat_r  = (| (\demuxWriteResult_CTmain_map'_Bool_Nat_onehotd  & {\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_r ,
                                                                                                            \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_r }));
  assign \writeMerge_choice_CTmain_map'_Bool_Nat_r  = \demuxWriteResult_CTmain_map'_Bool_Nat_r ;
  
  /* dcon (Ty MemIn_CTmain_map'_Bool_Nat,
      Dcon WriteIn_CTmain_map'_Bool_Nat) : [(forkHP1_CTmain_map'_Bool_Na2,Word16#),
                                            (writeMerge_data_CTmain_map'_Bool_Nat,CTmain_map'_Bool_Nat)] > (dconWriteIn_CTmain_map'_Bool_Nat,MemIn_CTmain_map'_Bool_Nat) */
  assign \dconWriteIn_CTmain_map'_Bool_Nat_d  = \WriteIn_CTmain_map'_Bool_Nat_dc ((& {\forkHP1_CTmain_map'_Bool_Na2_d [0],
                                                                                      \writeMerge_data_CTmain_map'_Bool_Nat_d [0]}), \forkHP1_CTmain_map'_Bool_Na2_d , \writeMerge_data_CTmain_map'_Bool_Nat_d );
  assign {\forkHP1_CTmain_map'_Bool_Na2_r ,
          \writeMerge_data_CTmain_map'_Bool_Nat_r } = {2 {(\dconWriteIn_CTmain_map'_Bool_Nat_r  && \dconWriteIn_CTmain_map'_Bool_Nat_d [0])}};
  
  /* dcon (Ty Pointer_CTmain_map'_Bool_Nat,
      Dcon Pointer_CTmain_map'_Bool_Nat) : [(forkHP1_CTmain_map'_Bool_Na3,Word16#)] > (dconPtr_CTmain_map'_Bool_Nat,Pointer_CTmain_map'_Bool_Nat) */
  assign \dconPtr_CTmain_map'_Bool_Nat_d  = \Pointer_CTmain_map'_Bool_Nat_dc ((& {\forkHP1_CTmain_map'_Bool_Na3_d [0]}), \forkHP1_CTmain_map'_Bool_Na3_d );
  assign {\forkHP1_CTmain_map'_Bool_Na3_r } = {1 {(\dconPtr_CTmain_map'_Bool_Nat_r  && \dconPtr_CTmain_map'_Bool_Nat_d [0])}};
  
  /* demux (Ty MemOut_CTmain_map'_Bool_Nat,
       Ty Pointer_CTmain_map'_Bool_Nat) : (memWriteOut_CTmain_map'_Bool_Nat,MemOut_CTmain_map'_Bool_Nat) (dconPtr_CTmain_map'_Bool_Nat,Pointer_CTmain_map'_Bool_Nat) > [(_39,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                                                                        (demuxWriteResult_CTmain_map'_Bool_Nat,Pointer_CTmain_map'_Bool_Nat)] */
  logic [1:0] \dconPtr_CTmain_map'_Bool_Nat_onehotd ;
  always_comb
    if ((\memWriteOut_CTmain_map'_Bool_Nat_d [0] && \dconPtr_CTmain_map'_Bool_Nat_d [0]))
      unique case (\memWriteOut_CTmain_map'_Bool_Nat_d [1:1])
        1'd0: \dconPtr_CTmain_map'_Bool_Nat_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmain_map'_Bool_Nat_onehotd  = 2'd2;
        default: \dconPtr_CTmain_map'_Bool_Nat_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmain_map'_Bool_Nat_onehotd  = 2'd0;
  assign _39_d = {\dconPtr_CTmain_map'_Bool_Nat_d [16:1],
                  \dconPtr_CTmain_map'_Bool_Nat_onehotd [0]};
  assign \demuxWriteResult_CTmain_map'_Bool_Nat_d  = {\dconPtr_CTmain_map'_Bool_Nat_d [16:1],
                                                      \dconPtr_CTmain_map'_Bool_Nat_onehotd [1]};
  assign \dconPtr_CTmain_map'_Bool_Nat_r  = (| (\dconPtr_CTmain_map'_Bool_Nat_onehotd  & {\demuxWriteResult_CTmain_map'_Bool_Nat_r ,
                                                                                          _39_r}));
  assign \memWriteOut_CTmain_map'_Bool_Nat_r  = \dconPtr_CTmain_map'_Bool_Nat_r ;
  
  /* const (Ty Word16#,Lit 0) : (go__11,Go) > (initHP_QTree_Nat,Word16#) */
  assign initHP_QTree_Nat_d = {16'd0, go__11_d[0]};
  assign go__11_r = initHP_QTree_Nat_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Nat1,Go) > (incrHP_QTree_Nat,Word16#) */
  assign incrHP_QTree_Nat_d = {16'd1, incrHP_QTree_Nat1_d[0]};
  assign incrHP_QTree_Nat1_r = incrHP_QTree_Nat_r;
  
  /* merge (Ty Go) : [(go__12,Go),
                 (incrHP_QTree_Nat2,Go)] > (incrHP_mergeQTree_Nat,Go) */
  logic [1:0] incrHP_mergeQTree_Nat_selected;
  logic [1:0] incrHP_mergeQTree_Nat_select;
  always_comb
    begin
      incrHP_mergeQTree_Nat_selected = 2'd0;
      if ((| incrHP_mergeQTree_Nat_select))
        incrHP_mergeQTree_Nat_selected = incrHP_mergeQTree_Nat_select;
      else
        if (go__12_d[0]) incrHP_mergeQTree_Nat_selected[0] = 1'd1;
        else if (incrHP_QTree_Nat2_d[0])
          incrHP_mergeQTree_Nat_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Nat_select <= 2'd0;
    else
      incrHP_mergeQTree_Nat_select <= (incrHP_mergeQTree_Nat_r ? 2'd0 :
                                       incrHP_mergeQTree_Nat_selected);
  always_comb
    if (incrHP_mergeQTree_Nat_selected[0])
      incrHP_mergeQTree_Nat_d = go__12_d;
    else if (incrHP_mergeQTree_Nat_selected[1])
      incrHP_mergeQTree_Nat_d = incrHP_QTree_Nat2_d;
    else incrHP_mergeQTree_Nat_d = 1'd0;
  assign {incrHP_QTree_Nat2_r,
          go__12_r} = (incrHP_mergeQTree_Nat_r ? incrHP_mergeQTree_Nat_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Nat_buf,Go) > [(incrHP_QTree_Nat1,Go),
                                                 (incrHP_QTree_Nat2,Go)] */
  logic [1:0] incrHP_mergeQTree_Nat_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Nat_buf_done;
  assign incrHP_QTree_Nat1_d = (incrHP_mergeQTree_Nat_buf_d[0] && (! incrHP_mergeQTree_Nat_buf_emitted[0]));
  assign incrHP_QTree_Nat2_d = (incrHP_mergeQTree_Nat_buf_d[0] && (! incrHP_mergeQTree_Nat_buf_emitted[1]));
  assign incrHP_mergeQTree_Nat_buf_done = (incrHP_mergeQTree_Nat_buf_emitted | ({incrHP_QTree_Nat2_d[0],
                                                                                 incrHP_QTree_Nat1_d[0]} & {incrHP_QTree_Nat2_r,
                                                                                                            incrHP_QTree_Nat1_r}));
  assign incrHP_mergeQTree_Nat_buf_r = (& incrHP_mergeQTree_Nat_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Nat_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Nat_buf_emitted <= (incrHP_mergeQTree_Nat_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Nat_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Nat,Word16#) (forkHP1_QTree_Nat,Word16#) > (addHP_QTree_Nat,Word16#) */
  assign addHP_QTree_Nat_d = {(incrHP_QTree_Nat_d[16:1] + forkHP1_QTree_Nat_d[16:1]),
                              (incrHP_QTree_Nat_d[0] && forkHP1_QTree_Nat_d[0])};
  assign {incrHP_QTree_Nat_r,
          forkHP1_QTree_Nat_r} = {2 {(addHP_QTree_Nat_r && addHP_QTree_Nat_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Nat,Word16#),
                      (addHP_QTree_Nat,Word16#)] > (mergeHP_QTree_Nat,Word16#) */
  logic [1:0] mergeHP_QTree_Nat_selected;
  logic [1:0] mergeHP_QTree_Nat_select;
  always_comb
    begin
      mergeHP_QTree_Nat_selected = 2'd0;
      if ((| mergeHP_QTree_Nat_select))
        mergeHP_QTree_Nat_selected = mergeHP_QTree_Nat_select;
      else
        if (initHP_QTree_Nat_d[0]) mergeHP_QTree_Nat_selected[0] = 1'd1;
        else if (addHP_QTree_Nat_d[0])
          mergeHP_QTree_Nat_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Nat_select <= 2'd0;
    else
      mergeHP_QTree_Nat_select <= (mergeHP_QTree_Nat_r ? 2'd0 :
                                   mergeHP_QTree_Nat_selected);
  always_comb
    if (mergeHP_QTree_Nat_selected[0])
      mergeHP_QTree_Nat_d = initHP_QTree_Nat_d;
    else if (mergeHP_QTree_Nat_selected[1])
      mergeHP_QTree_Nat_d = addHP_QTree_Nat_d;
    else mergeHP_QTree_Nat_d = {16'd0, 1'd0};
  assign {addHP_QTree_Nat_r,
          initHP_QTree_Nat_r} = (mergeHP_QTree_Nat_r ? mergeHP_QTree_Nat_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Nat,Go) > (incrHP_mergeQTree_Nat_buf,Go) */
  Go_t incrHP_mergeQTree_Nat_bufchan_d;
  logic incrHP_mergeQTree_Nat_bufchan_r;
  assign incrHP_mergeQTree_Nat_r = ((! incrHP_mergeQTree_Nat_bufchan_d[0]) || incrHP_mergeQTree_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Nat_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Nat_r)
        incrHP_mergeQTree_Nat_bufchan_d <= incrHP_mergeQTree_Nat_d;
  Go_t incrHP_mergeQTree_Nat_bufchan_buf;
  assign incrHP_mergeQTree_Nat_bufchan_r = (! incrHP_mergeQTree_Nat_bufchan_buf[0]);
  assign incrHP_mergeQTree_Nat_buf_d = (incrHP_mergeQTree_Nat_bufchan_buf[0] ? incrHP_mergeQTree_Nat_bufchan_buf :
                                        incrHP_mergeQTree_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Nat_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Nat_buf_r && incrHP_mergeQTree_Nat_bufchan_buf[0]))
        incrHP_mergeQTree_Nat_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Nat_buf_r) && (! incrHP_mergeQTree_Nat_bufchan_buf[0])))
        incrHP_mergeQTree_Nat_bufchan_buf <= incrHP_mergeQTree_Nat_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Nat,Word16#) > (mergeHP_QTree_Nat_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Nat_bufchan_d;
  logic mergeHP_QTree_Nat_bufchan_r;
  assign mergeHP_QTree_Nat_r = ((! mergeHP_QTree_Nat_bufchan_d[0]) || mergeHP_QTree_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Nat_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Nat_r)
        mergeHP_QTree_Nat_bufchan_d <= mergeHP_QTree_Nat_d;
  \Word16#_t  mergeHP_QTree_Nat_bufchan_buf;
  assign mergeHP_QTree_Nat_bufchan_r = (! mergeHP_QTree_Nat_bufchan_buf[0]);
  assign mergeHP_QTree_Nat_buf_d = (mergeHP_QTree_Nat_bufchan_buf[0] ? mergeHP_QTree_Nat_bufchan_buf :
                                    mergeHP_QTree_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Nat_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Nat_buf_r && mergeHP_QTree_Nat_bufchan_buf[0]))
        mergeHP_QTree_Nat_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Nat_buf_r) && (! mergeHP_QTree_Nat_bufchan_buf[0])))
        mergeHP_QTree_Nat_bufchan_buf <= mergeHP_QTree_Nat_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Nat_buf,Word16#) > [(forkHP1_QTree_Nat,Word16#),
                                                       (forkHP1_QTree_Na2,Word16#),
                                                       (forkHP1_QTree_Na3,Word16#)] */
  logic [2:0] mergeHP_QTree_Nat_buf_emitted;
  logic [2:0] mergeHP_QTree_Nat_buf_done;
  assign forkHP1_QTree_Nat_d = {mergeHP_QTree_Nat_buf_d[16:1],
                                (mergeHP_QTree_Nat_buf_d[0] && (! mergeHP_QTree_Nat_buf_emitted[0]))};
  assign forkHP1_QTree_Na2_d = {mergeHP_QTree_Nat_buf_d[16:1],
                                (mergeHP_QTree_Nat_buf_d[0] && (! mergeHP_QTree_Nat_buf_emitted[1]))};
  assign forkHP1_QTree_Na3_d = {mergeHP_QTree_Nat_buf_d[16:1],
                                (mergeHP_QTree_Nat_buf_d[0] && (! mergeHP_QTree_Nat_buf_emitted[2]))};
  assign mergeHP_QTree_Nat_buf_done = (mergeHP_QTree_Nat_buf_emitted | ({forkHP1_QTree_Na3_d[0],
                                                                         forkHP1_QTree_Na2_d[0],
                                                                         forkHP1_QTree_Nat_d[0]} & {forkHP1_QTree_Na3_r,
                                                                                                    forkHP1_QTree_Na2_r,
                                                                                                    forkHP1_QTree_Nat_r}));
  assign mergeHP_QTree_Nat_buf_r = (& mergeHP_QTree_Nat_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Nat_buf_emitted <= 3'd0;
    else
      mergeHP_QTree_Nat_buf_emitted <= (mergeHP_QTree_Nat_buf_r ? 3'd0 :
                                        mergeHP_QTree_Nat_buf_done);
  
  /* bram (Ty MemIn_QTree_Nat,
      Ty MemOut_QTree_Nat) : (dconWriteIn_QTree_Nat,MemIn_QTree_Nat) > (memWriteOut_QTree_Nat,MemOut_QTree_Nat) */
  logic [65:0] dconWriteIn_QTree_Nat_mem[65535:0];
  logic [15:0] dconWriteIn_QTree_Nat_address;
  logic [65:0] dconWriteIn_QTree_Nat_din;
  logic [65:0] memWriteOut_QTree_Nat_q;
  logic memWriteOut_QTree_Nat_valid;
  logic dconWriteIn_QTree_Nat_we;
  logic memWriteOut_QTree_Nat_we;
  assign dconWriteIn_QTree_Nat_din = dconWriteIn_QTree_Nat_d[83:18];
  assign dconWriteIn_QTree_Nat_address = dconWriteIn_QTree_Nat_d[17:2];
  assign dconWriteIn_QTree_Nat_we = (dconWriteIn_QTree_Nat_d[1:1] && dconWriteIn_QTree_Nat_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memWriteOut_QTree_Nat_we <= 1'd0;
        memWriteOut_QTree_Nat_valid <= 1'd0;
      end
    else
      begin
        memWriteOut_QTree_Nat_we <= dconWriteIn_QTree_Nat_we;
        memWriteOut_QTree_Nat_valid <= dconWriteIn_QTree_Nat_d[0];
        if (dconWriteIn_QTree_Nat_we)
          begin
            dconWriteIn_QTree_Nat_mem[dconWriteIn_QTree_Nat_address] <= dconWriteIn_QTree_Nat_din;
            memWriteOut_QTree_Nat_q <= dconWriteIn_QTree_Nat_din;
          end
        else
          memWriteOut_QTree_Nat_q <= dconWriteIn_QTree_Nat_mem[dconWriteIn_QTree_Nat_address];
      end
  assign memWriteOut_QTree_Nat_d = {memWriteOut_QTree_Nat_q,
                                    memWriteOut_QTree_Nat_we,
                                    memWriteOut_QTree_Nat_valid};
  assign dconWriteIn_QTree_Nat_r = ((! memWriteOut_QTree_Nat_valid) || memWriteOut_QTree_Nat_r);
  logic [31:0] profiling_MemIn_QTree_Nat_read;
  logic [31:0] profiling_MemIn_QTree_Nat_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Nat_write <= 0;
        profiling_MemIn_QTree_Nat_read <= 0;
      end
    else
      if ((dconWriteIn_QTree_Nat_we == 1'd1))
        profiling_MemIn_QTree_Nat_write <= (profiling_MemIn_QTree_Nat_write + 1);
      else
        if ((memWriteOut_QTree_Nat_valid == 1'd1))
          profiling_MemIn_QTree_Nat_read <= (profiling_MemIn_QTree_Nat_read + 1);
  
  /* mergectrl (Ty C5,
           Ty QTree_Nat) : [(lizzieLet11_1_1_argbuf,QTree_Nat),
                            (lizzieLet33_1_argbuf,QTree_Nat),
                            (lizzieLet7_1_argbuf,QTree_Nat),
                            (lizzieLet8_1_argbuf,QTree_Nat),
                            (lizzieLet9_1_argbuf,QTree_Nat)] > (writeMerge_choice_QTree_Nat,C5) (writeMerge_data_QTree_Nat,QTree_Nat) */
  logic [4:0] lizzieLet11_1_1_argbuf_select_d;
  assign lizzieLet11_1_1_argbuf_select_d = ((| lizzieLet11_1_1_argbuf_select_q) ? lizzieLet11_1_1_argbuf_select_q :
                                            (lizzieLet11_1_1_argbuf_d[0] ? 5'd1 :
                                             (lizzieLet33_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet7_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet8_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet9_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] lizzieLet11_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet11_1_1_argbuf_select_q <= (lizzieLet11_1_1_argbuf_done ? 5'd0 :
                                          lizzieLet11_1_1_argbuf_select_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_1_1_argbuf_emit_q <= (lizzieLet11_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet11_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_1_1_argbuf_emit_d;
  assign lizzieLet11_1_1_argbuf_emit_d = (lizzieLet11_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Nat_d[0],
                                                                            writeMerge_data_QTree_Nat_d[0]} & {writeMerge_choice_QTree_Nat_r,
                                                                                                               writeMerge_data_QTree_Nat_r}));
  logic lizzieLet11_1_1_argbuf_done;
  assign lizzieLet11_1_1_argbuf_done = (& lizzieLet11_1_1_argbuf_emit_d);
  assign {lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet33_1_argbuf_r,
          lizzieLet11_1_1_argbuf_r} = (lizzieLet11_1_1_argbuf_done ? lizzieLet11_1_1_argbuf_select_d :
                                       5'd0);
  assign writeMerge_data_QTree_Nat_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet11_1_1_argbuf_d :
                                        ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet33_1_argbuf_d :
                                         ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                          ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                           ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                            {66'd0, 1'd0})))));
  assign writeMerge_choice_QTree_Nat_d = ((lizzieLet11_1_1_argbuf_select_d[0] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                          ((lizzieLet11_1_1_argbuf_select_d[1] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                           ((lizzieLet11_1_1_argbuf_select_d[2] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                            ((lizzieLet11_1_1_argbuf_select_d[3] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                             ((lizzieLet11_1_1_argbuf_select_d[4] && (! lizzieLet11_1_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_QTree_Nat) : (writeMerge_choice_QTree_Nat,C5) (demuxWriteResult_QTree_Nat,Pointer_QTree_Nat) > [(writeQTree_NatlizzieLet11_1_1_argbuf,Pointer_QTree_Nat),
                                                                                                                  (writeQTree_NatlizzieLet33_1_argbuf,Pointer_QTree_Nat),
                                                                                                                  (writeQTree_NatlizzieLet7_1_argbuf,Pointer_QTree_Nat),
                                                                                                                  (writeQTree_NatlizzieLet8_1_argbuf,Pointer_QTree_Nat),
                                                                                                                  (writeQTree_NatlizzieLet9_1_argbuf,Pointer_QTree_Nat)] */
  logic [4:0] demuxWriteResult_QTree_Nat_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Nat_d[0] && demuxWriteResult_QTree_Nat_d[0]))
      unique case (writeMerge_choice_QTree_Nat_d[3:1])
        3'd0: demuxWriteResult_QTree_Nat_onehotd = 5'd1;
        3'd1: demuxWriteResult_QTree_Nat_onehotd = 5'd2;
        3'd2: demuxWriteResult_QTree_Nat_onehotd = 5'd4;
        3'd3: demuxWriteResult_QTree_Nat_onehotd = 5'd8;
        3'd4: demuxWriteResult_QTree_Nat_onehotd = 5'd16;
        default: demuxWriteResult_QTree_Nat_onehotd = 5'd0;
      endcase
    else demuxWriteResult_QTree_Nat_onehotd = 5'd0;
  assign writeQTree_NatlizzieLet11_1_1_argbuf_d = {demuxWriteResult_QTree_Nat_d[16:1],
                                                   demuxWriteResult_QTree_Nat_onehotd[0]};
  assign writeQTree_NatlizzieLet33_1_argbuf_d = {demuxWriteResult_QTree_Nat_d[16:1],
                                                 demuxWriteResult_QTree_Nat_onehotd[1]};
  assign writeQTree_NatlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Nat_d[16:1],
                                                demuxWriteResult_QTree_Nat_onehotd[2]};
  assign writeQTree_NatlizzieLet8_1_argbuf_d = {demuxWriteResult_QTree_Nat_d[16:1],
                                                demuxWriteResult_QTree_Nat_onehotd[3]};
  assign writeQTree_NatlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Nat_d[16:1],
                                                demuxWriteResult_QTree_Nat_onehotd[4]};
  assign demuxWriteResult_QTree_Nat_r = (| (demuxWriteResult_QTree_Nat_onehotd & {writeQTree_NatlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_NatlizzieLet8_1_argbuf_r,
                                                                                  writeQTree_NatlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_NatlizzieLet33_1_argbuf_r,
                                                                                  writeQTree_NatlizzieLet11_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Nat_r = demuxWriteResult_QTree_Nat_r;
  
  /* dcon (Ty MemIn_QTree_Nat,
      Dcon WriteIn_QTree_Nat) : [(forkHP1_QTree_Na2,Word16#),
                                 (writeMerge_data_QTree_Nat,QTree_Nat)] > (dconWriteIn_QTree_Nat,MemIn_QTree_Nat) */
  assign dconWriteIn_QTree_Nat_d = WriteIn_QTree_Nat_dc((& {forkHP1_QTree_Na2_d[0],
                                                            writeMerge_data_QTree_Nat_d[0]}), forkHP1_QTree_Na2_d, writeMerge_data_QTree_Nat_d);
  assign {forkHP1_QTree_Na2_r,
          writeMerge_data_QTree_Nat_r} = {2 {(dconWriteIn_QTree_Nat_r && dconWriteIn_QTree_Nat_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Nat,
      Dcon Pointer_QTree_Nat) : [(forkHP1_QTree_Na3,Word16#)] > (dconPtr_QTree_Nat,Pointer_QTree_Nat) */
  assign dconPtr_QTree_Nat_d = Pointer_QTree_Nat_dc((& {forkHP1_QTree_Na3_d[0]}), forkHP1_QTree_Na3_d);
  assign {forkHP1_QTree_Na3_r} = {1 {(dconPtr_QTree_Nat_r && dconPtr_QTree_Nat_d[0])}};
  
  /* demux (Ty MemOut_QTree_Nat,
       Ty Pointer_QTree_Nat) : (memWriteOut_QTree_Nat,MemOut_QTree_Nat) (dconPtr_QTree_Nat,Pointer_QTree_Nat) > [(_38,Pointer_QTree_Nat),
                                                                                                                 (demuxWriteResult_QTree_Nat,Pointer_QTree_Nat)] */
  logic [1:0] dconPtr_QTree_Nat_onehotd;
  always_comb
    if ((memWriteOut_QTree_Nat_d[0] && dconPtr_QTree_Nat_d[0]))
      unique case (memWriteOut_QTree_Nat_d[1:1])
        1'd0: dconPtr_QTree_Nat_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Nat_onehotd = 2'd2;
        default: dconPtr_QTree_Nat_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Nat_onehotd = 2'd0;
  assign _38_d = {dconPtr_QTree_Nat_d[16:1],
                  dconPtr_QTree_Nat_onehotd[0]};
  assign demuxWriteResult_QTree_Nat_d = {dconPtr_QTree_Nat_d[16:1],
                                         dconPtr_QTree_Nat_onehotd[1]};
  assign dconPtr_QTree_Nat_r = (| (dconPtr_QTree_Nat_onehotd & {demuxWriteResult_QTree_Nat_r,
                                                                _38_r}));
  assign memWriteOut_QTree_Nat_r = dconPtr_QTree_Nat_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Bool,Go) > (initHP_QTree_Bool,Word16#) */
  assign initHP_QTree_Bool_d = {16'd0,
                                go_1_dummy_write_QTree_Bool_d[0]};
  assign go_1_dummy_write_QTree_Bool_r = initHP_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Bool1,Go) > (incrHP_QTree_Bool,Word16#) */
  assign incrHP_QTree_Bool_d = {16'd1, incrHP_QTree_Bool1_d[0]};
  assign incrHP_QTree_Bool1_r = incrHP_QTree_Bool_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Bool,Go),
                 (incrHP_QTree_Bool2,Go)] > (incrHP_mergeQTree_Bool,Go) */
  logic [1:0] incrHP_mergeQTree_Bool_selected;
  logic [1:0] incrHP_mergeQTree_Bool_select;
  always_comb
    begin
      incrHP_mergeQTree_Bool_selected = 2'd0;
      if ((| incrHP_mergeQTree_Bool_select))
        incrHP_mergeQTree_Bool_selected = incrHP_mergeQTree_Bool_select;
      else
        if (go_2_dummy_write_QTree_Bool_d[0])
          incrHP_mergeQTree_Bool_selected[0] = 1'd1;
        else if (incrHP_QTree_Bool2_d[0])
          incrHP_mergeQTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_select <= 2'd0;
    else
      incrHP_mergeQTree_Bool_select <= (incrHP_mergeQTree_Bool_r ? 2'd0 :
                                        incrHP_mergeQTree_Bool_selected);
  always_comb
    if (incrHP_mergeQTree_Bool_selected[0])
      incrHP_mergeQTree_Bool_d = go_2_dummy_write_QTree_Bool_d;
    else if (incrHP_mergeQTree_Bool_selected[1])
      incrHP_mergeQTree_Bool_d = incrHP_QTree_Bool2_d;
    else incrHP_mergeQTree_Bool_d = 1'd0;
  assign {incrHP_QTree_Bool2_r,
          go_2_dummy_write_QTree_Bool_r} = (incrHP_mergeQTree_Bool_r ? incrHP_mergeQTree_Bool_selected :
                                            2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Bool_buf,Go) > [(incrHP_QTree_Bool1,Go),
                                                  (incrHP_QTree_Bool2,Go)] */
  logic [1:0] incrHP_mergeQTree_Bool_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Bool_buf_done;
  assign incrHP_QTree_Bool1_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[0]));
  assign incrHP_QTree_Bool2_d = (incrHP_mergeQTree_Bool_buf_d[0] && (! incrHP_mergeQTree_Bool_buf_emitted[1]));
  assign incrHP_mergeQTree_Bool_buf_done = (incrHP_mergeQTree_Bool_buf_emitted | ({incrHP_QTree_Bool2_d[0],
                                                                                   incrHP_QTree_Bool1_d[0]} & {incrHP_QTree_Bool2_r,
                                                                                                               incrHP_QTree_Bool1_r}));
  assign incrHP_mergeQTree_Bool_buf_r = (& incrHP_mergeQTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Bool_buf_emitted <= (incrHP_mergeQTree_Bool_buf_r ? 2'd0 :
                                             incrHP_mergeQTree_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Bool,Word16#) (forkHP1_QTree_Bool,Word16#) > (addHP_QTree_Bool,Word16#) */
  assign addHP_QTree_Bool_d = {(incrHP_QTree_Bool_d[16:1] + forkHP1_QTree_Bool_d[16:1]),
                               (incrHP_QTree_Bool_d[0] && forkHP1_QTree_Bool_d[0])};
  assign {incrHP_QTree_Bool_r,
          forkHP1_QTree_Bool_r} = {2 {(addHP_QTree_Bool_r && addHP_QTree_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Bool,Word16#),
                      (addHP_QTree_Bool,Word16#)] > (mergeHP_QTree_Bool,Word16#) */
  logic [1:0] mergeHP_QTree_Bool_selected;
  logic [1:0] mergeHP_QTree_Bool_select;
  always_comb
    begin
      mergeHP_QTree_Bool_selected = 2'd0;
      if ((| mergeHP_QTree_Bool_select))
        mergeHP_QTree_Bool_selected = mergeHP_QTree_Bool_select;
      else
        if (initHP_QTree_Bool_d[0]) mergeHP_QTree_Bool_selected[0] = 1'd1;
        else if (addHP_QTree_Bool_d[0])
          mergeHP_QTree_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_select <= 2'd0;
    else
      mergeHP_QTree_Bool_select <= (mergeHP_QTree_Bool_r ? 2'd0 :
                                    mergeHP_QTree_Bool_selected);
  always_comb
    if (mergeHP_QTree_Bool_selected[0])
      mergeHP_QTree_Bool_d = initHP_QTree_Bool_d;
    else if (mergeHP_QTree_Bool_selected[1])
      mergeHP_QTree_Bool_d = addHP_QTree_Bool_d;
    else mergeHP_QTree_Bool_d = {16'd0, 1'd0};
  assign {addHP_QTree_Bool_r,
          initHP_QTree_Bool_r} = (mergeHP_QTree_Bool_r ? mergeHP_QTree_Bool_selected :
                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Bool,Go) > (incrHP_mergeQTree_Bool_buf,Go) */
  Go_t incrHP_mergeQTree_Bool_bufchan_d;
  logic incrHP_mergeQTree_Bool_bufchan_r;
  assign incrHP_mergeQTree_Bool_r = ((! incrHP_mergeQTree_Bool_bufchan_d[0]) || incrHP_mergeQTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Bool_r)
        incrHP_mergeQTree_Bool_bufchan_d <= incrHP_mergeQTree_Bool_d;
  Go_t incrHP_mergeQTree_Bool_bufchan_buf;
  assign incrHP_mergeQTree_Bool_bufchan_r = (! incrHP_mergeQTree_Bool_bufchan_buf[0]);
  assign incrHP_mergeQTree_Bool_buf_d = (incrHP_mergeQTree_Bool_bufchan_buf[0] ? incrHP_mergeQTree_Bool_bufchan_buf :
                                         incrHP_mergeQTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Bool_buf_r && incrHP_mergeQTree_Bool_bufchan_buf[0]))
        incrHP_mergeQTree_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Bool_buf_r) && (! incrHP_mergeQTree_Bool_bufchan_buf[0])))
        incrHP_mergeQTree_Bool_bufchan_buf <= incrHP_mergeQTree_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Bool,Word16#) > (mergeHP_QTree_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Bool_bufchan_d;
  logic mergeHP_QTree_Bool_bufchan_r;
  assign mergeHP_QTree_Bool_r = ((! mergeHP_QTree_Bool_bufchan_d[0]) || mergeHP_QTree_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Bool_r)
        mergeHP_QTree_Bool_bufchan_d <= mergeHP_QTree_Bool_d;
  \Word16#_t  mergeHP_QTree_Bool_bufchan_buf;
  assign mergeHP_QTree_Bool_bufchan_r = (! mergeHP_QTree_Bool_bufchan_buf[0]);
  assign mergeHP_QTree_Bool_buf_d = (mergeHP_QTree_Bool_bufchan_buf[0] ? mergeHP_QTree_Bool_bufchan_buf :
                                     mergeHP_QTree_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Bool_buf_r && mergeHP_QTree_Bool_bufchan_buf[0]))
        mergeHP_QTree_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Bool_buf_r) && (! mergeHP_QTree_Bool_bufchan_buf[0])))
        mergeHP_QTree_Bool_bufchan_buf <= mergeHP_QTree_Bool_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Bool_snk,Word16#) > */
  assign {forkHP1_QTree_Bool_snk_r,
          forkHP1_QTree_Bool_snk_dout} = {forkHP1_QTree_Bool_snk_rout,
                                          forkHP1_QTree_Bool_snk_d};
  
  /* source (Ty Go) : > (\QTree_Bool_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Bool_src,Go) > [(go_1_dummy_write_QTree_Bool,Go),
                                       (go_2_dummy_write_QTree_Bool,Go)] */
  logic [1:0] \\QTree_Bool_src_emitted ;
  logic [1:0] \\QTree_Bool_src_done ;
  assign go_1_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [0]));
  assign go_2_dummy_write_QTree_Bool_d = (\\QTree_Bool_src_d [0] && (! \\QTree_Bool_src_emitted [1]));
  assign \\QTree_Bool_src_done  = (\\QTree_Bool_src_emitted  | ({go_2_dummy_write_QTree_Bool_d[0],
                                                                 go_1_dummy_write_QTree_Bool_d[0]} & {go_2_dummy_write_QTree_Bool_r,
                                                                                                      go_1_dummy_write_QTree_Bool_r}));
  assign \\QTree_Bool_src_r  = (& \\QTree_Bool_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Bool_src_emitted  <= 2'd0;
    else
      \\QTree_Bool_src_emitted  <= (\\QTree_Bool_src_r  ? 2'd0 :
                                    \\QTree_Bool_src_done );
  
  /* source (Ty QTree_Bool) : > (dummy_write_QTree_Bool,QTree_Bool) */
  
  /* sink (Ty Pointer_QTree_Bool) : (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool) > */
  assign {dummy_write_QTree_Bool_sink_r,
          dummy_write_QTree_Bool_sink_dout} = {dummy_write_QTree_Bool_sink_rout,
                                               dummy_write_QTree_Bool_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Bool_buf,Word16#) > [(forkHP1_QTree_Bool,Word16#),
                                                        (forkHP1_QTree_Bool_snk,Word16#),
                                                        (forkHP1_QTree_Boo3,Word16#),
                                                        (forkHP1_QTree_Boo4,Word16#)] */
  logic [3:0] mergeHP_QTree_Bool_buf_emitted;
  logic [3:0] mergeHP_QTree_Bool_buf_done;
  assign forkHP1_QTree_Bool_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[0]))};
  assign forkHP1_QTree_Bool_snk_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                     (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[1]))};
  assign forkHP1_QTree_Boo3_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[2]))};
  assign forkHP1_QTree_Boo4_d = {mergeHP_QTree_Bool_buf_d[16:1],
                                 (mergeHP_QTree_Bool_buf_d[0] && (! mergeHP_QTree_Bool_buf_emitted[3]))};
  assign mergeHP_QTree_Bool_buf_done = (mergeHP_QTree_Bool_buf_emitted | ({forkHP1_QTree_Boo4_d[0],
                                                                           forkHP1_QTree_Boo3_d[0],
                                                                           forkHP1_QTree_Bool_snk_d[0],
                                                                           forkHP1_QTree_Bool_d[0]} & {forkHP1_QTree_Boo4_r,
                                                                                                       forkHP1_QTree_Boo3_r,
                                                                                                       forkHP1_QTree_Bool_snk_r,
                                                                                                       forkHP1_QTree_Bool_r}));
  assign mergeHP_QTree_Bool_buf_r = (& mergeHP_QTree_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Bool_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Bool_buf_emitted <= (mergeHP_QTree_Bool_buf_r ? 4'd0 :
                                         mergeHP_QTree_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Bool) : [(dconReadIn_QTree_Bool,MemIn_QTree_Bool),
                                   (dconWriteIn_QTree_Bool,MemIn_QTree_Bool)] > (memMergeChoice_QTree_Bool,C2) (memMergeIn_QTree_Bool,MemIn_QTree_Bool) */
  logic [1:0] dconReadIn_QTree_Bool_select_d;
  assign dconReadIn_QTree_Bool_select_d = ((| dconReadIn_QTree_Bool_select_q) ? dconReadIn_QTree_Bool_select_q :
                                           (dconReadIn_QTree_Bool_d[0] ? 2'd1 :
                                            (dconWriteIn_QTree_Bool_d[0] ? 2'd2 :
                                             2'd0)));
  logic [1:0] dconReadIn_QTree_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_select_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_select_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                         dconReadIn_QTree_Bool_select_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Bool_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Bool_emit_q <= (dconReadIn_QTree_Bool_done ? 2'd0 :
                                       dconReadIn_QTree_Bool_emit_d);
  logic [1:0] dconReadIn_QTree_Bool_emit_d;
  assign dconReadIn_QTree_Bool_emit_d = (dconReadIn_QTree_Bool_emit_q | ({memMergeChoice_QTree_Bool_d[0],
                                                                          memMergeIn_QTree_Bool_d[0]} & {memMergeChoice_QTree_Bool_r,
                                                                                                         memMergeIn_QTree_Bool_r}));
  logic dconReadIn_QTree_Bool_done;
  assign dconReadIn_QTree_Bool_done = (& dconReadIn_QTree_Bool_emit_d);
  assign {dconWriteIn_QTree_Bool_r,
          dconReadIn_QTree_Bool_r} = (dconReadIn_QTree_Bool_done ? dconReadIn_QTree_Bool_select_d :
                                      2'd0);
  assign memMergeIn_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconReadIn_QTree_Bool_d :
                                    ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[0])) ? dconWriteIn_QTree_Bool_d :
                                     {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Bool_d = ((dconReadIn_QTree_Bool_select_d[0] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                        ((dconReadIn_QTree_Bool_select_d[1] && (! dconReadIn_QTree_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Bool,
      Ty MemOut_QTree_Bool) : (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) > (memOut_QTree_Bool,MemOut_QTree_Bool) */
  logic [65:0] memMergeIn_QTree_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Bool_dbuf_address;
  logic [65:0] memMergeIn_QTree_Bool_dbuf_din;
  logic [65:0] memOut_QTree_Bool_q;
  logic memOut_QTree_Bool_valid;
  logic memMergeIn_QTree_Bool_dbuf_we;
  logic memOut_QTree_Bool_we;
  assign memMergeIn_QTree_Bool_dbuf_din = memMergeIn_QTree_Bool_dbuf_d[83:18];
  assign memMergeIn_QTree_Bool_dbuf_address = memMergeIn_QTree_Bool_dbuf_d[17:2];
  assign memMergeIn_QTree_Bool_dbuf_we = (memMergeIn_QTree_Bool_dbuf_d[1:1] && memMergeIn_QTree_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Bool_we <= 1'd0;
        memOut_QTree_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Bool_we <= memMergeIn_QTree_Bool_dbuf_we;
        memOut_QTree_Bool_valid <= memMergeIn_QTree_Bool_dbuf_d[0];
        if (memMergeIn_QTree_Bool_dbuf_we)
          begin
            memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address] <= memMergeIn_QTree_Bool_dbuf_din;
            memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_din;
          end
        else
          memOut_QTree_Bool_q <= memMergeIn_QTree_Bool_dbuf_mem[memMergeIn_QTree_Bool_dbuf_address];
      end
  assign memOut_QTree_Bool_d = {memOut_QTree_Bool_q,
                                memOut_QTree_Bool_we,
                                memOut_QTree_Bool_valid};
  assign memMergeIn_QTree_Bool_dbuf_r = ((! memOut_QTree_Bool_valid) || memOut_QTree_Bool_r);
  logic [31:0] profiling_MemIn_QTree_Bool_read;
  logic [31:0] profiling_MemIn_QTree_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Bool_write <= 0;
        profiling_MemIn_QTree_Bool_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Bool_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Bool_write <= (profiling_MemIn_QTree_Bool_write + 1);
      else
        if ((memOut_QTree_Bool_valid == 1'd1))
          profiling_MemIn_QTree_Bool_read <= (profiling_MemIn_QTree_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Bool) : (memMergeChoice_QTree_Bool,C2) (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) > [(memReadOut_QTree_Bool,MemOut_QTree_Bool),
                                                                                                            (memWriteOut_QTree_Bool,MemOut_QTree_Bool)] */
  logic [1:0] memOut_QTree_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Bool_d[0] && memOut_QTree_Bool_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Bool_d[1:1])
        1'd0: memOut_QTree_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Bool_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                    memOut_QTree_Bool_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Bool_d = {memOut_QTree_Bool_dbuf_d[67:1],
                                     memOut_QTree_Bool_dbuf_onehotd[1]};
  assign memOut_QTree_Bool_dbuf_r = (| (memOut_QTree_Bool_dbuf_onehotd & {memWriteOut_QTree_Bool_r,
                                                                          memReadOut_QTree_Bool_r}));
  assign memMergeChoice_QTree_Bool_r = memOut_QTree_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_dbuf,MemIn_QTree_Bool) */
  assign memMergeIn_QTree_Bool_rbuf_r = ((! memMergeIn_QTree_Bool_dbuf_d[0]) || memMergeIn_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Bool_rbuf_r)
        memMergeIn_QTree_Bool_dbuf_d <= memMergeIn_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Bool) : (memMergeIn_QTree_Bool,MemIn_QTree_Bool) > (memMergeIn_QTree_Bool_rbuf,MemIn_QTree_Bool) */
  MemIn_QTree_Bool_t memMergeIn_QTree_Bool_buf;
  assign memMergeIn_QTree_Bool_r = (! memMergeIn_QTree_Bool_buf[0]);
  assign memMergeIn_QTree_Bool_rbuf_d = (memMergeIn_QTree_Bool_buf[0] ? memMergeIn_QTree_Bool_buf :
                                         memMergeIn_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Bool_rbuf_r && memMergeIn_QTree_Bool_buf[0]))
        memMergeIn_QTree_Bool_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Bool_rbuf_r) && (! memMergeIn_QTree_Bool_buf[0])))
        memMergeIn_QTree_Bool_buf <= memMergeIn_QTree_Bool_d;
  
  /* dbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) > (memOut_QTree_Bool_dbuf,MemOut_QTree_Bool) */
  assign memOut_QTree_Bool_rbuf_r = ((! memOut_QTree_Bool_dbuf_d[0]) || memOut_QTree_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Bool_rbuf_r)
        memOut_QTree_Bool_dbuf_d <= memOut_QTree_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Bool) : (memOut_QTree_Bool,MemOut_QTree_Bool) > (memOut_QTree_Bool_rbuf,MemOut_QTree_Bool) */
  MemOut_QTree_Bool_t memOut_QTree_Bool_buf;
  assign memOut_QTree_Bool_r = (! memOut_QTree_Bool_buf[0]);
  assign memOut_QTree_Bool_rbuf_d = (memOut_QTree_Bool_buf[0] ? memOut_QTree_Bool_buf :
                                     memOut_QTree_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Bool_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Bool_rbuf_r && memOut_QTree_Bool_buf[0]))
        memOut_QTree_Bool_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Bool_rbuf_r) && (! memOut_QTree_Bool_buf[0])))
        memOut_QTree_Bool_buf <= memOut_QTree_Bool_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Bool) : [(m1ad9_1_argbuf,Pointer_QTree_Bool),
                                     (macS_1_argbuf,Pointer_QTree_Bool),
                                     (mad1_1_argbuf,Pointer_QTree_Bool)] > (readMerge_choice_QTree_Bool,C3) (readMerge_data_QTree_Bool,Pointer_QTree_Bool) */
  logic [2:0] m1ad9_1_argbuf_select_d;
  assign m1ad9_1_argbuf_select_d = ((| m1ad9_1_argbuf_select_q) ? m1ad9_1_argbuf_select_q :
                                    (m1ad9_1_argbuf_d[0] ? 3'd1 :
                                     (macS_1_argbuf_d[0] ? 3'd2 :
                                      (mad1_1_argbuf_d[0] ? 3'd4 :
                                       3'd0))));
  logic [2:0] m1ad9_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad9_1_argbuf_select_q <= 3'd0;
    else
      m1ad9_1_argbuf_select_q <= (m1ad9_1_argbuf_done ? 3'd0 :
                                  m1ad9_1_argbuf_select_d);
  logic [1:0] m1ad9_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad9_1_argbuf_emit_q <= 2'd0;
    else
      m1ad9_1_argbuf_emit_q <= (m1ad9_1_argbuf_done ? 2'd0 :
                                m1ad9_1_argbuf_emit_d);
  logic [1:0] m1ad9_1_argbuf_emit_d;
  assign m1ad9_1_argbuf_emit_d = (m1ad9_1_argbuf_emit_q | ({readMerge_choice_QTree_Bool_d[0],
                                                            readMerge_data_QTree_Bool_d[0]} & {readMerge_choice_QTree_Bool_r,
                                                                                               readMerge_data_QTree_Bool_r}));
  logic m1ad9_1_argbuf_done;
  assign m1ad9_1_argbuf_done = (& m1ad9_1_argbuf_emit_d);
  assign {mad1_1_argbuf_r,
          macS_1_argbuf_r,
          m1ad9_1_argbuf_r} = (m1ad9_1_argbuf_done ? m1ad9_1_argbuf_select_d :
                               3'd0);
  assign readMerge_data_QTree_Bool_d = ((m1ad9_1_argbuf_select_d[0] && (! m1ad9_1_argbuf_emit_q[0])) ? m1ad9_1_argbuf_d :
                                        ((m1ad9_1_argbuf_select_d[1] && (! m1ad9_1_argbuf_emit_q[0])) ? macS_1_argbuf_d :
                                         ((m1ad9_1_argbuf_select_d[2] && (! m1ad9_1_argbuf_emit_q[0])) ? mad1_1_argbuf_d :
                                          {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Bool_d = ((m1ad9_1_argbuf_select_d[0] && (! m1ad9_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((m1ad9_1_argbuf_select_d[1] && (! m1ad9_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((m1ad9_1_argbuf_select_d[2] && (! m1ad9_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Bool) : (readMerge_choice_QTree_Bool,C3) (destructReadOut_QTree_Bool,QTree_Bool) > [(readPointer_QTree_Boolm1ad9_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_BoolmacS_1_argbuf,QTree_Bool),
                                                                                                    (readPointer_QTree_Boolmad1_1_argbuf,QTree_Bool)] */
  logic [2:0] destructReadOut_QTree_Bool_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Bool_d[0] && destructReadOut_QTree_Bool_d[0]))
      unique case (readMerge_choice_QTree_Bool_d[2:1])
        2'd0: destructReadOut_QTree_Bool_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Bool_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Bool_onehotd = 3'd4;
        default: destructReadOut_QTree_Bool_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Bool_onehotd = 3'd0;
  assign readPointer_QTree_Boolm1ad9_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                   destructReadOut_QTree_Bool_onehotd[0]};
  assign readPointer_QTree_BoolmacS_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                  destructReadOut_QTree_Bool_onehotd[1]};
  assign readPointer_QTree_Boolmad1_1_argbuf_d = {destructReadOut_QTree_Bool_d[66:1],
                                                  destructReadOut_QTree_Bool_onehotd[2]};
  assign destructReadOut_QTree_Bool_r = (| (destructReadOut_QTree_Bool_onehotd & {readPointer_QTree_Boolmad1_1_argbuf_r,
                                                                                  readPointer_QTree_BoolmacS_1_argbuf_r,
                                                                                  readPointer_QTree_Boolm1ad9_1_argbuf_r}));
  assign readMerge_choice_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* destruct (Ty Pointer_QTree_Bool,
          Dcon Pointer_QTree_Bool) : (readMerge_data_QTree_Bool,Pointer_QTree_Bool) > [(destructReadIn_QTree_Bool,Word16#)] */
  assign destructReadIn_QTree_Bool_d = {readMerge_data_QTree_Bool_d[16:1],
                                        readMerge_data_QTree_Bool_d[0]};
  assign readMerge_data_QTree_Bool_r = destructReadIn_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon ReadIn_QTree_Bool) : [(destructReadIn_QTree_Bool,Word16#)] > (dconReadIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconReadIn_QTree_Bool_d = ReadIn_QTree_Bool_dc((& {destructReadIn_QTree_Bool_d[0]}), destructReadIn_QTree_Bool_d);
  assign {destructReadIn_QTree_Bool_r} = {1 {(dconReadIn_QTree_Bool_r && dconReadIn_QTree_Bool_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Bool,
          Dcon ReadOut_QTree_Bool) : (memReadOut_QTree_Bool,MemOut_QTree_Bool) > [(destructReadOut_QTree_Bool,QTree_Bool)] */
  assign destructReadOut_QTree_Bool_d = {memReadOut_QTree_Bool_d[67:2],
                                         memReadOut_QTree_Bool_d[0]};
  assign memReadOut_QTree_Bool_r = destructReadOut_QTree_Bool_r;
  
  /* mergectrl (Ty C9,
           Ty QTree_Bool) : [(lizzieLet13_1_1_argbuf,QTree_Bool),
                             (lizzieLet14_1_argbuf,QTree_Bool),
                             (lizzieLet15_1_argbuf,QTree_Bool),
                             (lizzieLet17_1_argbuf,QTree_Bool),
                             (lizzieLet28_1_argbuf,QTree_Bool),
                             (lizzieLet38_1_argbuf,QTree_Bool),
                             (lizzieLet3_1_argbuf,QTree_Bool),
                             (lizzieLet5_1_argbuf,QTree_Bool),
                             (dummy_write_QTree_Bool,QTree_Bool)] > (writeMerge_choice_QTree_Bool,C9) (writeMerge_data_QTree_Bool,QTree_Bool) */
  logic [8:0] lizzieLet13_1_1_argbuf_select_d;
  assign lizzieLet13_1_1_argbuf_select_d = ((| lizzieLet13_1_1_argbuf_select_q) ? lizzieLet13_1_1_argbuf_select_q :
                                            (lizzieLet13_1_1_argbuf_d[0] ? 9'd1 :
                                             (lizzieLet14_1_argbuf_d[0] ? 9'd2 :
                                              (lizzieLet15_1_argbuf_d[0] ? 9'd4 :
                                               (lizzieLet17_1_argbuf_d[0] ? 9'd8 :
                                                (lizzieLet28_1_argbuf_d[0] ? 9'd16 :
                                                 (lizzieLet38_1_argbuf_d[0] ? 9'd32 :
                                                  (lizzieLet3_1_argbuf_d[0] ? 9'd64 :
                                                   (lizzieLet5_1_argbuf_d[0] ? 9'd128 :
                                                    (dummy_write_QTree_Bool_d[0] ? 9'd256 :
                                                     9'd0))))))))));
  logic [8:0] lizzieLet13_1_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_1_argbuf_select_q <= 9'd0;
    else
      lizzieLet13_1_1_argbuf_select_q <= (lizzieLet13_1_1_argbuf_done ? 9'd0 :
                                          lizzieLet13_1_1_argbuf_select_d);
  logic [1:0] lizzieLet13_1_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet13_1_1_argbuf_emit_q <= (lizzieLet13_1_1_argbuf_done ? 2'd0 :
                                        lizzieLet13_1_1_argbuf_emit_d);
  logic [1:0] lizzieLet13_1_1_argbuf_emit_d;
  assign lizzieLet13_1_1_argbuf_emit_d = (lizzieLet13_1_1_argbuf_emit_q | ({writeMerge_choice_QTree_Bool_d[0],
                                                                            writeMerge_data_QTree_Bool_d[0]} & {writeMerge_choice_QTree_Bool_r,
                                                                                                                writeMerge_data_QTree_Bool_r}));
  logic lizzieLet13_1_1_argbuf_done;
  assign lizzieLet13_1_1_argbuf_done = (& lizzieLet13_1_1_argbuf_emit_d);
  assign {dummy_write_QTree_Bool_r,
          lizzieLet5_1_argbuf_r,
          lizzieLet3_1_argbuf_r,
          lizzieLet38_1_argbuf_r,
          lizzieLet28_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet15_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet13_1_1_argbuf_r} = (lizzieLet13_1_1_argbuf_done ? lizzieLet13_1_1_argbuf_select_d :
                                       9'd0);
  assign writeMerge_data_QTree_Bool_d = ((lizzieLet13_1_1_argbuf_select_d[0] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet13_1_1_argbuf_d :
                                         ((lizzieLet13_1_1_argbuf_select_d[1] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                          ((lizzieLet13_1_1_argbuf_select_d[2] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                           ((lizzieLet13_1_1_argbuf_select_d[3] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                            ((lizzieLet13_1_1_argbuf_select_d[4] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet28_1_argbuf_d :
                                             ((lizzieLet13_1_1_argbuf_select_d[5] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet38_1_argbuf_d :
                                              ((lizzieLet13_1_1_argbuf_select_d[6] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet3_1_argbuf_d :
                                               ((lizzieLet13_1_1_argbuf_select_d[7] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                                ((lizzieLet13_1_1_argbuf_select_d[8] && (! lizzieLet13_1_1_argbuf_emit_q[0])) ? dummy_write_QTree_Bool_d :
                                                 {66'd0, 1'd0})))))))));
  assign writeMerge_choice_QTree_Bool_d = ((lizzieLet13_1_1_argbuf_select_d[0] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C1_9_dc(1'd1) :
                                           ((lizzieLet13_1_1_argbuf_select_d[1] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C2_9_dc(1'd1) :
                                            ((lizzieLet13_1_1_argbuf_select_d[2] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C3_9_dc(1'd1) :
                                             ((lizzieLet13_1_1_argbuf_select_d[3] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C4_9_dc(1'd1) :
                                              ((lizzieLet13_1_1_argbuf_select_d[4] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C5_9_dc(1'd1) :
                                               ((lizzieLet13_1_1_argbuf_select_d[5] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C6_9_dc(1'd1) :
                                                ((lizzieLet13_1_1_argbuf_select_d[6] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C7_9_dc(1'd1) :
                                                 ((lizzieLet13_1_1_argbuf_select_d[7] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C8_9_dc(1'd1) :
                                                  ((lizzieLet13_1_1_argbuf_select_d[8] && (! lizzieLet13_1_1_argbuf_emit_q[1])) ? C9_9_dc(1'd1) :
                                                   {4'd0, 1'd0})))))))));
  
  /* demux (Ty C9,
       Ty Pointer_QTree_Bool) : (writeMerge_choice_QTree_Bool,C9) (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool) > [(writeQTree_BoollizzieLet13_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet15_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet17_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet38_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool),
                                                                                                                      (dummy_write_QTree_Bool_sink,Pointer_QTree_Bool)] */
  logic [8:0] demuxWriteResult_QTree_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Bool_d[0] && demuxWriteResult_QTree_Bool_d[0]))
      unique case (writeMerge_choice_QTree_Bool_d[4:1])
        4'd0: demuxWriteResult_QTree_Bool_onehotd = 9'd1;
        4'd1: demuxWriteResult_QTree_Bool_onehotd = 9'd2;
        4'd2: demuxWriteResult_QTree_Bool_onehotd = 9'd4;
        4'd3: demuxWriteResult_QTree_Bool_onehotd = 9'd8;
        4'd4: demuxWriteResult_QTree_Bool_onehotd = 9'd16;
        4'd5: demuxWriteResult_QTree_Bool_onehotd = 9'd32;
        4'd6: demuxWriteResult_QTree_Bool_onehotd = 9'd64;
        4'd7: demuxWriteResult_QTree_Bool_onehotd = 9'd128;
        4'd8: demuxWriteResult_QTree_Bool_onehotd = 9'd256;
        default: demuxWriteResult_QTree_Bool_onehotd = 9'd0;
      endcase
    else demuxWriteResult_QTree_Bool_onehotd = 9'd0;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                    demuxWriteResult_QTree_Bool_onehotd[0]};
  assign writeQTree_BoollizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[1]};
  assign writeQTree_BoollizzieLet15_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[2]};
  assign writeQTree_BoollizzieLet17_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[3]};
  assign writeQTree_BoollizzieLet28_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[4]};
  assign writeQTree_BoollizzieLet38_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                  demuxWriteResult_QTree_Bool_onehotd[5]};
  assign writeQTree_BoollizzieLet3_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[6]};
  assign writeQTree_BoollizzieLet5_1_argbuf_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                                 demuxWriteResult_QTree_Bool_onehotd[7]};
  assign dummy_write_QTree_Bool_sink_d = {demuxWriteResult_QTree_Bool_d[16:1],
                                          demuxWriteResult_QTree_Bool_onehotd[8]};
  assign demuxWriteResult_QTree_Bool_r = (| (demuxWriteResult_QTree_Bool_onehotd & {dummy_write_QTree_Bool_sink_r,
                                                                                    writeQTree_BoollizzieLet5_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet3_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet38_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet28_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet17_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet15_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet14_1_argbuf_r,
                                                                                    writeQTree_BoollizzieLet13_1_1_argbuf_r}));
  assign writeMerge_choice_QTree_Bool_r = demuxWriteResult_QTree_Bool_r;
  
  /* dcon (Ty MemIn_QTree_Bool,
      Dcon WriteIn_QTree_Bool) : [(forkHP1_QTree_Boo3,Word16#),
                                  (writeMerge_data_QTree_Bool,QTree_Bool)] > (dconWriteIn_QTree_Bool,MemIn_QTree_Bool) */
  assign dconWriteIn_QTree_Bool_d = WriteIn_QTree_Bool_dc((& {forkHP1_QTree_Boo3_d[0],
                                                              writeMerge_data_QTree_Bool_d[0]}), forkHP1_QTree_Boo3_d, writeMerge_data_QTree_Bool_d);
  assign {forkHP1_QTree_Boo3_r,
          writeMerge_data_QTree_Bool_r} = {2 {(dconWriteIn_QTree_Bool_r && dconWriteIn_QTree_Bool_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Bool,
      Dcon Pointer_QTree_Bool) : [(forkHP1_QTree_Boo4,Word16#)] > (dconPtr_QTree_Bool,Pointer_QTree_Bool) */
  assign dconPtr_QTree_Bool_d = Pointer_QTree_Bool_dc((& {forkHP1_QTree_Boo4_d[0]}), forkHP1_QTree_Boo4_d);
  assign {forkHP1_QTree_Boo4_r} = {1 {(dconPtr_QTree_Bool_r && dconPtr_QTree_Bool_d[0])}};
  
  /* demux (Ty MemOut_QTree_Bool,
       Ty Pointer_QTree_Bool) : (memWriteOut_QTree_Bool,MemOut_QTree_Bool) (dconPtr_QTree_Bool,Pointer_QTree_Bool) > [(_37,Pointer_QTree_Bool),
                                                                                                                      (demuxWriteResult_QTree_Bool,Pointer_QTree_Bool)] */
  logic [1:0] dconPtr_QTree_Bool_onehotd;
  always_comb
    if ((memWriteOut_QTree_Bool_d[0] && dconPtr_QTree_Bool_d[0]))
      unique case (memWriteOut_QTree_Bool_d[1:1])
        1'd0: dconPtr_QTree_Bool_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Bool_onehotd = 2'd2;
        default: dconPtr_QTree_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Bool_onehotd = 2'd0;
  assign _37_d = {dconPtr_QTree_Bool_d[16:1],
                  dconPtr_QTree_Bool_onehotd[0]};
  assign demuxWriteResult_QTree_Bool_d = {dconPtr_QTree_Bool_d[16:1],
                                          dconPtr_QTree_Bool_onehotd[1]};
  assign dconPtr_QTree_Bool_r = (| (dconPtr_QTree_Bool_onehotd & {demuxWriteResult_QTree_Bool_r,
                                                                  _37_r}));
  assign memWriteOut_QTree_Bool_r = dconPtr_QTree_Bool_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__13,Go) > (initHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \initHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd0,
                                                    go__13_d[0]};
  assign go__13_r = \initHP_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTmap''_map''_Bool_Bool_Bool1,Go) > (incrHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd1,
                                                    \incrHP_CTmap''_map''_Bool_Bool_Bool1_d [0]};
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool1_r  = \incrHP_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* merge (Ty Go) : [(go__14,Go),
                 (incrHP_CTmap''_map''_Bool_Bool_Bool2,Go)] > (incrHP_mergeCTmap''_map''_Bool_Bool_Bool,Go) */
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ;
  always_comb
    begin
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  = 2'd0;
      if ((| \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  = \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select ;
      else
        if (go__14_d[0])
          \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [0] = 1'd1;
        else if (\incrHP_CTmap''_map''_Bool_Bool_Bool2_d [0])
          \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_select  <= (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  ? 2'd0 :
                                                            \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected );
  always_comb
    if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [0])
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = go__14_d;
    else if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected [1])
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = \incrHP_CTmap''_map''_Bool_Bool_Bool2_d ;
    else \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d  = 1'd0;
  assign {\incrHP_CTmap''_map''_Bool_Bool_Bool2_r ,
          go__14_r} = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  ? \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf,Go) > [(incrHP_CTmap''_map''_Bool_Bool_Bool1,Go),
                                                                    (incrHP_CTmap''_map''_Bool_Bool_Bool2,Go)] */
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted ;
  logic [1:0] \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done ;
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool1_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted [0]));
  assign \incrHP_CTmap''_map''_Bool_Bool_Bool2_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted [1]));
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  | ({\incrHP_CTmap''_map''_Bool_Bool_Bool2_d [0],
                                                                                                                           \incrHP_CTmap''_map''_Bool_Bool_Bool1_d [0]} & {\incrHP_CTmap''_map''_Bool_Bool_Bool2_r ,
                                                                                                                                                                           \incrHP_CTmap''_map''_Bool_Bool_Bool1_r }));
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  = (& \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_emitted  <= (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  ? 2'd0 :
                                                                 \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTmap''_map''_Bool_Bool_Bool,Word16#) (forkHP1_CTmap''_map''_Bool_Bool_Bool,Word16#) > (addHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  assign \addHP_CTmap''_map''_Bool_Bool_Bool_d  = {(\incrHP_CTmap''_map''_Bool_Bool_Bool_d [16:1] + \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [16:1]),
                                                   (\incrHP_CTmap''_map''_Bool_Bool_Bool_d [0] && \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [0])};
  assign {\incrHP_CTmap''_map''_Bool_Bool_Bool_r ,
          \forkHP1_CTmap''_map''_Bool_Bool_Bool_r } = {2 {(\addHP_CTmap''_map''_Bool_Bool_Bool_r  && \addHP_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTmap''_map''_Bool_Bool_Bool,Word16#),
                      (addHP_CTmap''_map''_Bool_Bool_Bool,Word16#)] > (mergeHP_CTmap''_map''_Bool_Bool_Bool,Word16#) */
  logic [1:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected ;
  logic [1:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ;
  always_comb
    begin
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  = 2'd0;
      if ((| \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  = \mergeHP_CTmap''_map''_Bool_Bool_Bool_select ;
      else
        if (\initHP_CTmap''_map''_Bool_Bool_Bool_d [0])
          \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [0] = 1'd1;
        else if (\addHP_CTmap''_map''_Bool_Bool_Bool_d [0])
          \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_select  <= 2'd0;
    else
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_select  <= (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r  ? 2'd0 :
                                                        \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected );
  always_comb
    if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [0])
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = \initHP_CTmap''_map''_Bool_Bool_Bool_d ;
    else if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_selected [1])
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = \addHP_CTmap''_map''_Bool_Bool_Bool_d ;
    else \mergeHP_CTmap''_map''_Bool_Bool_Bool_d  = {16'd0, 1'd0};
  assign {\addHP_CTmap''_map''_Bool_Bool_Bool_r ,
          \initHP_CTmap''_map''_Bool_Bool_Bool_r } = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r  ? \mergeHP_CTmap''_map''_Bool_Bool_Bool_selected  :
                                                      2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTmap''_map''_Bool_Bool_Bool,Go) > (incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf,Go) */
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  logic \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r ;
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r  = ((! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d [0]) || \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_r )
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d  <= \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_d ;
  Go_t \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf ;
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_r  = (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]);
  assign \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_d  = (\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0] ? \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  :
                                                             \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r  && \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_buf_r ) && (! \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf [0])))
        \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= \incrHP_mergeCTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTmap''_map''_Bool_Bool_Bool,Word16#) > (mergeHP_CTmap''_map''_Bool_Bool_Bool_buf,Word16#) */
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  logic \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r ;
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_r  = ((! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d [0]) || \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTmap''_map''_Bool_Bool_Bool_r )
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d  <= \mergeHP_CTmap''_map''_Bool_Bool_Bool_d ;
  \Word16#_t  \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf ;
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_r  = (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]);
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d  = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0] ? \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  :
                                                         \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= {16'd0,
                                                             1'd0};
    else
      if ((\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  && \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0]))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= {16'd0,
                                                               1'd0};
      else if (((! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r ) && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf [0])))
        \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_buf  <= \mergeHP_CTmap''_map''_Bool_Bool_Bool_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTmap''_map''_Bool_Bool_Bool_buf,Word16#) > [(forkHP1_CTmap''_map''_Bool_Bool_Bool,Word16#),
                                                                          (forkHP1_CTmap''_map''_Bool_Bool_Boo2,Word16#),
                                                                          (forkHP1_CTmap''_map''_Bool_Bool_Boo3,Word16#)] */
  logic [2:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted ;
  logic [2:0] \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done ;
  assign \forkHP1_CTmap''_map''_Bool_Bool_Bool_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [0]))};
  assign \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [1]))};
  assign \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d  = {\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [16:1],
                                                     (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_d [0] && (! \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted [2]))};
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done  = (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  | ({\forkHP1_CTmap''_map''_Bool_Bool_Boo3_d [0],
                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d [0],
                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_r ,
                                                                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ,
                                                                                                                                                                   \forkHP1_CTmap''_map''_Bool_Bool_Bool_r }));
  assign \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  = (& \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_emitted  <= (\mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_r  ? 3'd0 :
                                                             \mergeHP_CTmap''_map''_Bool_Bool_Bool_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : [(dconReadIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool),
                                                     (dconWriteIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool)] > (memMergeChoice_CTmap''_map''_Bool_Bool_Bool,C2) (memMergeIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d  = ((| \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q ) ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  :
                                                               (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_d [0] ? 2'd1 :
                                                                (\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d [0] ? 2'd2 :
                                                                 2'd0)));
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_q  <= (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? 2'd0 :
                                                             \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  <= 2'd0;
    else
      \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  <= (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? 2'd0 :
                                                           \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d );
  logic [1:0] \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d  = (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q  | ({\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [0],
                                                                                                                  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                                                                     \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r }));
  logic \dconReadIn_CTmap''_map''_Bool_Bool_Bool_done ;
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  = (& \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_d );
  assign {\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r ,
          \dconReadIn_CTmap''_map''_Bool_Bool_Bool_r } = (\dconReadIn_CTmap''_map''_Bool_Bool_Bool_done  ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d  :
                                                          2'd0);
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d  = ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [0] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [0])) ? \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d  :
                                                        ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [1] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [0])) ? \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d  :
                                                         {85'd0, 1'd0}));
  assign \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d  = ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [0] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [1])) ? C1_2_dc(1'd1) :
                                                            ((\dconReadIn_CTmap''_map''_Bool_Bool_Bool_select_d [1] && (! \dconReadIn_CTmap''_map''_Bool_Bool_Bool_emit_q [1])) ? C2_2_dc(1'd1) :
                                                             {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  logic [67:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ;
  logic [67:0] \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
  logic [67:0] \memOut_CTmap''_map''_Bool_Bool_Bool_q ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_valid ;
  logic \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we ;
  logic \memOut_CTmap''_map''_Bool_Bool_Bool_we ;
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din  = \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [85:18];
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address  = \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [17:2];
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we  = (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [1:1] && \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTmap''_map''_Bool_Bool_Bool_we  <= 1'd0;
        \memOut_CTmap''_map''_Bool_Bool_Bool_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTmap''_map''_Bool_Bool_Bool_we  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we ;
        \memOut_CTmap''_map''_Bool_Bool_Bool_valid  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0];
        if (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we )
          begin
            \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ] <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
            \memOut_CTmap''_map''_Bool_Bool_Bool_q  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_din ;
          end
        else
          \memOut_CTmap''_map''_Bool_Bool_Bool_q  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_mem [\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_address ];
      end
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_q ,
                                                    \memOut_CTmap''_map''_Bool_Bool_Bool_we ,
                                                    \memOut_CTmap''_map''_Bool_Bool_Bool_valid };
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r  = ((! \memOut_CTmap''_map''_Bool_Bool_Bool_valid ) || \memOut_CTmap''_map''_Bool_Bool_Bool_r );
  logic [31:0] \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read ;
  logic [31:0] \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  <= 0;
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  <= 0;
      end
    else
      if ((\memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_we  == 1'd1))
        \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  <= (\profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_write  + 1);
      else
        if ((\memOut_CTmap''_map''_Bool_Bool_Bool_valid  == 1'd1))
          \profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  <= (\profiling_MemIn_CTmap''_map''_Bool_Bool_Bool_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memMergeChoice_CTmap''_map''_Bool_Bool_Bool,C2) (memOut_CTmap''_map''_Bool_Bool_Bool_dbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) > [(memReadOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                    (memWriteOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [0] && \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]))
      unique case (\memMergeChoice_CTmap''_map''_Bool_Bool_Bool_d [1:1])
        1'd0: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd2;
        default: \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [69:1],
                                                        \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd [0]};
  assign \memWriteOut_CTmap''_map''_Bool_Bool_Bool_d  = {\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [69:1],
                                                         \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd [1]};
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r  = (| (\memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_onehotd  & {\memWriteOut_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                  \memReadOut_CTmap''_map''_Bool_Bool_Bool_r }));
  assign \memMergeChoice_CTmap''_map''_Bool_Bool_Bool_r  = \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r  = ((! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]) || \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= {85'd0, 1'd0};
    else
      if (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r )
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTmap''_map''_Bool_Bool_Bool) : (memMergeIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) > (memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  \MemIn_CTmap''_map''_Bool_Bool_Bool_t  \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf ;
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_r  = (! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0]);
  assign \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_d  = (\memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0] ? \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  :
                                                             \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= {85'd0, 1'd0};
    else
      if ((\memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r  && \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0]))
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= {85'd0, 1'd0};
      else if (((! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_rbuf_r ) && (! \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf [0])))
        \memMergeIn_CTmap''_map''_Bool_Bool_Bool_buf  <= \memMergeIn_CTmap''_map''_Bool_Bool_Bool_d ;
  
  /* dbuf (Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memOut_CTmap''_map''_Bool_Bool_Bool_rbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool_dbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r  = ((! \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d [0]) || \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= {69'd0, 1'd0};
    else
      if (\memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r )
        \memOut_CTmap''_map''_Bool_Bool_Bool_dbuf_d  <= \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTmap''_map''_Bool_Bool_Bool) : (memOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) > (memOut_CTmap''_map''_Bool_Bool_Bool_rbuf,MemOut_CTmap''_map''_Bool_Bool_Bool) */
  \MemOut_CTmap''_map''_Bool_Bool_Bool_t  \memOut_CTmap''_map''_Bool_Bool_Bool_buf ;
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_r  = (! \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0]);
  assign \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_d  = (\memOut_CTmap''_map''_Bool_Bool_Bool_buf [0] ? \memOut_CTmap''_map''_Bool_Bool_Bool_buf  :
                                                         \memOut_CTmap''_map''_Bool_Bool_Bool_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= {69'd0, 1'd0};
    else
      if ((\memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r  && \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0]))
        \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= {69'd0, 1'd0};
      else if (((! \memOut_CTmap''_map''_Bool_Bool_Bool_rbuf_r ) && (! \memOut_CTmap''_map''_Bool_Bool_Bool_buf [0])))
        \memOut_CTmap''_map''_Bool_Bool_Bool_buf  <= \memOut_CTmap''_map''_Bool_Bool_Bool_d ;
  
  /* destruct (Ty Pointer_CTmap''_map''_Bool_Bool_Bool,
          Dcon Pointer_CTmap''_map''_Bool_Bool_Bool) : (scfarg_0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(destructReadIn_CTmap''_map''_Bool_Bool_Bool,Word16#)] */
  assign \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d  = {scfarg_0_2_1_argbuf_d[16:1],
                                                            scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = \destructReadIn_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Dcon ReadIn_CTmap''_map''_Bool_Bool_Bool) : [(destructReadIn_CTmap''_map''_Bool_Bool_Bool,Word16#)] > (dconReadIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d  = \ReadIn_CTmap''_map''_Bool_Bool_Bool_dc ((& {\destructReadIn_CTmap''_map''_Bool_Bool_Bool_d [0]}), \destructReadIn_CTmap''_map''_Bool_Bool_Bool_d );
  assign {\destructReadIn_CTmap''_map''_Bool_Bool_Bool_r } = {1 {(\dconReadIn_CTmap''_map''_Bool_Bool_Bool_r  && \dconReadIn_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* destruct (Ty MemOut_CTmap''_map''_Bool_Bool_Bool,
          Dcon ReadOut_CTmap''_map''_Bool_Bool_Bool) : (memReadOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) > [(readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf,CTmap''_map''_Bool_Bool_Bool)] */
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d  = {\memReadOut_CTmap''_map''_Bool_Bool_Bool_d [69:2],
                                                                            \memReadOut_CTmap''_map''_Bool_Bool_Bool_d [0]};
  assign \memReadOut_CTmap''_map''_Bool_Bool_Bool_r  = \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTmap''_map''_Bool_Bool_Bool) : [(lizzieLet16_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet23_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet35_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet36_1_argbuf,CTmap''_map''_Bool_Bool_Bool),
                                               (lizzieLet37_1_argbuf,CTmap''_map''_Bool_Bool_Bool)] > (writeMerge_choice_CTmap''_map''_Bool_Bool_Bool,C5) (writeMerge_data_CTmap''_map''_Bool_Bool_Bool,CTmap''_map''_Bool_Bool_Bool) */
  logic [4:0] lizzieLet16_1_argbuf_select_d;
  assign lizzieLet16_1_argbuf_select_d = ((| lizzieLet16_1_argbuf_select_q) ? lizzieLet16_1_argbuf_select_q :
                                          (lizzieLet16_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet23_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet35_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet36_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet37_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet16_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet16_1_argbuf_select_q <= (lizzieLet16_1_argbuf_done ? 5'd0 :
                                        lizzieLet16_1_argbuf_select_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet16_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet16_1_argbuf_emit_q <= (lizzieLet16_1_argbuf_done ? 2'd0 :
                                      lizzieLet16_1_argbuf_emit_d);
  logic [1:0] lizzieLet16_1_argbuf_emit_d;
  assign lizzieLet16_1_argbuf_emit_d = (lizzieLet16_1_argbuf_emit_q | ({\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [0],
                                                                        \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d [0]} & {\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                                                \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r }));
  logic lizzieLet16_1_argbuf_done;
  assign lizzieLet16_1_argbuf_done = (& lizzieLet16_1_argbuf_emit_d);
  assign {lizzieLet37_1_argbuf_r,
          lizzieLet36_1_argbuf_r,
          lizzieLet35_1_argbuf_r,
          lizzieLet23_1_argbuf_r,
          lizzieLet16_1_argbuf_r} = (lizzieLet16_1_argbuf_done ? lizzieLet16_1_argbuf_select_d :
                                     5'd0);
  assign \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d  = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                                             ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet23_1_argbuf_d :
                                                              ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet35_1_argbuf_d :
                                                               ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet36_1_argbuf_d :
                                                                ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[0])) ? lizzieLet37_1_argbuf_d :
                                                                 {68'd0, 1'd0})))));
  assign \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d  = ((lizzieLet16_1_argbuf_select_d[0] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                               ((lizzieLet16_1_argbuf_select_d[1] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                                ((lizzieLet16_1_argbuf_select_d[2] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                                 ((lizzieLet16_1_argbuf_select_d[3] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                                  ((lizzieLet16_1_argbuf_select_d[4] && (! lizzieLet16_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                                   {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeMerge_choice_CTmap''_map''_Bool_Bool_Bool,C5) (demuxWriteResult_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                              (writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [4:0] \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [0] && \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [0]))
      unique case (\writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_d [3:1])
        3'd0:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd1;
        3'd1:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd2;
        3'd2:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd4;
        3'd3:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd8;
        3'd4:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd16;
        default:
          \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd0;
      endcase
    else
      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  = 5'd0;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [0]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [1]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [2]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [3]};
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_d  = {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                                      \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd [4]};
  assign \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r  = (| (\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_onehotd  & {\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_r ,
                                                                                                                            \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_r }));
  assign \writeMerge_choice_CTmap''_map''_Bool_Bool_Bool_r  = \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* dcon (Ty MemIn_CTmap''_map''_Bool_Bool_Bool,
      Dcon WriteIn_CTmap''_map''_Bool_Bool_Bool) : [(forkHP1_CTmap''_map''_Bool_Bool_Boo2,Word16#),
                                                    (writeMerge_data_CTmap''_map''_Bool_Bool_Bool,CTmap''_map''_Bool_Bool_Bool)] > (dconWriteIn_CTmap''_map''_Bool_Bool_Bool,MemIn_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d  = \WriteIn_CTmap''_map''_Bool_Bool_Bool_dc ((& {\forkHP1_CTmap''_map''_Bool_Bool_Boo2_d [0],
                                                                                                      \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d [0]}), \forkHP1_CTmap''_map''_Bool_Bool_Boo2_d , \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_d );
  assign {\forkHP1_CTmap''_map''_Bool_Bool_Boo2_r ,
          \writeMerge_data_CTmap''_map''_Bool_Bool_Bool_r } = {2 {(\dconWriteIn_CTmap''_map''_Bool_Bool_Bool_r  && \dconWriteIn_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* dcon (Ty Pointer_CTmap''_map''_Bool_Bool_Bool,
      Dcon Pointer_CTmap''_map''_Bool_Bool_Bool) : [(forkHP1_CTmap''_map''_Bool_Bool_Boo3,Word16#)] > (dconPtr_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \dconPtr_CTmap''_map''_Bool_Bool_Bool_d  = \Pointer_CTmap''_map''_Bool_Bool_Bool_dc ((& {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_d [0]}), \forkHP1_CTmap''_map''_Bool_Bool_Boo3_d );
  assign {\forkHP1_CTmap''_map''_Bool_Bool_Boo3_r } = {1 {(\dconPtr_CTmap''_map''_Bool_Bool_Bool_r  && \dconPtr_CTmap''_map''_Bool_Bool_Bool_d [0])}};
  
  /* demux (Ty MemOut_CTmap''_map''_Bool_Bool_Bool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (memWriteOut_CTmap''_map''_Bool_Bool_Bool,MemOut_CTmap''_map''_Bool_Bool_Bool) (dconPtr_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(_36,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                                                                                                (demuxWriteResult_CTmap''_map''_Bool_Bool_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd ;
  always_comb
    if ((\memWriteOut_CTmap''_map''_Bool_Bool_Bool_d [0] && \dconPtr_CTmap''_map''_Bool_Bool_Bool_d [0]))
      unique case (\memWriteOut_CTmap''_map''_Bool_Bool_Bool_d [1:1])
        1'd0: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd1;
        1'd1: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd2;
        default: \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  = 2'd0;
  assign _36_d = {\dconPtr_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                  \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd [0]};
  assign \demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_d  = {\dconPtr_CTmap''_map''_Bool_Bool_Bool_d [16:1],
                                                              \dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd [1]};
  assign \dconPtr_CTmap''_map''_Bool_Bool_Bool_r  = (| (\dconPtr_CTmap''_map''_Bool_Bool_Bool_onehotd  & {\demuxWriteResult_CTmap''_map''_Bool_Bool_Bool_r ,
                                                                                                          _36_r}));
  assign \memWriteOut_CTmap''_map''_Bool_Bool_Bool_r  = \dconPtr_CTmap''_map''_Bool_Bool_Bool_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go__15,Go) > (initHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign initHP_CTkron_kron_Bool_Bool_Bool_d = {16'd0, go__15_d[0]};
  assign go__15_r = initHP_CTkron_kron_Bool_Bool_Bool_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTkron_kron_Bool_Bool_Bool1,Go) > (incrHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign incrHP_CTkron_kron_Bool_Bool_Bool_d = {16'd1,
                                                incrHP_CTkron_kron_Bool_Bool_Bool1_d[0]};
  assign incrHP_CTkron_kron_Bool_Bool_Bool1_r = incrHP_CTkron_kron_Bool_Bool_Bool_r;
  
  /* merge (Ty Go) : [(go__16,Go),
                 (incrHP_CTkron_kron_Bool_Bool_Bool2,Go)] > (incrHP_mergeCTkron_kron_Bool_Bool_Bool,Go) */
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected;
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_select;
  always_comb
    begin
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected = 2'd0;
      if ((| incrHP_mergeCTkron_kron_Bool_Bool_Bool_select))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected = incrHP_mergeCTkron_kron_Bool_Bool_Bool_select;
      else
        if (go__16_d[0])
          incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[0] = 1'd1;
        else if (incrHP_CTkron_kron_Bool_Bool_Bool2_d[0])
          incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_select <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_select <= (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r ? 2'd0 :
                                                        incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected);
  always_comb
    if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[0])
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = go__16_d;
    else if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected[1])
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = incrHP_CTkron_kron_Bool_Bool_Bool2_d;
    else incrHP_mergeCTkron_kron_Bool_Bool_Bool_d = 1'd0;
  assign {incrHP_CTkron_kron_Bool_Bool_Bool2_r,
          go__16_r} = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r ? incrHP_mergeCTkron_kron_Bool_Bool_Bool_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf,Go) > [(incrHP_CTkron_kron_Bool_Bool_Bool1,Go),
                                                                  (incrHP_CTkron_kron_Bool_Bool_Bool2,Go)] */
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted;
  logic [1:0] incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done;
  assign incrHP_CTkron_kron_Bool_Bool_Bool1_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d[0] && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted[0]));
  assign incrHP_CTkron_kron_Bool_Bool_Bool2_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d[0] && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted[1]));
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted | ({incrHP_CTkron_kron_Bool_Bool_Bool2_d[0],
                                                                                                                   incrHP_CTkron_kron_Bool_Bool_Bool1_d[0]} & {incrHP_CTkron_kron_Bool_Bool_Bool2_r,
                                                                                                                                                               incrHP_CTkron_kron_Bool_Bool_Bool1_r}));
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r = (& incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_emitted <= (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r ? 2'd0 :
                                                             incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTkron_kron_Bool_Bool_Bool,Word16#) (forkHP1_CTkron_kron_Bool_Bool_Bool,Word16#) > (addHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  assign addHP_CTkron_kron_Bool_Bool_Bool_d = {(incrHP_CTkron_kron_Bool_Bool_Bool_d[16:1] + forkHP1_CTkron_kron_Bool_Bool_Bool_d[16:1]),
                                               (incrHP_CTkron_kron_Bool_Bool_Bool_d[0] && forkHP1_CTkron_kron_Bool_Bool_Bool_d[0])};
  assign {incrHP_CTkron_kron_Bool_Bool_Bool_r,
          forkHP1_CTkron_kron_Bool_Bool_Bool_r} = {2 {(addHP_CTkron_kron_Bool_Bool_Bool_r && addHP_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTkron_kron_Bool_Bool_Bool,Word16#),
                      (addHP_CTkron_kron_Bool_Bool_Bool,Word16#)] > (mergeHP_CTkron_kron_Bool_Bool_Bool,Word16#) */
  logic [1:0] mergeHP_CTkron_kron_Bool_Bool_Bool_selected;
  logic [1:0] mergeHP_CTkron_kron_Bool_Bool_Bool_select;
  always_comb
    begin
      mergeHP_CTkron_kron_Bool_Bool_Bool_selected = 2'd0;
      if ((| mergeHP_CTkron_kron_Bool_Bool_Bool_select))
        mergeHP_CTkron_kron_Bool_Bool_Bool_selected = mergeHP_CTkron_kron_Bool_Bool_Bool_select;
      else
        if (initHP_CTkron_kron_Bool_Bool_Bool_d[0])
          mergeHP_CTkron_kron_Bool_Bool_Bool_selected[0] = 1'd1;
        else if (addHP_CTkron_kron_Bool_Bool_Bool_d[0])
          mergeHP_CTkron_kron_Bool_Bool_Bool_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_select <= 2'd0;
    else
      mergeHP_CTkron_kron_Bool_Bool_Bool_select <= (mergeHP_CTkron_kron_Bool_Bool_Bool_r ? 2'd0 :
                                                    mergeHP_CTkron_kron_Bool_Bool_Bool_selected);
  always_comb
    if (mergeHP_CTkron_kron_Bool_Bool_Bool_selected[0])
      mergeHP_CTkron_kron_Bool_Bool_Bool_d = initHP_CTkron_kron_Bool_Bool_Bool_d;
    else if (mergeHP_CTkron_kron_Bool_Bool_Bool_selected[1])
      mergeHP_CTkron_kron_Bool_Bool_Bool_d = addHP_CTkron_kron_Bool_Bool_Bool_d;
    else mergeHP_CTkron_kron_Bool_Bool_Bool_d = {16'd0, 1'd0};
  assign {addHP_CTkron_kron_Bool_Bool_Bool_r,
          initHP_CTkron_kron_Bool_Bool_Bool_r} = (mergeHP_CTkron_kron_Bool_Bool_Bool_r ? mergeHP_CTkron_kron_Bool_Bool_Bool_selected :
                                                  2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTkron_kron_Bool_Bool_Bool,Go) > (incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf,Go) */
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d;
  logic incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r;
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_r = ((! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d[0]) || incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTkron_kron_Bool_Bool_Bool_r)
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d <= incrHP_mergeCTkron_kron_Bool_Bool_Bool_d;
  Go_t incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf;
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_r = (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0]);
  assign incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_d = (incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0] ? incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf :
                                                         incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r && incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0]))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTkron_kron_Bool_Bool_Bool_buf_r) && (! incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf[0])))
        incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_buf <= incrHP_mergeCTkron_kron_Bool_Bool_Bool_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTkron_kron_Bool_Bool_Bool,Word16#) > (mergeHP_CTkron_kron_Bool_Bool_Bool_buf,Word16#) */
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d;
  logic mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r;
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_r = ((! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d[0]) || mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTkron_kron_Bool_Bool_Bool_r)
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d <= mergeHP_CTkron_kron_Bool_Bool_Bool_d;
  \Word16#_t  mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf;
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_r = (! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0]);
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d = (mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0] ? mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf :
                                                     mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r && mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0]))
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r) && (! mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf[0])))
        mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_buf <= mergeHP_CTkron_kron_Bool_Bool_Bool_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTkron_kron_Bool_Bool_Bool_buf,Word16#) > [(forkHP1_CTkron_kron_Bool_Bool_Bool,Word16#),
                                                                        (forkHP1_CTkron_kron_Bool_Bool_Boo2,Word16#),
                                                                        (forkHP1_CTkron_kron_Bool_Bool_Boo3,Word16#)] */
  logic [2:0] mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted;
  logic [2:0] mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done;
  assign forkHP1_CTkron_kron_Bool_Bool_Bool_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[0]))};
  assign forkHP1_CTkron_kron_Bool_Bool_Boo2_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[1]))};
  assign forkHP1_CTkron_kron_Bool_Bool_Boo3_d = {mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[16:1],
                                                 (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_d[0] && (! mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted[2]))};
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done = (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted | ({forkHP1_CTkron_kron_Bool_Bool_Boo3_d[0],
                                                                                                           forkHP1_CTkron_kron_Bool_Bool_Boo2_d[0],
                                                                                                           forkHP1_CTkron_kron_Bool_Bool_Bool_d[0]} & {forkHP1_CTkron_kron_Bool_Bool_Boo3_r,
                                                                                                                                                       forkHP1_CTkron_kron_Bool_Bool_Boo2_r,
                                                                                                                                                       forkHP1_CTkron_kron_Bool_Bool_Bool_r}));
  assign mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r = (& mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted <= 3'd0;
    else
      mergeHP_CTkron_kron_Bool_Bool_Bool_buf_emitted <= (mergeHP_CTkron_kron_Bool_Bool_Bool_buf_r ? 3'd0 :
                                                         mergeHP_CTkron_kron_Bool_Bool_Bool_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTkron_kron_Bool_Bool_Bool) : [(dconReadIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool),
                                                   (dconWriteIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool)] > (memMergeChoice_CTkron_kron_Bool_Bool_Bool,C2) (memMergeIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d = ((| dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q) ? dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q :
                                                           (dconReadIn_CTkron_kron_Bool_Bool_Bool_d[0] ? 2'd1 :
                                                            (dconWriteIn_CTkron_kron_Bool_Bool_Bool_d[0] ? 2'd2 :
                                                             2'd0)));
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Bool_Bool_Bool_select_q <= (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? 2'd0 :
                                                         dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d);
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q <= 2'd0;
    else
      dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q <= (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? 2'd0 :
                                                       dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d);
  logic [1:0] dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d = (dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q | ({memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[0],
                                                                                                          memMergeIn_CTkron_kron_Bool_Bool_Bool_d[0]} & {memMergeChoice_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                                                                         memMergeIn_CTkron_kron_Bool_Bool_Bool_r}));
  logic dconReadIn_CTkron_kron_Bool_Bool_Bool_done;
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_done = (& dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_d);
  assign {dconWriteIn_CTkron_kron_Bool_Bool_Bool_r,
          dconReadIn_CTkron_kron_Bool_Bool_Bool_r} = (dconReadIn_CTkron_kron_Bool_Bool_Bool_done ? dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d :
                                                      2'd0);
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_d = ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[0] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[0])) ? dconReadIn_CTkron_kron_Bool_Bool_Bool_d :
                                                    ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[1] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[0])) ? dconWriteIn_CTkron_kron_Bool_Bool_Bool_d :
                                                     {100'd0, 1'd0}));
  assign memMergeChoice_CTkron_kron_Bool_Bool_Bool_d = ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[0] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[1])) ? C1_2_dc(1'd1) :
                                                        ((dconReadIn_CTkron_kron_Bool_Bool_Bool_select_d[1] && (! dconReadIn_CTkron_kron_Bool_Bool_Bool_emit_q[1])) ? C2_2_dc(1'd1) :
                                                         {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf,MemIn_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) */
  logic [82:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address;
  logic [82:0] memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
  logic [82:0] memOut_CTkron_kron_Bool_Bool_Bool_q;
  logic memOut_CTkron_kron_Bool_Bool_Bool_valid;
  logic memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we;
  logic memOut_CTkron_kron_Bool_Bool_Bool_we;
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din = memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[100:18];
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address = memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[17:2];
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we = (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[1:1] && memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTkron_kron_Bool_Bool_Bool_we <= 1'd0;
        memOut_CTkron_kron_Bool_Bool_Bool_valid <= 1'd0;
      end
    else
      begin
        memOut_CTkron_kron_Bool_Bool_Bool_we <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we;
        memOut_CTkron_kron_Bool_Bool_Bool_valid <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0];
        if (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we)
          begin
            memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address] <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
            memOut_CTkron_kron_Bool_Bool_Bool_q <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_din;
          end
        else
          memOut_CTkron_kron_Bool_Bool_Bool_q <= memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_mem[memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_address];
      end
  assign memOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_q,
                                                memOut_CTkron_kron_Bool_Bool_Bool_we,
                                                memOut_CTkron_kron_Bool_Bool_Bool_valid};
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r = ((! memOut_CTkron_kron_Bool_Bool_Bool_valid) || memOut_CTkron_kron_Bool_Bool_Bool_r);
  logic [31:0] profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read;
  logic [31:0] profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write <= 0;
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read <= 0;
      end
    else
      if ((memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_we == 1'd1))
        profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write <= (profiling_MemIn_CTkron_kron_Bool_Bool_Bool_write + 1);
      else
        if ((memOut_CTkron_kron_Bool_Bool_Bool_valid == 1'd1))
          profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read <= (profiling_MemIn_CTkron_kron_Bool_Bool_Bool_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memMergeChoice_CTkron_kron_Bool_Bool_Bool,C2) (memOut_CTkron_kron_Bool_Bool_Bool_dbuf,MemOut_CTkron_kron_Bool_Bool_Bool) > [(memReadOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                            (memWriteOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool)] */
  logic [1:0] memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[0] && memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]))
      unique case (memMergeChoice_CTkron_kron_Bool_Bool_Bool_d[1:1])
        1'd0: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd2;
        default: memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd = 2'd0;
  assign memReadOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[84:1],
                                                    memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd[0]};
  assign memWriteOut_CTkron_kron_Bool_Bool_Bool_d = {memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[84:1],
                                                     memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd[1]};
  assign memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r = (| (memOut_CTkron_kron_Bool_Bool_Bool_dbuf_onehotd & {memWriteOut_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                          memReadOut_CTkron_kron_Bool_Bool_Bool_r}));
  assign memMergeChoice_CTkron_kron_Bool_Bool_Bool_r = memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r;
  
  /* dbuf (Ty MemIn_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf,MemIn_CTkron_kron_Bool_Bool_Bool) > (memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r = ((! memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]) || memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d <= {100'd0, 1'd0};
    else
      if (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r)
        memMergeIn_CTkron_kron_Bool_Bool_Bool_dbuf_d <= memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  
  /* rbuf (Ty MemIn_CTkron_kron_Bool_Bool_Bool) : (memMergeIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) > (memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf,MemIn_CTkron_kron_Bool_Bool_Bool) */
  MemIn_CTkron_kron_Bool_Bool_Bool_t memMergeIn_CTkron_kron_Bool_Bool_Bool_buf;
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_r = (! memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0]);
  assign memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_d = (memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0] ? memMergeIn_CTkron_kron_Bool_Bool_Bool_buf :
                                                         memMergeIn_CTkron_kron_Bool_Bool_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= {100'd0, 1'd0};
    else
      if ((memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r && memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0]))
        memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= {100'd0, 1'd0};
      else if (((! memMergeIn_CTkron_kron_Bool_Bool_Bool_rbuf_r) && (! memMergeIn_CTkron_kron_Bool_Bool_Bool_buf[0])))
        memMergeIn_CTkron_kron_Bool_Bool_Bool_buf <= memMergeIn_CTkron_kron_Bool_Bool_Bool_d;
  
  /* dbuf (Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memOut_CTkron_kron_Bool_Bool_Bool_rbuf,MemOut_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool_dbuf,MemOut_CTkron_kron_Bool_Bool_Bool) */
  assign memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r = ((! memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d[0]) || memOut_CTkron_kron_Bool_Bool_Bool_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d <= {84'd0, 1'd0};
    else
      if (memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r)
        memOut_CTkron_kron_Bool_Bool_Bool_dbuf_d <= memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d;
  
  /* rbuf (Ty MemOut_CTkron_kron_Bool_Bool_Bool) : (memOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) > (memOut_CTkron_kron_Bool_Bool_Bool_rbuf,MemOut_CTkron_kron_Bool_Bool_Bool) */
  MemOut_CTkron_kron_Bool_Bool_Bool_t memOut_CTkron_kron_Bool_Bool_Bool_buf;
  assign memOut_CTkron_kron_Bool_Bool_Bool_r = (! memOut_CTkron_kron_Bool_Bool_Bool_buf[0]);
  assign memOut_CTkron_kron_Bool_Bool_Bool_rbuf_d = (memOut_CTkron_kron_Bool_Bool_Bool_buf[0] ? memOut_CTkron_kron_Bool_Bool_Bool_buf :
                                                     memOut_CTkron_kron_Bool_Bool_Bool_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTkron_kron_Bool_Bool_Bool_buf <= {84'd0, 1'd0};
    else
      if ((memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r && memOut_CTkron_kron_Bool_Bool_Bool_buf[0]))
        memOut_CTkron_kron_Bool_Bool_Bool_buf <= {84'd0, 1'd0};
      else if (((! memOut_CTkron_kron_Bool_Bool_Bool_rbuf_r) && (! memOut_CTkron_kron_Bool_Bool_Bool_buf[0])))
        memOut_CTkron_kron_Bool_Bool_Bool_buf <= memOut_CTkron_kron_Bool_Bool_Bool_d;
  
  /* destruct (Ty Pointer_CTkron_kron_Bool_Bool_Bool,
          Dcon Pointer_CTkron_kron_Bool_Bool_Bool) : (scfarg_0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > [(destructReadIn_CTkron_kron_Bool_Bool_Bool,Word16#)] */
  assign destructReadIn_CTkron_kron_Bool_Bool_Bool_d = {scfarg_0_1_argbuf_d[16:1],
                                                        scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CTkron_kron_Bool_Bool_Bool_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Dcon ReadIn_CTkron_kron_Bool_Bool_Bool) : [(destructReadIn_CTkron_kron_Bool_Bool_Bool,Word16#)] > (dconReadIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign dconReadIn_CTkron_kron_Bool_Bool_Bool_d = ReadIn_CTkron_kron_Bool_Bool_Bool_dc((& {destructReadIn_CTkron_kron_Bool_Bool_Bool_d[0]}), destructReadIn_CTkron_kron_Bool_Bool_Bool_d);
  assign {destructReadIn_CTkron_kron_Bool_Bool_Bool_r} = {1 {(dconReadIn_CTkron_kron_Bool_Bool_Bool_r && dconReadIn_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* destruct (Ty MemOut_CTkron_kron_Bool_Bool_Bool,
          Dcon ReadOut_CTkron_kron_Bool_Bool_Bool) : (memReadOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) > [(readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf,CTkron_kron_Bool_Bool_Bool)] */
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d = {memReadOut_CTkron_kron_Bool_Bool_Bool_d[84:2],
                                                                      memReadOut_CTkron_kron_Bool_Bool_Bool_d[0]};
  assign memReadOut_CTkron_kron_Bool_Bool_Bool_r = readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTkron_kron_Bool_Bool_Bool) : [(lizzieLet21_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet25_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet26_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet27_1_argbuf,CTkron_kron_Bool_Bool_Bool),
                                             (lizzieLet4_1_argbuf,CTkron_kron_Bool_Bool_Bool)] > (writeMerge_choice_CTkron_kron_Bool_Bool_Bool,C5) (writeMerge_data_CTkron_kron_Bool_Bool_Bool,CTkron_kron_Bool_Bool_Bool) */
  logic [4:0] lizzieLet21_1_argbuf_select_d;
  assign lizzieLet21_1_argbuf_select_d = ((| lizzieLet21_1_argbuf_select_q) ? lizzieLet21_1_argbuf_select_q :
                                          (lizzieLet21_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet25_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet26_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet27_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet4_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet21_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet21_1_argbuf_select_q <= (lizzieLet21_1_argbuf_done ? 5'd0 :
                                        lizzieLet21_1_argbuf_select_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet21_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet21_1_argbuf_emit_q <= (lizzieLet21_1_argbuf_done ? 2'd0 :
                                      lizzieLet21_1_argbuf_emit_d);
  logic [1:0] lizzieLet21_1_argbuf_emit_d;
  assign lizzieLet21_1_argbuf_emit_d = (lizzieLet21_1_argbuf_emit_q | ({writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[0],
                                                                        writeMerge_data_CTkron_kron_Bool_Bool_Bool_d[0]} & {writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                                            writeMerge_data_CTkron_kron_Bool_Bool_Bool_r}));
  logic lizzieLet21_1_argbuf_done;
  assign lizzieLet21_1_argbuf_done = (& lizzieLet21_1_argbuf_emit_d);
  assign {lizzieLet4_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet21_1_argbuf_r} = (lizzieLet21_1_argbuf_done ? lizzieLet21_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTkron_kron_Bool_Bool_Bool_d = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                                         ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                          ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                           ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                                            ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[0])) ? lizzieLet4_1_argbuf_d :
                                                             {83'd0, 1'd0})))));
  assign writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d = ((lizzieLet21_1_argbuf_select_d[0] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                           ((lizzieLet21_1_argbuf_select_d[1] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                            ((lizzieLet21_1_argbuf_select_d[2] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                             ((lizzieLet21_1_argbuf_select_d[3] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                              ((lizzieLet21_1_argbuf_select_d[4] && (! lizzieLet21_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                               {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeMerge_choice_CTkron_kron_Bool_Bool_Bool,C5) (demuxWriteResult_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > [(writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                      (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [4:0] demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd;
  always_comb
    if ((writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[0] && demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[0]))
      unique case (writeMerge_choice_CTkron_kron_Bool_Bool_Bool_d[3:1])
        3'd0: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd16;
        default:
          demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd = 5'd0;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[0]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[1]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[2]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                  demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[3]};
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_d = {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                                 demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd[4]};
  assign demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r = (| (demuxWriteResult_CTkron_kron_Bool_Bool_Bool_onehotd & {writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_r,
                                                                                                                    writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r}));
  assign writeMerge_choice_CTkron_kron_Bool_Bool_Bool_r = demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r;
  
  /* dcon (Ty MemIn_CTkron_kron_Bool_Bool_Bool,
      Dcon WriteIn_CTkron_kron_Bool_Bool_Bool) : [(forkHP1_CTkron_kron_Bool_Bool_Boo2,Word16#),
                                                  (writeMerge_data_CTkron_kron_Bool_Bool_Bool,CTkron_kron_Bool_Bool_Bool)] > (dconWriteIn_CTkron_kron_Bool_Bool_Bool,MemIn_CTkron_kron_Bool_Bool_Bool) */
  assign dconWriteIn_CTkron_kron_Bool_Bool_Bool_d = WriteIn_CTkron_kron_Bool_Bool_Bool_dc((& {forkHP1_CTkron_kron_Bool_Bool_Boo2_d[0],
                                                                                              writeMerge_data_CTkron_kron_Bool_Bool_Bool_d[0]}), forkHP1_CTkron_kron_Bool_Bool_Boo2_d, writeMerge_data_CTkron_kron_Bool_Bool_Bool_d);
  assign {forkHP1_CTkron_kron_Bool_Bool_Boo2_r,
          writeMerge_data_CTkron_kron_Bool_Bool_Bool_r} = {2 {(dconWriteIn_CTkron_kron_Bool_Bool_Bool_r && dconWriteIn_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* dcon (Ty Pointer_CTkron_kron_Bool_Bool_Bool,
      Dcon Pointer_CTkron_kron_Bool_Bool_Bool) : [(forkHP1_CTkron_kron_Bool_Bool_Boo3,Word16#)] > (dconPtr_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign dconPtr_CTkron_kron_Bool_Bool_Bool_d = Pointer_CTkron_kron_Bool_Bool_Bool_dc((& {forkHP1_CTkron_kron_Bool_Bool_Boo3_d[0]}), forkHP1_CTkron_kron_Bool_Bool_Boo3_d);
  assign {forkHP1_CTkron_kron_Bool_Bool_Boo3_r} = {1 {(dconPtr_CTkron_kron_Bool_Bool_Bool_r && dconPtr_CTkron_kron_Bool_Bool_Bool_d[0])}};
  
  /* demux (Ty MemOut_CTkron_kron_Bool_Bool_Bool,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (memWriteOut_CTkron_kron_Bool_Bool_Bool,MemOut_CTkron_kron_Bool_Bool_Bool) (dconPtr_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > [(_35,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                                                                                      (demuxWriteResult_CTkron_kron_Bool_Bool_Bool,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [1:0] dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd;
  always_comb
    if ((memWriteOut_CTkron_kron_Bool_Bool_Bool_d[0] && dconPtr_CTkron_kron_Bool_Bool_Bool_d[0]))
      unique case (memWriteOut_CTkron_kron_Bool_Bool_Bool_d[1:1])
        1'd0: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd1;
        1'd1: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd2;
        default: dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd0;
      endcase
    else dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd = 2'd0;
  assign _35_d = {dconPtr_CTkron_kron_Bool_Bool_Bool_d[16:1],
                  dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd[0]};
  assign demuxWriteResult_CTkron_kron_Bool_Bool_Bool_d = {dconPtr_CTkron_kron_Bool_Bool_Bool_d[16:1],
                                                          dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd[1]};
  assign dconPtr_CTkron_kron_Bool_Bool_Bool_r = (| (dconPtr_CTkron_kron_Bool_Bool_Bool_onehotd & {demuxWriteResult_CTkron_kron_Bool_Bool_Bool_r,
                                                                                                  _35_r}));
  assign memWriteOut_CTkron_kron_Bool_Bool_Bool_r = dconPtr_CTkron_kron_Bool_Bool_Bool_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m1adn_0,Pointer_QTree_Bool) */
  
  /* source (Ty Pointer_QTree_Bool) : > (m2ado_1,Pointer_QTree_Bool) */
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyBool,
          Dcon TupGo___MyDTBool_Bool___MyBool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) > [(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2,Go),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool),
                                                                                                                                        (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done;
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[1:1],
                                                                   (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted | ({applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0],
                                                                                                                                   applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]} & {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r,
                                                                                                                                                                                                 applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r ? 3'd0 :
                                                                     applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool) : (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0,MyDTBool_Bool) > [(arg0_1,MyDTBool_Bool),
                                                                                                  (arg0_2,MyDTBool_Bool),
                                                                                                  (arg0_3,MyDTBool_Bool)] */
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted;
  logic [2:0] applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done;
  assign arg0_1_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[0]));
  assign arg0_2_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[1]));
  assign arg0_3_d = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_d[0] && (! applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted[2]));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done = (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted | ({arg0_3_d[0],
                                                                                                                                       arg0_2_d[0],
                                                                                                                                       arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                                       arg0_2_r,
                                                                                                                                                       arg0_1_r}));
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r = (& applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= 3'd0;
    else
      applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_emitted <= (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_r ? 3'd0 :
                                                                       applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg0_done);
  
  /* fork (Ty MyBool) : (applyfnBool_Bool_5_resbuf,MyBool) > [(es_0_2_1,MyBool),
                                                         (es_0_2_2,MyBool),
                                                         (es_0_2_3,MyBool)] */
  logic [2:0] applyfnBool_Bool_5_resbuf_emitted;
  logic [2:0] applyfnBool_Bool_5_resbuf_done;
  assign es_0_2_1_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[0]))};
  assign es_0_2_2_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[1]))};
  assign es_0_2_3_d = {applyfnBool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_5_resbuf_emitted[2]))};
  assign applyfnBool_Bool_5_resbuf_done = (applyfnBool_Bool_5_resbuf_emitted | ({es_0_2_3_d[0],
                                                                                 es_0_2_2_d[0],
                                                                                 es_0_2_1_d[0]} & {es_0_2_3_r,
                                                                                                   es_0_2_2_r,
                                                                                                   es_0_2_1_r}));
  assign applyfnBool_Bool_5_resbuf_r = (& applyfnBool_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnBool_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnBool_Bool_5_resbuf_emitted <= (applyfnBool_Bool_5_resbuf_r ? 3'd0 :
                                            applyfnBool_Bool_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
          Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) > [(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4,MyDTBool_Bool_Bool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool),
                                                                                                                                                                                       (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2,MyBool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done;
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[0]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[1]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[1:1],
                                                                                      (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[2]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[2:2],
                                                                                        (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted[3]))};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted | ({applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d[0],
                                                                                                                                                                         applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]} & {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_r,
                                                                                                                                                                                                                                                          applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r ? 4'd0 :
                                                                                        applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Bool_Bool) : (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4,MyDTBool_Bool_Bool) > [(arg0_4_1,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_4_2,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_4_3,MyDTBool_Bool_Bool),
                                                                                                                                 (arg0_4_4,MyDTBool_Bool_Bool)] */
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted;
  logic [3:0] applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_done;
  assign arg0_4_1_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted[0]));
  assign arg0_4_2_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted[1]));
  assign arg0_4_3_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted[2]));
  assign arg0_4_4_d = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_d[0] && (! applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted[3]));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_done = (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted | ({arg0_4_4_d[0],
                                                                                                                                                                                 arg0_4_3_d[0],
                                                                                                                                                                                 arg0_4_2_d[0],
                                                                                                                                                                                 arg0_4_1_d[0]} & {arg0_4_4_r,
                                                                                                                                                                                                   arg0_4_3_r,
                                                                                                                                                                                                   arg0_4_2_r,
                                                                                                                                                                                                   arg0_4_1_r}));
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_r = (& applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted <= 4'd0;
    else
      applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_emitted <= (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_r ? 4'd0 :
                                                                                            applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg0_4_done);
  
  /* fork (Ty MyBool) : (applyfnBool_Bool_Bool_5_resbuf,MyBool) > [(xacw_1_1,MyBool),
                                                              (xacw_1_2,MyBool)] */
  logic [1:0] applyfnBool_Bool_Bool_5_resbuf_emitted;
  logic [1:0] applyfnBool_Bool_Bool_5_resbuf_done;
  assign xacw_1_1_d = {applyfnBool_Bool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_Bool_5_resbuf_emitted[0]))};
  assign xacw_1_2_d = {applyfnBool_Bool_Bool_5_resbuf_d[1:1],
                       (applyfnBool_Bool_Bool_5_resbuf_d[0] && (! applyfnBool_Bool_Bool_5_resbuf_emitted[1]))};
  assign applyfnBool_Bool_Bool_5_resbuf_done = (applyfnBool_Bool_Bool_5_resbuf_emitted | ({xacw_1_2_d[0],
                                                                                           xacw_1_1_d[0]} & {xacw_1_2_r,
                                                                                                             xacw_1_1_r}));
  assign applyfnBool_Bool_Bool_5_resbuf_r = (& applyfnBool_Bool_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Bool_Bool_5_resbuf_emitted <= 2'd0;
    else
      applyfnBool_Bool_Bool_5_resbuf_emitted <= (applyfnBool_Bool_Bool_5_resbuf_r ? 2'd0 :
                                                 applyfnBool_Bool_Bool_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTBool_Nat___MyBool,
          Dcon TupGo___MyDTBool_Nat___MyBool) : (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1,TupGo___MyDTBool_Nat___MyBool) > [(applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4,Go),
                                                                                                                                    (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2,MyDTBool_Nat),
                                                                                                                                    (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1,MyBool)] */
  logic [2:0] applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted;
  logic [2:0] applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_done;
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted[0]));
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted[1]));
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d = {applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d[1:1],
                                                                   (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted[2]))};
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_done = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted | ({applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d[0],
                                                                                                                               applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d[0],
                                                                                                                               applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d[0]} & {applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_r,
                                                                                                                                                                                           applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_r,
                                                                                                                                                                                           applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_r}));
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_r = (& applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted <= 3'd0;
    else
      applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_emitted <= (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_r ? 3'd0 :
                                                                   applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_done);
  
  /* fork (Ty MyDTBool_Nat) : (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2,MyDTBool_Nat) > [(arg0_2_1,MyDTBool_Nat),
                                                                                                (arg0_2_2,MyDTBool_Nat),
                                                                                                (arg0_2_3,MyDTBool_Nat)] */
  logic [2:0] applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted;
  logic [2:0] applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_done;
  assign arg0_2_1_d = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_d[0] && (! applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted[2]));
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_done = (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                                       arg0_2_2_d[0],
                                                                                                                                       arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                                         arg0_2_2_r,
                                                                                                                                                         arg0_2_1_r}));
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_r = (& applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted <= 3'd0;
    else
      applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_emitted <= (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_r ? 3'd0 :
                                                                       applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg0_2_done);
  
  /* fork (Ty Pointer_Nat) : (applyfnBool_Nat_5_resbuf,Pointer_Nat) > [(xacw_1,Pointer_Nat),
                                                                  (xacw_2,Pointer_Nat)] */
  logic [1:0] applyfnBool_Nat_5_resbuf_emitted;
  logic [1:0] applyfnBool_Nat_5_resbuf_done;
  assign xacw_1_d = {applyfnBool_Nat_5_resbuf_d[16:1],
                     (applyfnBool_Nat_5_resbuf_d[0] && (! applyfnBool_Nat_5_resbuf_emitted[0]))};
  assign xacw_2_d = {applyfnBool_Nat_5_resbuf_d[16:1],
                     (applyfnBool_Nat_5_resbuf_d[0] && (! applyfnBool_Nat_5_resbuf_emitted[1]))};
  assign applyfnBool_Nat_5_resbuf_done = (applyfnBool_Nat_5_resbuf_emitted | ({xacw_2_d[0],
                                                                               xacw_1_d[0]} & {xacw_2_r,
                                                                                               xacw_1_r}));
  assign applyfnBool_Nat_5_resbuf_r = (& applyfnBool_Nat_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnBool_Nat_5_resbuf_emitted <= 2'd0;
    else
      applyfnBool_Nat_5_resbuf_emitted <= (applyfnBool_Nat_5_resbuf_r ? 2'd0 :
                                           applyfnBool_Nat_5_resbuf_done);
  
  /* destruct (Ty TupGo___MyDTNat_Bool___Pointer_Nat,
          Dcon TupGo___MyDTNat_Bool___Pointer_Nat) : (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1,TupGo___MyDTNat_Bool___Pointer_Nat) > [(applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5,Go),
                                                                                                                                                   (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6,MyDTNat_Bool),
                                                                                                                                                   (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3,Pointer_Nat)] */
  logic [2:0] applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted;
  logic [2:0] applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_done;
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted[0]));
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted[1]));
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d = {applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d[16:1],
                                                                        (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted[2]))};
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_done = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted | ({applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d[0],
                                                                                                                                         applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d[0],
                                                                                                                                         applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d[0]} & {applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_r,
                                                                                                                                                                                                          applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_r,
                                                                                                                                                                                                          applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_r}));
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_r = (& applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted <= 3'd0;
    else
      applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_emitted <= (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_r ? 3'd0 :
                                                                        applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_done);
  
  /* fork (Ty MyDTNat_Bool) : (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6,MyDTNat_Bool) > [(arg0_6_1,MyDTNat_Bool),
                                                                                                     (arg0_6_2,MyDTNat_Bool),
                                                                                                     (arg0_6_3,MyDTNat_Bool)] */
  logic [2:0] applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted;
  logic [2:0] applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_done;
  assign arg0_6_1_d = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted[0]));
  assign arg0_6_2_d = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted[1]));
  assign arg0_6_3_d = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_d[0] && (! applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted[2]));
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_done = (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted | ({arg0_6_3_d[0],
                                                                                                                                                 arg0_6_2_d[0],
                                                                                                                                                 arg0_6_1_d[0]} & {arg0_6_3_r,
                                                                                                                                                                   arg0_6_2_r,
                                                                                                                                                                   arg0_6_1_r}));
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_r = (& applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted <= 3'd0;
    else
      applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_emitted <= (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_r ? 3'd0 :
                                                                            applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg0_6_done);
  
  /* fork (Ty MyBool) : (applyfnNat_Bool_5_resbuf,MyBool) > [(es_0_1_1,MyBool),
                                                        (es_0_1_2,MyBool),
                                                        (es_0_1_3,MyBool)] */
  logic [2:0] applyfnNat_Bool_5_resbuf_emitted;
  logic [2:0] applyfnNat_Bool_5_resbuf_done;
  assign es_0_1_1_d = {applyfnNat_Bool_5_resbuf_d[1:1],
                       (applyfnNat_Bool_5_resbuf_d[0] && (! applyfnNat_Bool_5_resbuf_emitted[0]))};
  assign es_0_1_2_d = {applyfnNat_Bool_5_resbuf_d[1:1],
                       (applyfnNat_Bool_5_resbuf_d[0] && (! applyfnNat_Bool_5_resbuf_emitted[1]))};
  assign es_0_1_3_d = {applyfnNat_Bool_5_resbuf_d[1:1],
                       (applyfnNat_Bool_5_resbuf_d[0] && (! applyfnNat_Bool_5_resbuf_emitted[2]))};
  assign applyfnNat_Bool_5_resbuf_done = (applyfnNat_Bool_5_resbuf_emitted | ({es_0_1_3_d[0],
                                                                               es_0_1_2_d[0],
                                                                               es_0_1_1_d[0]} & {es_0_1_3_r,
                                                                                                 es_0_1_2_r,
                                                                                                 es_0_1_1_r}));
  assign applyfnNat_Bool_5_resbuf_r = (& applyfnNat_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnNat_Bool_5_resbuf_emitted <= 3'd0;
    else
      applyfnNat_Bool_5_resbuf_emitted <= (applyfnNat_Bool_5_resbuf_r ? 3'd0 :
                                           applyfnNat_Bool_5_resbuf_done);
  
  /* demux (Ty MyDTBool_Bool,
       Ty MyBool) : (arg0_1,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1,MyBool) > [(arg0_1Dcon_main1,MyBool)] */
  assign arg0_1Dcon_main1_d = {applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[1:1],
                               (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0])};
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_main1_r && (arg0_1_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolarg1_d[0]));
  
  /* fork (Ty MyBool) : (arg0_1Dcon_main1,MyBool) > [(arg0_1Dcon_main1_1,MyBool),
                                                (arg0_1Dcon_main1_2,MyBool)] */
  logic [1:0] arg0_1Dcon_main1_emitted;
  logic [1:0] arg0_1Dcon_main1_done;
  assign arg0_1Dcon_main1_1_d = {arg0_1Dcon_main1_d[1:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[0]))};
  assign arg0_1Dcon_main1_2_d = {arg0_1Dcon_main1_d[1:1],
                                 (arg0_1Dcon_main1_d[0] && (! arg0_1Dcon_main1_emitted[1]))};
  assign arg0_1Dcon_main1_done = (arg0_1Dcon_main1_emitted | ({arg0_1Dcon_main1_2_d[0],
                                                               arg0_1Dcon_main1_1_d[0]} & {arg0_1Dcon_main1_2_r,
                                                                                           arg0_1Dcon_main1_1_r}));
  assign arg0_1Dcon_main1_r = (& arg0_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_main1_emitted <= 2'd0;
    else
      arg0_1Dcon_main1_emitted <= (arg0_1Dcon_main1_r ? 2'd0 :
                                   arg0_1Dcon_main1_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_1Dcon_main1_1,MyBool) (arg0_2Dcon_main1,Go) > [(arg0_1Dcon_main1_1MyFalse,Go),
                                                                     (arg0_1Dcon_main1_1MyTrue,Go)] */
  logic [1:0] arg0_2Dcon_main1_onehotd;
  always_comb
    if ((arg0_1Dcon_main1_1_d[0] && arg0_2Dcon_main1_d[0]))
      unique case (arg0_1Dcon_main1_1_d[1:1])
        1'd0: arg0_2Dcon_main1_onehotd = 2'd1;
        1'd1: arg0_2Dcon_main1_onehotd = 2'd2;
        default: arg0_2Dcon_main1_onehotd = 2'd0;
      endcase
    else arg0_2Dcon_main1_onehotd = 2'd0;
  assign arg0_1Dcon_main1_1MyFalse_d = arg0_2Dcon_main1_onehotd[0];
  assign arg0_1Dcon_main1_1MyTrue_d = arg0_2Dcon_main1_onehotd[1];
  assign arg0_2Dcon_main1_r = (| (arg0_2Dcon_main1_onehotd & {arg0_1Dcon_main1_1MyTrue_r,
                                                              arg0_1Dcon_main1_1MyFalse_r}));
  assign arg0_1Dcon_main1_1_r = arg0_2Dcon_main1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(arg0_1Dcon_main1_1MyFalse,Go)] > (arg0_1Dcon_main1_1MyFalse_1MyTrue,MyBool) */
  assign arg0_1Dcon_main1_1MyFalse_1MyTrue_d = MyTrue_dc((& {arg0_1Dcon_main1_1MyFalse_d[0]}), arg0_1Dcon_main1_1MyFalse_d);
  assign {arg0_1Dcon_main1_1MyFalse_r} = {1 {(arg0_1Dcon_main1_1MyFalse_1MyTrue_r && arg0_1Dcon_main1_1MyFalse_1MyTrue_d[0])}};
  
  /* buf (Ty MyBool) : (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux,MyBool) > (applyfnBool_Bool_5_resbuf,MyBool) */
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  logic arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r;
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r = ((! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d[0]) || arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d <= {1'd0,
                                                                                               1'd0};
    else
      if (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r)
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d <= arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d;
  MyBool_t arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf;
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_r = (! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]);
  assign applyfnBool_Bool_5_resbuf_d = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0] ? arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf :
                                        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                 1'd0};
    else
      if ((applyfnBool_Bool_5_resbuf_r && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0]))
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= {1'd0,
                                                                                                   1'd0};
      else if (((! applyfnBool_Bool_5_resbuf_r) && (! arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf[0])))
        arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_buf <= arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(arg0_1Dcon_main1_1MyTrue,Go)] > (arg0_1Dcon_main1_1MyTrue_1MyFalse,MyBool) */
  assign arg0_1Dcon_main1_1MyTrue_1MyFalse_d = MyFalse_dc((& {arg0_1Dcon_main1_1MyTrue_d[0]}), arg0_1Dcon_main1_1MyTrue_d);
  assign {arg0_1Dcon_main1_1MyTrue_r} = {1 {(arg0_1Dcon_main1_1MyTrue_1MyFalse_r && arg0_1Dcon_main1_1MyTrue_1MyFalse_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_1Dcon_main1_2,MyBool) [(arg0_1Dcon_main1_1MyFalse_1MyTrue,MyBool),
                                               (arg0_1Dcon_main1_1MyTrue_1MyFalse,MyBool)] > (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux,MyBool) */
  logic [1:0] arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux;
  logic [1:0] arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot;
  always_comb
    unique case (arg0_1Dcon_main1_2_d[1:1])
      1'd0:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd1,
                                                                                        arg0_1Dcon_main1_1MyFalse_1MyTrue_d};
      1'd1:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd2,
                                                                                        arg0_1Dcon_main1_1MyTrue_1MyFalse_d};
      default:
        {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot,
         arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux} = {2'd0,
                                                                                        {1'd0,
                                                                                         1'd0}};
    endcase
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d = {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux[1:1],
                                                                                     (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux[0] && arg0_1Dcon_main1_2_d[0])};
  assign arg0_1Dcon_main1_2_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r);
  assign {arg0_1Dcon_main1_1MyTrue_1MyFalse_r,
          arg0_1Dcon_main1_1MyFalse_1MyTrue_r} = (arg0_1Dcon_main1_2_r ? arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_onehot :
                                                  2'd0);
  
  /* demux (Ty MyDTBool_Bool,
       Ty Go) : (arg0_2,MyDTBool_Bool) (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2,Go) > [(arg0_2Dcon_main1,Go)] */
  assign arg0_2Dcon_main1_d = (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]);
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]));
  assign arg0_2_r = (arg0_2Dcon_main1_r && (arg0_2_d[0] && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBoolgo_2_d[0]));
  
  /* demux (Ty MyDTBool_Nat,
       Ty MyBool) : (arg0_2_1,MyDTBool_Nat) (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1,MyBool) > [(arg0_2_1Dcon_to_nat,MyBool)] */
  assign arg0_2_1Dcon_to_nat_d = {applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d[1:1],
                                  (arg0_2_1_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d[0])};
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_r = (arg0_2_1Dcon_to_nat_r && (arg0_2_1_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d[0]));
  assign arg0_2_1_r = (arg0_2_1Dcon_to_nat_r && (arg0_2_1_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolarg1_1_d[0]));
  
  /* fork (Ty MyBool) : (arg0_2_1Dcon_to_nat,MyBool) > [(arg0_2_1Dcon_to_nat_1,MyBool),
                                                   (arg0_2_1Dcon_to_nat_2,MyBool)] */
  logic [1:0] arg0_2_1Dcon_to_nat_emitted;
  logic [1:0] arg0_2_1Dcon_to_nat_done;
  assign arg0_2_1Dcon_to_nat_1_d = {arg0_2_1Dcon_to_nat_d[1:1],
                                    (arg0_2_1Dcon_to_nat_d[0] && (! arg0_2_1Dcon_to_nat_emitted[0]))};
  assign arg0_2_1Dcon_to_nat_2_d = {arg0_2_1Dcon_to_nat_d[1:1],
                                    (arg0_2_1Dcon_to_nat_d[0] && (! arg0_2_1Dcon_to_nat_emitted[1]))};
  assign arg0_2_1Dcon_to_nat_done = (arg0_2_1Dcon_to_nat_emitted | ({arg0_2_1Dcon_to_nat_2_d[0],
                                                                     arg0_2_1Dcon_to_nat_1_d[0]} & {arg0_2_1Dcon_to_nat_2_r,
                                                                                                    arg0_2_1Dcon_to_nat_1_r}));
  assign arg0_2_1Dcon_to_nat_r = (& arg0_2_1Dcon_to_nat_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_to_nat_emitted <= 2'd0;
    else
      arg0_2_1Dcon_to_nat_emitted <= (arg0_2_1Dcon_to_nat_r ? 2'd0 :
                                      arg0_2_1Dcon_to_nat_done);
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_2_1Dcon_to_nat_1,MyBool) (arg0_2_2Dcon_to_nat,Go) > [(arg0_2_1Dcon_to_nat_1MyFalse,Go),
                                                                           (arg0_2_1Dcon_to_nat_1MyTrue,Go)] */
  logic [1:0] arg0_2_2Dcon_to_nat_onehotd;
  always_comb
    if ((arg0_2_1Dcon_to_nat_1_d[0] && arg0_2_2Dcon_to_nat_d[0]))
      unique case (arg0_2_1Dcon_to_nat_1_d[1:1])
        1'd0: arg0_2_2Dcon_to_nat_onehotd = 2'd1;
        1'd1: arg0_2_2Dcon_to_nat_onehotd = 2'd2;
        default: arg0_2_2Dcon_to_nat_onehotd = 2'd0;
      endcase
    else arg0_2_2Dcon_to_nat_onehotd = 2'd0;
  assign arg0_2_1Dcon_to_nat_1MyFalse_d = arg0_2_2Dcon_to_nat_onehotd[0];
  assign arg0_2_1Dcon_to_nat_1MyTrue_d = arg0_2_2Dcon_to_nat_onehotd[1];
  assign arg0_2_2Dcon_to_nat_r = (| (arg0_2_2Dcon_to_nat_onehotd & {arg0_2_1Dcon_to_nat_1MyTrue_r,
                                                                    arg0_2_1Dcon_to_nat_1MyFalse_r}));
  assign arg0_2_1Dcon_to_nat_1_r = arg0_2_2Dcon_to_nat_r;
  
  /* dcon (Ty Nat,
      Dcon Zero) : [(arg0_2_1Dcon_to_nat_1MyFalse,Go)] > (arg0_2_1Dcon_to_nat_1MyFalse_1Zero,Nat) */
  assign arg0_2_1Dcon_to_nat_1MyFalse_1Zero_d = Zero_dc((& {arg0_2_1Dcon_to_nat_1MyFalse_d[0]}), arg0_2_1Dcon_to_nat_1MyFalse_d);
  assign {arg0_2_1Dcon_to_nat_1MyFalse_r} = {1 {(arg0_2_1Dcon_to_nat_1MyFalse_1Zero_r && arg0_2_1Dcon_to_nat_1MyFalse_1Zero_d[0])}};
  
  /* buf (Ty Nat) : (arg0_2_1Dcon_to_nat_1MyFalse_1Zero,Nat) > (lizzieLet0_1_argbuf,Nat) */
  Nat_t arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d;
  logic arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_r;
  assign arg0_2_1Dcon_to_nat_1MyFalse_1Zero_r = ((! arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d[0]) || arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d <= {17'd0, 1'd0};
    else
      if (arg0_2_1Dcon_to_nat_1MyFalse_1Zero_r)
        arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d <= arg0_2_1Dcon_to_nat_1MyFalse_1Zero_d;
  Nat_t arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf;
  assign arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_r = (! arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf[0] ? arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf :
                                  arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf[0]))
        arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf <= {17'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf[0])))
        arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_buf <= arg0_2_1Dcon_to_nat_1MyFalse_1Zero_bufchan_d;
  
  /* buf (Ty Go) : (arg0_2_1Dcon_to_nat_1MyTrue,Go) > (arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf,Go) */
  Go_t arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d;
  logic arg0_2_1Dcon_to_nat_1MyTrue_bufchan_r;
  assign arg0_2_1Dcon_to_nat_1MyTrue_r = ((! arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d[0]) || arg0_2_1Dcon_to_nat_1MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d <= 1'd0;
    else
      if (arg0_2_1Dcon_to_nat_1MyTrue_r)
        arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d <= arg0_2_1Dcon_to_nat_1MyTrue_d;
  Go_t arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf;
  assign arg0_2_1Dcon_to_nat_1MyTrue_bufchan_r = (! arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf[0]);
  assign arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_d = (arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf[0] ? arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf :
                                                   arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf <= 1'd0;
    else
      if ((arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_r && arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf[0]))
        arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf <= 1'd0;
      else if (((! arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_r) && (! arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf[0])))
        arg0_2_1Dcon_to_nat_1MyTrue_bufchan_buf <= arg0_2_1Dcon_to_nat_1MyTrue_bufchan_d;
  
  /* dcon (Ty TupGo,
      Dcon TupGo) : [(arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf,Go)] > (to_nat1TupGo_1,TupGo) */
  assign to_nat1TupGo_1_d = TupGo_dc((& {arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_d[0]}), arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_d);
  assign {arg0_2_1Dcon_to_nat_1MyTrue_1_argbuf_r} = {1 {(to_nat1TupGo_1_r && to_nat1TupGo_1_d[0])}};
  
  /* mux (Ty MyBool,
     Ty Pointer_Nat) : (arg0_2_1Dcon_to_nat_2,MyBool) [(writeNatlizzieLet0_1_argbuf_rwb,Pointer_Nat),
                                                       (to_nat1_resbuf,Pointer_Nat)] > (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux,Pointer_Nat) */
  logic [16:0] writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux;
  logic [1:0] writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_onehot;
  always_comb
    unique case (arg0_2_1Dcon_to_nat_2_d[1:1])
      1'd0:
        {writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_onehot,
         writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux} = {2'd1,
                                                                   writeNatlizzieLet0_1_argbuf_rwb_d};
      1'd1:
        {writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_onehot,
         writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux} = {2'd2,
                                                                   to_nat1_resbuf_d};
      default:
        {writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_onehot,
         writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux} = {2'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d = {writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux[16:1],
                                                                (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux[0] && arg0_2_1Dcon_to_nat_2_d[0])};
  assign arg0_2_1Dcon_to_nat_2_r = (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d[0] && writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_r);
  assign {to_nat1_resbuf_r,
          writeNatlizzieLet0_1_argbuf_rwb_r} = (arg0_2_1Dcon_to_nat_2_r ? writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_onehot :
                                                2'd0);
  
  /* demux (Ty MyDTBool_Nat,
       Ty Go) : (arg0_2_2,MyDTBool_Nat) (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4,Go) > [(arg0_2_2Dcon_to_nat,Go)] */
  assign arg0_2_2Dcon_to_nat_d = (arg0_2_2_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d[0]);
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_r = (arg0_2_2Dcon_to_nat_r && (arg0_2_2_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d[0]));
  assign arg0_2_2_r = (arg0_2_2Dcon_to_nat_r && (arg0_2_2_d[0] && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBoolgo_4_d[0]));
  
  /* mux (Ty MyDTBool_Nat,
     Ty Pointer_Nat) : (arg0_2_3,MyDTBool_Nat) [(writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux,Pointer_Nat)] > (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux,Pointer_Nat) */
  assign writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_d = {writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d[16:1],
                                                                    (arg0_2_3_d[0] && writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d[0])};
  assign writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_r = (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_r && (arg0_2_3_d[0] && writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d[0]));
  assign arg0_2_3_r = (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_r && (arg0_2_3_d[0] && writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_d[0]));
  
  /* mux (Ty MyDTBool_Bool,
     Ty MyBool) : (arg0_3,MyDTBool_Bool) [(arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux,MyBool)] > (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux,MyBool) */
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_d = {arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[1:1],
                                                                                         (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0])};
  assign arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0]));
  assign arg0_3_r = (arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_mux_r && (arg0_3_d[0] && arg0_1Dcon_main1_1MyFalse_1MyTruearg0_1Dcon_main1_1MyTrue_1MyFalse_mux_d[0]));
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_4_1,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2,MyBool) > [(arg0_4_1Dcon_&&,MyBool)] */
  assign \arg0_4_1Dcon_&&_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d[1:1],
                                (arg0_4_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_r = (\arg0_4_1Dcon_&&_r  && (arg0_4_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d[0]));
  assign arg0_4_1_r = (\arg0_4_1Dcon_&&_r  && (arg0_4_1_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg1_2_d[0]));
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty MyBool) : (arg0_4_2,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2,MyBool) > [(arg0_4_2Dcon_&&,MyBool)] */
  assign \arg0_4_2Dcon_&&_d  = {applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[1:1],
                                (arg0_4_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0])};
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_r = (\arg0_4_2Dcon_&&_r  && (arg0_4_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  assign arg0_4_2_r = (\arg0_4_2Dcon_&&_r  && (arg0_4_2_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolarg2_d[0]));
  
  /* fork (Ty MyBool) : (arg0_4_2Dcon_&&,MyBool) > [(arg0_4_2Dcon_&&_1,MyBool),
                                               (arg0_4_2Dcon_&&_2,MyBool),
                                               (arg0_4_2Dcon_&&_3,MyBool)] */
  logic [2:0] \arg0_4_2Dcon_&&_emitted ;
  logic [2:0] \arg0_4_2Dcon_&&_done ;
  assign \arg0_4_2Dcon_&&_1_d  = {\arg0_4_2Dcon_&&_d [1:1],
                                  (\arg0_4_2Dcon_&&_d [0] && (! \arg0_4_2Dcon_&&_emitted [0]))};
  assign \arg0_4_2Dcon_&&_2_d  = {\arg0_4_2Dcon_&&_d [1:1],
                                  (\arg0_4_2Dcon_&&_d [0] && (! \arg0_4_2Dcon_&&_emitted [1]))};
  assign \arg0_4_2Dcon_&&_3_d  = {\arg0_4_2Dcon_&&_d [1:1],
                                  (\arg0_4_2Dcon_&&_d [0] && (! \arg0_4_2Dcon_&&_emitted [2]))};
  assign \arg0_4_2Dcon_&&_done  = (\arg0_4_2Dcon_&&_emitted  | ({\arg0_4_2Dcon_&&_3_d [0],
                                                                 \arg0_4_2Dcon_&&_2_d [0],
                                                                 \arg0_4_2Dcon_&&_1_d [0]} & {\arg0_4_2Dcon_&&_3_r ,
                                                                                              \arg0_4_2Dcon_&&_2_r ,
                                                                                              \arg0_4_2Dcon_&&_1_r }));
  assign \arg0_4_2Dcon_&&_r  = (& \arg0_4_2Dcon_&&_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_4_2Dcon_&&_emitted  <= 3'd0;
    else
      \arg0_4_2Dcon_&&_emitted  <= (\arg0_4_2Dcon_&&_r  ? 3'd0 :
                                    \arg0_4_2Dcon_&&_done );
  
  /* demux (Ty MyBool,
       Ty MyBool) : (arg0_4_2Dcon_&&_1,MyBool) (arg0_4_1Dcon_&&,MyBool) > [(_34,MyBool),
                                                                           (arg0_4_2Dcon_&&_1MyTrue,MyBool)] */
  logic [1:0] \arg0_4_1Dcon_&&_onehotd ;
  always_comb
    if ((\arg0_4_2Dcon_&&_1_d [0] && \arg0_4_1Dcon_&&_d [0]))
      unique case (\arg0_4_2Dcon_&&_1_d [1:1])
        1'd0: \arg0_4_1Dcon_&&_onehotd  = 2'd1;
        1'd1: \arg0_4_1Dcon_&&_onehotd  = 2'd2;
        default: \arg0_4_1Dcon_&&_onehotd  = 2'd0;
      endcase
    else \arg0_4_1Dcon_&&_onehotd  = 2'd0;
  assign _34_d = {\arg0_4_1Dcon_&&_d [1:1],
                  \arg0_4_1Dcon_&&_onehotd [0]};
  assign \arg0_4_2Dcon_&&_1MyTrue_d  = {\arg0_4_1Dcon_&&_d [1:1],
                                        \arg0_4_1Dcon_&&_onehotd [1]};
  assign \arg0_4_1Dcon_&&_r  = (| (\arg0_4_1Dcon_&&_onehotd  & {\arg0_4_2Dcon_&&_1MyTrue_r ,
                                                                _34_r}));
  assign \arg0_4_2Dcon_&&_1_r  = \arg0_4_1Dcon_&&_r ;
  
  /* demux (Ty MyBool,
       Ty Go) : (arg0_4_2Dcon_&&_2,MyBool) (arg0_4_3Dcon_&&,Go) > [(arg0_4_2Dcon_&&_2MyFalse,Go),
                                                                   (_33,Go)] */
  logic [1:0] \arg0_4_3Dcon_&&_onehotd ;
  always_comb
    if ((\arg0_4_2Dcon_&&_2_d [0] && \arg0_4_3Dcon_&&_d [0]))
      unique case (\arg0_4_2Dcon_&&_2_d [1:1])
        1'd0: \arg0_4_3Dcon_&&_onehotd  = 2'd1;
        1'd1: \arg0_4_3Dcon_&&_onehotd  = 2'd2;
        default: \arg0_4_3Dcon_&&_onehotd  = 2'd0;
      endcase
    else \arg0_4_3Dcon_&&_onehotd  = 2'd0;
  assign \arg0_4_2Dcon_&&_2MyFalse_d  = \arg0_4_3Dcon_&&_onehotd [0];
  assign _33_d = \arg0_4_3Dcon_&&_onehotd [1];
  assign \arg0_4_3Dcon_&&_r  = (| (\arg0_4_3Dcon_&&_onehotd  & {_33_r,
                                                                \arg0_4_2Dcon_&&_2MyFalse_r }));
  assign \arg0_4_2Dcon_&&_2_r  = \arg0_4_3Dcon_&&_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(arg0_4_2Dcon_&&_2MyFalse,Go)] > (arg0_4_2Dcon_&&_2MyFalse_1MyFalse,MyBool) */
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_d  = MyFalse_dc((& {\arg0_4_2Dcon_&&_2MyFalse_d [0]}), \arg0_4_2Dcon_&&_2MyFalse_d );
  assign {\arg0_4_2Dcon_&&_2MyFalse_r } = {1 {(\arg0_4_2Dcon_&&_2MyFalse_1MyFalse_r  && \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_d [0])}};
  
  /* buf (Ty MyBool) : (arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux,MyBool) > (applyfnBool_Bool_Bool_5_resbuf,MyBool) */
  MyBool_t \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d ;
  logic \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r ;
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_r  = ((! \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d [0]) || \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d  <= {1'd0,
                                                                                         1'd0};
    else
      if (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_r )
        \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d  <= \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_d ;
  MyBool_t \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf ;
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_r  = (! \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0]);
  assign applyfnBool_Bool_Bool_5_resbuf_d = (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0] ? \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  :
                                             \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= {1'd0,
                                                                                           1'd0};
    else
      if ((applyfnBool_Bool_Bool_5_resbuf_r && \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0]))
        \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= {1'd0,
                                                                                             1'd0};
      else if (((! applyfnBool_Bool_Bool_5_resbuf_r) && (! \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf [0])))
        \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_buf  <= \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_bufchan_d ;
  
  /* mux (Ty MyBool,
     Ty MyBool) : (arg0_4_2Dcon_&&_3,MyBool) [(arg0_4_2Dcon_&&_2MyFalse_1MyFalse,MyBool),
                                              (arg0_4_2Dcon_&&_1MyTrue,MyBool)] > (arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux,MyBool) */
  logic [1:0] \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux ;
  logic [1:0] \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_onehot ;
  always_comb
    unique case (\arg0_4_2Dcon_&&_3_d [1:1])
      1'd0:
        {\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd1,
                                                                                  \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_d };
      1'd1:
        {\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd2,
                                                                                  \arg0_4_2Dcon_&&_1MyTrue_d };
      default:
        {\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_onehot ,
         \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux } = {2'd0,
                                                                                  {1'd0, 1'd0}};
    endcase
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d  = {\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux [1:1],
                                                                               (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux [0] && \arg0_4_2Dcon_&&_3_d [0])};
  assign \arg0_4_2Dcon_&&_3_r  = (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d [0] && \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_r );
  assign {\arg0_4_2Dcon_&&_1MyTrue_r ,
          \arg0_4_2Dcon_&&_2MyFalse_1MyFalse_r } = (\arg0_4_2Dcon_&&_3_r  ? \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_onehot  :
                                                    2'd0);
  
  /* demux (Ty MyDTBool_Bool_Bool,
       Ty Go) : (arg0_4_3,MyDTBool_Bool_Bool) (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3,Go) > [(arg0_4_3Dcon_&&,Go)] */
  assign \arg0_4_3Dcon_&&_d  = (arg0_4_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]);
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_r = (\arg0_4_3Dcon_&&_r  && (arg0_4_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  assign arg0_4_3_r = (\arg0_4_3Dcon_&&_r  && (arg0_4_3_d[0] && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBoolgo_3_d[0]));
  
  /* mux (Ty MyDTBool_Bool_Bool,
     Ty MyBool) : (arg0_4_4,MyDTBool_Bool_Bool) [(arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux,MyBool)] > (arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux,MyBool) */
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_d  = {\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d [1:1],
                                                                                   (arg0_4_4_d[0] && \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d [0])};
  assign \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_r  = (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_r  && (arg0_4_4_d[0] && \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d [0]));
  assign arg0_4_4_r = (\arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_mux_r  && (arg0_4_4_d[0] && \arg0_4_2Dcon_&&_2MyFalse_1MyFalsearg0_4_2Dcon_&&_1MyTrue_1_mux_d [0]));
  
  /* demux (Ty MyDTNat_Bool,
       Ty Pointer_Nat) : (arg0_6_1,MyDTNat_Bool) (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3,Pointer_Nat) > [(arg0_6_1Dcon_is_z_nut,Pointer_Nat)] */
  assign arg0_6_1Dcon_is_z_nut_d = {applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d[16:1],
                                    (arg0_6_1_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d[0])};
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_r = (arg0_6_1Dcon_is_z_nut_r && (arg0_6_1_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d[0]));
  assign arg0_6_1_r = (arg0_6_1Dcon_is_z_nut_r && (arg0_6_1_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natarg1_3_d[0]));
  
  /* buf (Ty Pointer_Nat) : (arg0_6_1Dcon_is_z_nut,Pointer_Nat) > (arg0_6_1Dcon_is_z_nut_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t arg0_6_1Dcon_is_z_nut_bufchan_d;
  logic arg0_6_1Dcon_is_z_nut_bufchan_r;
  assign arg0_6_1Dcon_is_z_nut_r = ((! arg0_6_1Dcon_is_z_nut_bufchan_d[0]) || arg0_6_1Dcon_is_z_nut_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_6_1Dcon_is_z_nut_bufchan_d <= {16'd0, 1'd0};
    else
      if (arg0_6_1Dcon_is_z_nut_r)
        arg0_6_1Dcon_is_z_nut_bufchan_d <= arg0_6_1Dcon_is_z_nut_d;
  Pointer_Nat_t arg0_6_1Dcon_is_z_nut_bufchan_buf;
  assign arg0_6_1Dcon_is_z_nut_bufchan_r = (! arg0_6_1Dcon_is_z_nut_bufchan_buf[0]);
  assign arg0_6_1Dcon_is_z_nut_1_argbuf_d = (arg0_6_1Dcon_is_z_nut_bufchan_buf[0] ? arg0_6_1Dcon_is_z_nut_bufchan_buf :
                                             arg0_6_1Dcon_is_z_nut_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_6_1Dcon_is_z_nut_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((arg0_6_1Dcon_is_z_nut_1_argbuf_r && arg0_6_1Dcon_is_z_nut_bufchan_buf[0]))
        arg0_6_1Dcon_is_z_nut_bufchan_buf <= {16'd0, 1'd0};
      else if (((! arg0_6_1Dcon_is_z_nut_1_argbuf_r) && (! arg0_6_1Dcon_is_z_nut_bufchan_buf[0])))
        arg0_6_1Dcon_is_z_nut_bufchan_buf <= arg0_6_1Dcon_is_z_nut_bufchan_d;
  
  /* demux (Ty MyDTNat_Bool,
       Ty Go) : (arg0_6_2,MyDTNat_Bool) (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5,Go) > [(arg0_6_2Dcon_is_z_nut,Go)] */
  assign arg0_6_2Dcon_is_z_nut_d = (arg0_6_2_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d[0]);
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_r = (arg0_6_2Dcon_is_z_nut_r && (arg0_6_2_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d[0]));
  assign arg0_6_2_r = (arg0_6_2Dcon_is_z_nut_r && (arg0_6_2_d[0] && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Natgo_5_d[0]));
  
  /* fork (Ty Go) : (arg0_6_2Dcon_is_z_nut,Go) > [(arg0_6_2Dcon_is_z_nut_1,Go),
                                             (arg0_6_2Dcon_is_z_nut_2,Go)] */
  logic [1:0] arg0_6_2Dcon_is_z_nut_emitted;
  logic [1:0] arg0_6_2Dcon_is_z_nut_done;
  assign arg0_6_2Dcon_is_z_nut_1_d = (arg0_6_2Dcon_is_z_nut_d[0] && (! arg0_6_2Dcon_is_z_nut_emitted[0]));
  assign arg0_6_2Dcon_is_z_nut_2_d = (arg0_6_2Dcon_is_z_nut_d[0] && (! arg0_6_2Dcon_is_z_nut_emitted[1]));
  assign arg0_6_2Dcon_is_z_nut_done = (arg0_6_2Dcon_is_z_nut_emitted | ({arg0_6_2Dcon_is_z_nut_2_d[0],
                                                                         arg0_6_2Dcon_is_z_nut_1_d[0]} & {arg0_6_2Dcon_is_z_nut_2_r,
                                                                                                          arg0_6_2Dcon_is_z_nut_1_r}));
  assign arg0_6_2Dcon_is_z_nut_r = (& arg0_6_2Dcon_is_z_nut_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_6_2Dcon_is_z_nut_emitted <= 2'd0;
    else
      arg0_6_2Dcon_is_z_nut_emitted <= (arg0_6_2Dcon_is_z_nut_r ? 2'd0 :
                                        arg0_6_2Dcon_is_z_nut_done);
  
  /* dcon (Ty Nat,
      Dcon Zero) : [(arg0_6_2Dcon_is_z_nut_1,Go)] > (arg0_6_2Dcon_is_z_nut_1Zero,Nat) */
  assign arg0_6_2Dcon_is_z_nut_1Zero_d = Zero_dc((& {arg0_6_2Dcon_is_z_nut_1_d[0]}), arg0_6_2Dcon_is_z_nut_1_d);
  assign {arg0_6_2Dcon_is_z_nut_1_r} = {1 {(arg0_6_2Dcon_is_z_nut_1Zero_r && arg0_6_2Dcon_is_z_nut_1Zero_d[0])}};
  
  /* buf (Ty Nat) : (arg0_6_2Dcon_is_z_nut_1Zero,Nat) > (lizzieLet1_1_argbuf,Nat) */
  Nat_t arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d;
  logic arg0_6_2Dcon_is_z_nut_1Zero_bufchan_r;
  assign arg0_6_2Dcon_is_z_nut_1Zero_r = ((! arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d[0]) || arg0_6_2Dcon_is_z_nut_1Zero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d <= {17'd0, 1'd0};
    else
      if (arg0_6_2Dcon_is_z_nut_1Zero_r)
        arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d <= arg0_6_2Dcon_is_z_nut_1Zero_d;
  Nat_t arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf;
  assign arg0_6_2Dcon_is_z_nut_1Zero_bufchan_r = (! arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf[0]);
  assign lizzieLet1_1_argbuf_d = (arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf[0] ? arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf :
                                  arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((lizzieLet1_1_argbuf_r && arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf[0]))
        arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf <= {17'd0, 1'd0};
      else if (((! lizzieLet1_1_argbuf_r) && (! arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf[0])))
        arg0_6_2Dcon_is_z_nut_1Zero_bufchan_buf <= arg0_6_2Dcon_is_z_nut_1Zero_bufchan_d;
  
  /* buf (Ty Go) : (arg0_6_2Dcon_is_z_nut_2,Go) > (arg0_6_2Dcon_is_z_nut_2_argbuf,Go) */
  Go_t arg0_6_2Dcon_is_z_nut_2_bufchan_d;
  logic arg0_6_2Dcon_is_z_nut_2_bufchan_r;
  assign arg0_6_2Dcon_is_z_nut_2_r = ((! arg0_6_2Dcon_is_z_nut_2_bufchan_d[0]) || arg0_6_2Dcon_is_z_nut_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_6_2Dcon_is_z_nut_2_bufchan_d <= 1'd0;
    else
      if (arg0_6_2Dcon_is_z_nut_2_r)
        arg0_6_2Dcon_is_z_nut_2_bufchan_d <= arg0_6_2Dcon_is_z_nut_2_d;
  Go_t arg0_6_2Dcon_is_z_nut_2_bufchan_buf;
  assign arg0_6_2Dcon_is_z_nut_2_bufchan_r = (! arg0_6_2Dcon_is_z_nut_2_bufchan_buf[0]);
  assign arg0_6_2Dcon_is_z_nut_2_argbuf_d = (arg0_6_2Dcon_is_z_nut_2_bufchan_buf[0] ? arg0_6_2Dcon_is_z_nut_2_bufchan_buf :
                                             arg0_6_2Dcon_is_z_nut_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_6_2Dcon_is_z_nut_2_bufchan_buf <= 1'd0;
    else
      if ((arg0_6_2Dcon_is_z_nut_2_argbuf_r && arg0_6_2Dcon_is_z_nut_2_bufchan_buf[0]))
        arg0_6_2Dcon_is_z_nut_2_bufchan_buf <= 1'd0;
      else if (((! arg0_6_2Dcon_is_z_nut_2_argbuf_r) && (! arg0_6_2Dcon_is_z_nut_2_bufchan_buf[0])))
        arg0_6_2Dcon_is_z_nut_2_bufchan_buf <= arg0_6_2Dcon_is_z_nut_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_Nat___Pointer_Nat,
      Dcon TupGo___Pointer_Nat___Pointer_Nat) : [(arg0_6_2Dcon_is_z_nut_2_argbuf,Go),
                                                 (arg0_6_1Dcon_is_z_nut_1_argbuf,Pointer_Nat),
                                                 (es_1_1_1_argbuf,Pointer_Nat)] > (eqNatTupGo___Pointer_Nat___Pointer_Nat_1,TupGo___Pointer_Nat___Pointer_Nat) */
  assign eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d = TupGo___Pointer_Nat___Pointer_Nat_dc((& {arg0_6_2Dcon_is_z_nut_2_argbuf_d[0],
                                                                                               arg0_6_1Dcon_is_z_nut_1_argbuf_d[0],
                                                                                               es_1_1_1_argbuf_d[0]}), arg0_6_2Dcon_is_z_nut_2_argbuf_d, arg0_6_1Dcon_is_z_nut_1_argbuf_d, es_1_1_1_argbuf_d);
  assign {arg0_6_2Dcon_is_z_nut_2_argbuf_r,
          arg0_6_1Dcon_is_z_nut_1_argbuf_r,
          es_1_1_1_argbuf_r} = {3 {(eqNatTupGo___Pointer_Nat___Pointer_Nat_1_r && eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[0])}};
  
  /* mux (Ty MyDTNat_Bool,
     Ty MyBool) : (arg0_6_3,MyDTNat_Bool) [(lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2,MyBool)] > (eqNat_1_mux,MyBool) */
  assign eqNat_1_mux_d = {lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d[1:1],
                          (arg0_6_3_d[0] && lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d[0])};
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_r = (eqNat_1_mux_r && (arg0_6_3_d[0] && lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d[0]));
  assign arg0_6_3_r = (eqNat_1_mux_r && (arg0_6_3_d[0] && lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d[0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) : (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) > [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                    (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [5:0] call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted;
  logic [5:0] call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done;
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[0]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[1]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[2]));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[16:1],
                                                                                                                                                                          (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[3]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[32:17],
                                                                                                                                                                          (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[4]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[48:33],
                                                                                                                                                                         (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0] && (! call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted[5]))};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done = (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted | ({call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d[0],
                                                                                                                                                                                                                                                                                                                                               call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d[0]} & {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_r}));
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r = (& call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted <= 6'd0;
    else
      call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_emitted <= (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r ? 6'd0 :
                                                                                                                                                                           call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_done);
  
  /* rbuf (Ty Go) : (call_kron_kron_Bool_Bool_Bool_goConst,Go) > (call_kron_kron_Bool_Bool_Bool_initBufi,Go) */
  Go_t call_kron_kron_Bool_Bool_Bool_goConst_buf;
  assign call_kron_kron_Bool_Bool_Bool_goConst_r = (! call_kron_kron_Bool_Bool_Bool_goConst_buf[0]);
  assign call_kron_kron_Bool_Bool_Bool_initBufi_d = (call_kron_kron_Bool_Bool_Bool_goConst_buf[0] ? call_kron_kron_Bool_Bool_Bool_goConst_buf :
                                                     call_kron_kron_Bool_Bool_Bool_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goConst_buf <= 1'd0;
    else
      if ((call_kron_kron_Bool_Bool_Bool_initBufi_r && call_kron_kron_Bool_Bool_Bool_goConst_buf[0]))
        call_kron_kron_Bool_Bool_Bool_goConst_buf <= 1'd0;
      else if (((! call_kron_kron_Bool_Bool_Bool_initBufi_r) && (! call_kron_kron_Bool_Bool_Bool_goConst_buf[0])))
        call_kron_kron_Bool_Bool_Bool_goConst_buf <= call_kron_kron_Bool_Bool_Bool_goConst_d;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_kron_kron_Bool_Bool_Bool_goMux1,Go),
                     (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf,Go),
                     (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf,Go),
                     (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf,Go),
                     (lizzieLet2_4QNode_Bool_1_argbuf,Go)] > (go_6_goMux_choice,C5) (go_6_goMux_data,Go) */
  logic [4:0] call_kron_kron_Bool_Bool_Bool_goMux1_select_d;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_select_d = ((| call_kron_kron_Bool_Bool_Bool_goMux1_select_q) ? call_kron_kron_Bool_Bool_Bool_goMux1_select_q :
                                                          (call_kron_kron_Bool_Bool_Bool_goMux1_d[0] ? 5'd1 :
                                                           (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d[0] ? 5'd2 :
                                                            (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d[0] ? 5'd4 :
                                                             (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d[0] ? 5'd8 :
                                                              (lizzieLet2_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                               5'd0))))));
  logic [4:0] call_kron_kron_Bool_Bool_Bool_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goMux1_select_q <= 5'd0;
    else
      call_kron_kron_Bool_Bool_Bool_goMux1_select_q <= (call_kron_kron_Bool_Bool_Bool_goMux1_done ? 5'd0 :
                                                        call_kron_kron_Bool_Bool_Bool_goMux1_select_d);
  logic [1:0] call_kron_kron_Bool_Bool_Bool_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_goMux1_emit_q <= 2'd0;
    else
      call_kron_kron_Bool_Bool_Bool_goMux1_emit_q <= (call_kron_kron_Bool_Bool_Bool_goMux1_done ? 2'd0 :
                                                      call_kron_kron_Bool_Bool_Bool_goMux1_emit_d);
  logic [1:0] call_kron_kron_Bool_Bool_Bool_goMux1_emit_d;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_emit_d = (call_kron_kron_Bool_Bool_Bool_goMux1_emit_q | ({go_6_goMux_choice_d[0],
                                                                                                        go_6_goMux_data_d[0]} & {go_6_goMux_choice_r,
                                                                                                                                 go_6_goMux_data_r}));
  logic call_kron_kron_Bool_Bool_Bool_goMux1_done;
  assign call_kron_kron_Bool_Bool_Bool_goMux1_done = (& call_kron_kron_Bool_Bool_Bool_goMux1_emit_d);
  assign {lizzieLet2_4QNode_Bool_1_argbuf_r,
          lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r,
          lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r,
          lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux1_r} = (call_kron_kron_Bool_Bool_Bool_goMux1_done ? call_kron_kron_Bool_Bool_Bool_goMux1_select_d :
                                                     5'd0);
  assign go_6_goMux_data_d = ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[0] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? call_kron_kron_Bool_Bool_Bool_goMux1_d :
                              ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[1] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d :
                               ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[2] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d :
                                ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[3] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d :
                                 ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[4] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[0])) ? lizzieLet2_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_6_goMux_choice_d = ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[0] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[1] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                 ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[2] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                  ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[3] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                   ((call_kron_kron_Bool_Bool_Bool_goMux1_select_d[4] && (! call_kron_kron_Bool_Bool_Bool_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_kron_kron_Bool_Bool_Bool_initBuf,Go) > [(call_kron_kron_Bool_Bool_Bool_unlockFork1,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork2,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork3,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork4,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork5,Go),
                                                             (call_kron_kron_Bool_Bool_Bool_unlockFork6,Go)] */
  logic [5:0] call_kron_kron_Bool_Bool_Bool_initBuf_emitted;
  logic [5:0] call_kron_kron_Bool_Bool_Bool_initBuf_done;
  assign call_kron_kron_Bool_Bool_Bool_unlockFork1_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork2_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[1]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork3_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[2]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork4_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[3]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork5_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[4]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork6_d = (call_kron_kron_Bool_Bool_Bool_initBuf_d[0] && (! call_kron_kron_Bool_Bool_Bool_initBuf_emitted[5]));
  assign call_kron_kron_Bool_Bool_Bool_initBuf_done = (call_kron_kron_Bool_Bool_Bool_initBuf_emitted | ({call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0],
                                                                                                         call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0]} & {call_kron_kron_Bool_Bool_Bool_unlockFork6_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork5_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork4_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork3_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork2_r,
                                                                                                                                                            call_kron_kron_Bool_Bool_Bool_unlockFork1_r}));
  assign call_kron_kron_Bool_Bool_Bool_initBuf_r = (& call_kron_kron_Bool_Bool_Bool_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_initBuf_emitted <= 6'd0;
    else
      call_kron_kron_Bool_Bool_Bool_initBuf_emitted <= (call_kron_kron_Bool_Bool_Bool_initBuf_r ? 6'd0 :
                                                        call_kron_kron_Bool_Bool_Bool_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_kron_kron_Bool_Bool_Bool_initBufi,Go) > (call_kron_kron_Bool_Bool_Bool_initBuf,Go) */
  assign call_kron_kron_Bool_Bool_Bool_initBufi_r = ((! call_kron_kron_Bool_Bool_Bool_initBuf_d[0]) || call_kron_kron_Bool_Bool_Bool_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_kron_kron_Bool_Bool_Bool_initBuf_d <= Go_dc(1'd1);
    else
      if (call_kron_kron_Bool_Bool_Bool_initBufi_r)
        call_kron_kron_Bool_Bool_Bool_initBuf_d <= call_kron_kron_Bool_Bool_Bool_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_kron_kron_Bool_Bool_Bool_unlockFork1,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6,Go)] > (call_kron_kron_Bool_Bool_Bool_goMux1,Go) */
  assign call_kron_kron_Bool_Bool_Bool_goMux1_d = (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_r = (call_kron_kron_Bool_Bool_Bool_goMux1_r && (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork1_r = (call_kron_kron_Bool_Bool_Bool_goMux1_r && (call_kron_kron_Bool_Bool_Bool_unlockFork1_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgo_6_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork2,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7,MyDTBool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux2,MyDTBool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux2_d = (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_r = (call_kron_kron_Bool_Bool_Bool_goMux2_r && (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork2_r = (call_kron_kron_Bool_Bool_Bool_goMux2_r && (call_kron_kron_Bool_Bool_Bool_unlockFork2_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_BoolisZad7_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork3,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8,MyDTBool_Bool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux3_d = (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d[0]);
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_r = (call_kron_kron_Bool_Bool_Bool_goMux3_r && (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork3_r = (call_kron_kron_Bool_Bool_Bool_goMux3_r && (call_kron_kron_Bool_Bool_Bool_unlockFork3_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolgad8_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork4,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9,Pointer_QTree_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux4,Pointer_QTree_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux4_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_r = (call_kron_kron_Bool_Bool_Bool_goMux4_r && (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork4_r = (call_kron_kron_Bool_Bool_Bool_goMux4_r && (call_kron_kron_Bool_Bool_Bool_unlockFork4_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm1ad9_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork5,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada,Pointer_QTree_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux5_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_r = (call_kron_kron_Bool_Bool_Bool_goMux5_r && (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork5_r = (call_kron_kron_Bool_Bool_Bool_goMux5_r && (call_kron_kron_Bool_Bool_Bool_unlockFork5_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolm2ada_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (call_kron_kron_Bool_Bool_Bool_unlockFork6,Go) [(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0,Pointer_CTkron_kron_Bool_Bool_Bool)] > (call_kron_kron_Bool_Bool_Bool_goMux6,Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_Bool_goMux6_d = {call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[16:1],
                                                   (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0])};
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_r = (call_kron_kron_Bool_Bool_Bool_goMux6_r && (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0]));
  assign call_kron_kron_Bool_Bool_Bool_unlockFork6_r = (call_kron_kron_Bool_Bool_Bool_goMux6_r && (call_kron_kron_Bool_Bool_Bool_unlockFork6_d[0] && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Boolsc_0_d[0]));
  
  /* destruct (Ty TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat,
          Dcon TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat) : (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1,TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat) > [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7,Go),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ,MyDTNat_Bool),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR,MyDTBool_Nat),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                        (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1,Pointer_CTmain_map'_Bool_Nat)] */
  logic [4:0] \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted ;
  logic [4:0] \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_done ;
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d  = (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0] && (! \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted [0]));
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d  = (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0] && (! \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted [1]));
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d  = (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0] && (! \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted [2]));
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d  = {\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [16:1],
                                                                                                                                   (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0] && (! \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted [3]))};
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d  = {\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [32:17],
                                                                                                                                     (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0] && (! \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted [4]))};
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_done  = (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted  | ({\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d [0],
                                                                                                                                                                                                                                                                   \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d [0]} & {\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                 \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_r ,
                                                                                                                                                                                                                                                                                                                                                                                                 \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_r ,
                                                                                                                                                                                                                                                                                                                                                                                                 \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_r ,
                                                                                                                                                                                                                                                                                                                                                                                                 \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_r }));
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_r  = (& \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted  <= 5'd0;
    else
      \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_emitted  <= (\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_r  ? 5'd0 :
                                                                                                                                     \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_done );
  
  /* rbuf (Ty Go) : (call_main_map'_Bool_Nat_goConst,Go) > (call_main_map'_Bool_Nat_initBufi,Go) */
  Go_t \call_main_map'_Bool_Nat_goConst_buf ;
  assign \call_main_map'_Bool_Nat_goConst_r  = (! \call_main_map'_Bool_Nat_goConst_buf [0]);
  assign \call_main_map'_Bool_Nat_initBufi_d  = (\call_main_map'_Bool_Nat_goConst_buf [0] ? \call_main_map'_Bool_Nat_goConst_buf  :
                                                 \call_main_map'_Bool_Nat_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \call_main_map'_Bool_Nat_goConst_buf  <= 1'd0;
    else
      if ((\call_main_map'_Bool_Nat_initBufi_r  && \call_main_map'_Bool_Nat_goConst_buf [0]))
        \call_main_map'_Bool_Nat_goConst_buf  <= 1'd0;
      else if (((! \call_main_map'_Bool_Nat_initBufi_r ) && (! \call_main_map'_Bool_Nat_goConst_buf [0])))
        \call_main_map'_Bool_Nat_goConst_buf  <= \call_main_map'_Bool_Nat_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_main_map'_Bool_Nat_goMux1,Go),
                           (lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf,Go),
                           (lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf,Go),
                           (lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf,Go),
                           (lizzieLet6_4QNode_Bool_1_argbuf,Go)] > (go_7_goMux_choice,C5) (go_7_goMux_data,Go) */
  logic [4:0] \call_main_map'_Bool_Nat_goMux1_select_d ;
  assign \call_main_map'_Bool_Nat_goMux1_select_d  = ((| \call_main_map'_Bool_Nat_goMux1_select_q ) ? \call_main_map'_Bool_Nat_goMux1_select_q  :
                                                      (\call_main_map'_Bool_Nat_goMux1_d [0] ? 5'd1 :
                                                       (\lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_d [0] ? 5'd2 :
                                                        (\lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_d [0] ? 5'd4 :
                                                         (\lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_d [0] ? 5'd8 :
                                                          (lizzieLet6_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                           5'd0))))));
  logic [4:0] \call_main_map'_Bool_Nat_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Bool_Nat_goMux1_select_q  <= 5'd0;
    else
      \call_main_map'_Bool_Nat_goMux1_select_q  <= (\call_main_map'_Bool_Nat_goMux1_done  ? 5'd0 :
                                                    \call_main_map'_Bool_Nat_goMux1_select_d );
  logic [1:0] \call_main_map'_Bool_Nat_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Bool_Nat_goMux1_emit_q  <= 2'd0;
    else
      \call_main_map'_Bool_Nat_goMux1_emit_q  <= (\call_main_map'_Bool_Nat_goMux1_done  ? 2'd0 :
                                                  \call_main_map'_Bool_Nat_goMux1_emit_d );
  logic [1:0] \call_main_map'_Bool_Nat_goMux1_emit_d ;
  assign \call_main_map'_Bool_Nat_goMux1_emit_d  = (\call_main_map'_Bool_Nat_goMux1_emit_q  | ({go_7_goMux_choice_d[0],
                                                                                                go_7_goMux_data_d[0]} & {go_7_goMux_choice_r,
                                                                                                                         go_7_goMux_data_r}));
  logic \call_main_map'_Bool_Nat_goMux1_done ;
  assign \call_main_map'_Bool_Nat_goMux1_done  = (& \call_main_map'_Bool_Nat_goMux1_emit_d );
  assign {lizzieLet6_4QNode_Bool_1_argbuf_r,
          \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_r ,
          \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_r ,
          \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_r ,
          \call_main_map'_Bool_Nat_goMux1_r } = (\call_main_map'_Bool_Nat_goMux1_done  ? \call_main_map'_Bool_Nat_goMux1_select_d  :
                                                 5'd0);
  assign go_7_goMux_data_d = ((\call_main_map'_Bool_Nat_goMux1_select_d [0] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [0])) ? \call_main_map'_Bool_Nat_goMux1_d  :
                              ((\call_main_map'_Bool_Nat_goMux1_select_d [1] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [0])) ? \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_d  :
                               ((\call_main_map'_Bool_Nat_goMux1_select_d [2] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [0])) ? \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_d  :
                                ((\call_main_map'_Bool_Nat_goMux1_select_d [3] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [0])) ? \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_d  :
                                 ((\call_main_map'_Bool_Nat_goMux1_select_d [4] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [0])) ? lizzieLet6_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_7_goMux_choice_d = ((\call_main_map'_Bool_Nat_goMux1_select_d [0] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_main_map'_Bool_Nat_goMux1_select_d [1] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_main_map'_Bool_Nat_goMux1_select_d [2] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_main_map'_Bool_Nat_goMux1_select_d [3] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_main_map'_Bool_Nat_goMux1_select_d [4] && (! \call_main_map'_Bool_Nat_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_main_map'_Bool_Nat_initBuf,Go) > [(call_main_map'_Bool_Nat_unlockFork1,Go),
                                                       (call_main_map'_Bool_Nat_unlockFork2,Go),
                                                       (call_main_map'_Bool_Nat_unlockFork3,Go),
                                                       (call_main_map'_Bool_Nat_unlockFork4,Go),
                                                       (call_main_map'_Bool_Nat_unlockFork5,Go)] */
  logic [4:0] \call_main_map'_Bool_Nat_initBuf_emitted ;
  logic [4:0] \call_main_map'_Bool_Nat_initBuf_done ;
  assign \call_main_map'_Bool_Nat_unlockFork1_d  = (\call_main_map'_Bool_Nat_initBuf_d [0] && (! \call_main_map'_Bool_Nat_initBuf_emitted [0]));
  assign \call_main_map'_Bool_Nat_unlockFork2_d  = (\call_main_map'_Bool_Nat_initBuf_d [0] && (! \call_main_map'_Bool_Nat_initBuf_emitted [1]));
  assign \call_main_map'_Bool_Nat_unlockFork3_d  = (\call_main_map'_Bool_Nat_initBuf_d [0] && (! \call_main_map'_Bool_Nat_initBuf_emitted [2]));
  assign \call_main_map'_Bool_Nat_unlockFork4_d  = (\call_main_map'_Bool_Nat_initBuf_d [0] && (! \call_main_map'_Bool_Nat_initBuf_emitted [3]));
  assign \call_main_map'_Bool_Nat_unlockFork5_d  = (\call_main_map'_Bool_Nat_initBuf_d [0] && (! \call_main_map'_Bool_Nat_initBuf_emitted [4]));
  assign \call_main_map'_Bool_Nat_initBuf_done  = (\call_main_map'_Bool_Nat_initBuf_emitted  | ({\call_main_map'_Bool_Nat_unlockFork5_d [0],
                                                                                                 \call_main_map'_Bool_Nat_unlockFork4_d [0],
                                                                                                 \call_main_map'_Bool_Nat_unlockFork3_d [0],
                                                                                                 \call_main_map'_Bool_Nat_unlockFork2_d [0],
                                                                                                 \call_main_map'_Bool_Nat_unlockFork1_d [0]} & {\call_main_map'_Bool_Nat_unlockFork5_r ,
                                                                                                                                                \call_main_map'_Bool_Nat_unlockFork4_r ,
                                                                                                                                                \call_main_map'_Bool_Nat_unlockFork3_r ,
                                                                                                                                                \call_main_map'_Bool_Nat_unlockFork2_r ,
                                                                                                                                                \call_main_map'_Bool_Nat_unlockFork1_r }));
  assign \call_main_map'_Bool_Nat_initBuf_r  = (& \call_main_map'_Bool_Nat_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Bool_Nat_initBuf_emitted  <= 5'd0;
    else
      \call_main_map'_Bool_Nat_initBuf_emitted  <= (\call_main_map'_Bool_Nat_initBuf_r  ? 5'd0 :
                                                    \call_main_map'_Bool_Nat_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_main_map'_Bool_Nat_initBufi,Go) > (call_main_map'_Bool_Nat_initBuf,Go) */
  assign \call_main_map'_Bool_Nat_initBufi_r  = ((! \call_main_map'_Bool_Nat_initBuf_d [0]) || \call_main_map'_Bool_Nat_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_main_map'_Bool_Nat_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_main_map'_Bool_Nat_initBufi_r )
        \call_main_map'_Bool_Nat_initBuf_d  <= \call_main_map'_Bool_Nat_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_main_map'_Bool_Nat_unlockFork1,Go) [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7,Go)] > (call_main_map'_Bool_Nat_goMux1,Go) */
  assign \call_main_map'_Bool_Nat_goMux1_d  = (\call_main_map'_Bool_Nat_unlockFork1_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d [0]);
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_r  = (\call_main_map'_Bool_Nat_goMux1_r  && (\call_main_map'_Bool_Nat_unlockFork1_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d [0]));
  assign \call_main_map'_Bool_Nat_unlockFork1_r  = (\call_main_map'_Bool_Nat_goMux1_r  && (\call_main_map'_Bool_Nat_unlockFork1_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natgo_7_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTNat_Bool) : (call_main_map'_Bool_Nat_unlockFork2,Go) [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ,MyDTNat_Bool)] > (call_main_map'_Bool_Nat_goMux2,MyDTNat_Bool) */
  assign \call_main_map'_Bool_Nat_goMux2_d  = (\call_main_map'_Bool_Nat_unlockFork2_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d [0]);
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_r  = (\call_main_map'_Bool_Nat_goMux2_r  && (\call_main_map'_Bool_Nat_unlockFork2_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d [0]));
  assign \call_main_map'_Bool_Nat_unlockFork2_r  = (\call_main_map'_Bool_Nat_goMux2_r  && (\call_main_map'_Bool_Nat_unlockFork2_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatisZacQ_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Nat) : (call_main_map'_Bool_Nat_unlockFork3,Go) [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR,MyDTBool_Nat)] > (call_main_map'_Bool_Nat_goMux3,MyDTBool_Nat) */
  assign \call_main_map'_Bool_Nat_goMux3_d  = (\call_main_map'_Bool_Nat_unlockFork3_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d [0]);
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_r  = (\call_main_map'_Bool_Nat_goMux3_r  && (\call_main_map'_Bool_Nat_unlockFork3_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d [0]));
  assign \call_main_map'_Bool_Nat_unlockFork3_r  = (\call_main_map'_Bool_Nat_goMux3_r  && (\call_main_map'_Bool_Nat_unlockFork3_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatgacR_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_main_map'_Bool_Nat_unlockFork4,Go) [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS,Pointer_QTree_Bool)] > (call_main_map'_Bool_Nat_goMux4,Pointer_QTree_Bool) */
  assign \call_main_map'_Bool_Nat_goMux4_d  = {\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d [16:1],
                                               (\call_main_map'_Bool_Nat_unlockFork4_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d [0])};
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_r  = (\call_main_map'_Bool_Nat_goMux4_r  && (\call_main_map'_Bool_Nat_unlockFork4_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d [0]));
  assign \call_main_map'_Bool_Nat_unlockFork4_r  = (\call_main_map'_Bool_Nat_goMux4_r  && (\call_main_map'_Bool_Nat_unlockFork4_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_NatmacS_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmain_map'_Bool_Nat) : (call_main_map'_Bool_Nat_unlockFork5,Go) [(call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1,Pointer_CTmain_map'_Bool_Nat)] > (call_main_map'_Bool_Nat_goMux5,Pointer_CTmain_map'_Bool_Nat) */
  assign \call_main_map'_Bool_Nat_goMux5_d  = {\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d [16:1],
                                               (\call_main_map'_Bool_Nat_unlockFork5_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d [0])};
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_r  = (\call_main_map'_Bool_Nat_goMux5_r  && (\call_main_map'_Bool_Nat_unlockFork5_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d [0]));
  assign \call_main_map'_Bool_Nat_unlockFork5_r  = (\call_main_map'_Bool_Nat_goMux5_r  && (\call_main_map'_Bool_Nat_unlockFork5_d [0] && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Natsc_0_1_d [0]));
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) : (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) > [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8,Go),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0,MyBool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                        (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [5:0] \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted ;
  logic [5:0] \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done ;
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [0]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [1]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [2]));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [1:1],
                                                                                                                                                                    (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [3]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [17:2],
                                                                                                                                                                   (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [4]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [33:18],
                                                                                                                                                                     (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0] && (! \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted [5]))};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done  = (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  | ({\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d [0],
                                                                                                                                                                                                                                                                                                                                   \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d [0]} & {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_r }));
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  = (& \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  <= 6'd0;
    else
      \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_emitted  <= (\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  ? 6'd0 :
                                                                                                                                                                     \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_done );
  
  /* rbuf (Ty Go) : (call_map''_map''_Bool_Bool_Bool_goConst,Go) > (call_map''_map''_Bool_Bool_Bool_initBufi,Go) */
  Go_t \call_map''_map''_Bool_Bool_Bool_goConst_buf ;
  assign \call_map''_map''_Bool_Bool_Bool_goConst_r  = (! \call_map''_map''_Bool_Bool_Bool_goConst_buf [0]);
  assign \call_map''_map''_Bool_Bool_Bool_initBufi_d  = (\call_map''_map''_Bool_Bool_Bool_goConst_buf [0] ? \call_map''_map''_Bool_Bool_Bool_goConst_buf  :
                                                         \call_map''_map''_Bool_Bool_Bool_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= 1'd0;
    else
      if ((\call_map''_map''_Bool_Bool_Bool_initBufi_r  && \call_map''_map''_Bool_Bool_Bool_goConst_buf [0]))
        \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= 1'd0;
      else if (((! \call_map''_map''_Bool_Bool_Bool_initBufi_r ) && (! \call_map''_map''_Bool_Bool_Bool_goConst_buf [0])))
        \call_map''_map''_Bool_Bool_Bool_goConst_buf  <= \call_map''_map''_Bool_Bool_Bool_goConst_d ;
  
  /* mergectrl (Ty C5,
           Ty Go) : [(call_map''_map''_Bool_Bool_Bool_goMux1,Go),
                     (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf,Go),
                     (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf,Go),
                     (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf,Go),
                     (lizzieLet12_1_4QNode_Bool_1_argbuf,Go)] > (go_8_goMux_choice,C5) (go_8_goMux_data,Go) */
  logic [4:0] \call_map''_map''_Bool_Bool_Bool_goMux1_select_d ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_select_d  = ((| \call_map''_map''_Bool_Bool_Bool_goMux1_select_q ) ? \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  :
                                                              (\call_map''_map''_Bool_Bool_Bool_goMux1_d [0] ? 5'd1 :
                                                               (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d [0] ? 5'd2 :
                                                                (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d [0] ? 5'd4 :
                                                                 (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d [0] ? 5'd8 :
                                                                  (lizzieLet12_1_4QNode_Bool_1_argbuf_d[0] ? 5'd16 :
                                                                   5'd0))))));
  logic [4:0] \call_map''_map''_Bool_Bool_Bool_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  <= 5'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_goMux1_select_q  <= (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? 5'd0 :
                                                            \call_map''_map''_Bool_Bool_Bool_goMux1_select_d );
  logic [1:0] \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  <= 2'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  <= (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? 2'd0 :
                                                          \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d );
  logic [1:0] \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d  = (\call_map''_map''_Bool_Bool_Bool_goMux1_emit_q  | ({go_8_goMux_choice_d[0],
                                                                                                                go_8_goMux_data_d[0]} & {go_8_goMux_choice_r,
                                                                                                                                         go_8_goMux_data_r}));
  logic \call_map''_map''_Bool_Bool_Bool_goMux1_done ;
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_done  = (& \call_map''_map''_Bool_Bool_Bool_goMux1_emit_d );
  assign {lizzieLet12_1_4QNode_Bool_1_argbuf_r,
          \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ,
          \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ,
          \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ,
          \call_map''_map''_Bool_Bool_Bool_goMux1_r } = (\call_map''_map''_Bool_Bool_Bool_goMux1_done  ? \call_map''_map''_Bool_Bool_Bool_goMux1_select_d  :
                                                         5'd0);
  assign go_8_goMux_data_d = ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [0] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \call_map''_map''_Bool_Bool_Bool_goMux1_d  :
                              ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [1] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d  :
                               ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [2] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d  :
                                ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [3] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d  :
                                 ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [4] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [0])) ? lizzieLet12_1_4QNode_Bool_1_argbuf_d :
                                  1'd0)))));
  assign go_8_goMux_choice_d = ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [0] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [1] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                 ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [2] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                  ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [3] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                   ((\call_map''_map''_Bool_Bool_Bool_goMux1_select_d [4] && (! \call_map''_map''_Bool_Bool_Bool_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                    {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_map''_map''_Bool_Bool_Bool_initBuf,Go) > [(call_map''_map''_Bool_Bool_Bool_unlockFork1,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork2,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork3,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork4,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork5,Go),
                                                               (call_map''_map''_Bool_Bool_Bool_unlockFork6,Go)] */
  logic [5:0] \call_map''_map''_Bool_Bool_Bool_initBuf_emitted ;
  logic [5:0] \call_map''_map''_Bool_Bool_Bool_initBuf_done ;
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork1_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork2_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [1]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork3_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [2]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork4_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [3]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork5_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [4]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork6_d  = (\call_map''_map''_Bool_Bool_Bool_initBuf_d [0] && (! \call_map''_map''_Bool_Bool_Bool_initBuf_emitted [5]));
  assign \call_map''_map''_Bool_Bool_Bool_initBuf_done  = (\call_map''_map''_Bool_Bool_Bool_initBuf_emitted  | ({\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0],
                                                                                                                 \call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0]} & {\call_map''_map''_Bool_Bool_Bool_unlockFork6_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork5_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork4_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork3_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork2_r ,
                                                                                                                                                                        \call_map''_map''_Bool_Bool_Bool_unlockFork1_r }));
  assign \call_map''_map''_Bool_Bool_Bool_initBuf_r  = (& \call_map''_map''_Bool_Bool_Bool_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_initBuf_emitted  <= 6'd0;
    else
      \call_map''_map''_Bool_Bool_Bool_initBuf_emitted  <= (\call_map''_map''_Bool_Bool_Bool_initBuf_r  ? 6'd0 :
                                                            \call_map''_map''_Bool_Bool_Bool_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_map''_map''_Bool_Bool_Bool_initBufi,Go) > (call_map''_map''_Bool_Bool_Bool_initBuf,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_initBufi_r  = ((! \call_map''_map''_Bool_Bool_Bool_initBuf_d [0]) || \call_map''_map''_Bool_Bool_Bool_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_map''_map''_Bool_Bool_Bool_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_map''_map''_Bool_Bool_Bool_initBufi_r )
        \call_map''_map''_Bool_Bool_Bool_initBuf_d  <= \call_map''_map''_Bool_Bool_Bool_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_map''_map''_Bool_Bool_Bool_unlockFork1,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8,Go)] > (call_map''_map''_Bool_Bool_Bool_goMux1,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux1_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_r  = (\call_map''_map''_Bool_Bool_Bool_goMux1_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork1_r  = (\call_map''_map''_Bool_Bool_Bool_goMux1_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork1_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolgo_8_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork2,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY,MyDTBool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux2,MyDTBool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux2_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_r  = (\call_map''_map''_Bool_Bool_Bool_goMux2_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork2_r  = (\call_map''_map''_Bool_Bool_Bool_goMux2_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork2_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolisZacY_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTBool_Bool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork3,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ,MyDTBool_Bool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux3_d  = (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d [0]);
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_r  = (\call_map''_map''_Bool_Bool_Bool_goMux3_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork3_r  = (\call_map''_map''_Bool_Bool_Bool_goMux3_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork3_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_BoolgacZ_d [0]));
  
  /* mux (Ty Go,
     Ty MyBool) : (call_map''_map''_Bool_Bool_Bool_unlockFork4,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0,MyBool)] > (call_map''_map''_Bool_Bool_Bool_goMux4,MyBool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux4_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d [1:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_r  = (\call_map''_map''_Bool_Bool_Bool_goMux4_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork4_r  = (\call_map''_map''_Bool_Bool_Bool_goMux4_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork4_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolv'ad0_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork5,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1,Pointer_QTree_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux5_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d [16:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_r  = (\call_map''_map''_Bool_Bool_Bool_goMux5_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork5_r  = (\call_map''_map''_Bool_Bool_Bool_goMux5_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork5_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolmad1_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (call_map''_map''_Bool_Bool_Bool_unlockFork6,Go) [(call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (call_map''_map''_Bool_Bool_Bool_goMux6,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_Bool_goMux6_d  = {\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [16:1],
                                                       (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0])};
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_r  = (\call_map''_map''_Bool_Bool_Bool_goMux6_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0]));
  assign \call_map''_map''_Bool_Bool_Bool_unlockFork6_r  = (\call_map''_map''_Bool_Bool_Bool_goMux6_r  && (\call_map''_map''_Bool_Bool_Bool_unlockFork6_d [0] && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Boolsc_0_2_d [0]));
  
  /* destruct (Ty TupGo___Pointer_Nat___Pointer_Nat,
          Dcon TupGo___Pointer_Nat___Pointer_Nat) : (eqNatTupGo___Pointer_Nat___Pointer_Nat_1,TupGo___Pointer_Nat___Pointer_Nat) > [(eqNatTupGo___Pointer_Nat___Pointer_Natgo_9,Go),
                                                                                                                                    (eqNatTupGo___Pointer_Nat___Pointer_Natxadg,Pointer_Nat),
                                                                                                                                    (eqNatTupGo___Pointer_Nat___Pointer_Natyadh,Pointer_Nat)] */
  logic [2:0] eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted;
  logic [2:0] eqNatTupGo___Pointer_Nat___Pointer_Nat_1_done;
  assign eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d = (eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[0] && (! eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted[0]));
  assign eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d = {eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[16:1],
                                                         (eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[0] && (! eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted[1]))};
  assign eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d = {eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[32:17],
                                                         (eqNatTupGo___Pointer_Nat___Pointer_Nat_1_d[0] && (! eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted[2]))};
  assign eqNatTupGo___Pointer_Nat___Pointer_Nat_1_done = (eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted | ({eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d[0],
                                                                                                               eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d[0],
                                                                                                               eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d[0]} & {eqNatTupGo___Pointer_Nat___Pointer_Natyadh_r,
                                                                                                                                                                   eqNatTupGo___Pointer_Nat___Pointer_Natxadg_r,
                                                                                                                                                                   eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_r}));
  assign eqNatTupGo___Pointer_Nat___Pointer_Nat_1_r = (& eqNatTupGo___Pointer_Nat___Pointer_Nat_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted <= 3'd0;
    else
      eqNatTupGo___Pointer_Nat___Pointer_Nat_1_emitted <= (eqNatTupGo___Pointer_Nat___Pointer_Nat_1_r ? 3'd0 :
                                                           eqNatTupGo___Pointer_Nat___Pointer_Nat_1_done);
  
  /* buf (Ty MyBool) : (eqNat_1_mux,MyBool) > (applyfnNat_Bool_5_resbuf,MyBool) */
  MyBool_t eqNat_1_mux_bufchan_d;
  logic eqNat_1_mux_bufchan_r;
  assign eqNat_1_mux_r = ((! eqNat_1_mux_bufchan_d[0]) || eqNat_1_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_1_mux_bufchan_d <= {1'd0, 1'd0};
    else if (eqNat_1_mux_r) eqNat_1_mux_bufchan_d <= eqNat_1_mux_d;
  MyBool_t eqNat_1_mux_bufchan_buf;
  assign eqNat_1_mux_bufchan_r = (! eqNat_1_mux_bufchan_buf[0]);
  assign applyfnNat_Bool_5_resbuf_d = (eqNat_1_mux_bufchan_buf[0] ? eqNat_1_mux_bufchan_buf :
                                       eqNat_1_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_1_mux_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnNat_Bool_5_resbuf_r && eqNat_1_mux_bufchan_buf[0]))
        eqNat_1_mux_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnNat_Bool_5_resbuf_r) && (! eqNat_1_mux_bufchan_buf[0])))
        eqNat_1_mux_bufchan_buf <= eqNat_1_mux_bufchan_d;
  
  /* rbuf (Ty Go) : (eqNat_goConst,Go) > (eqNat_initBufi,Go) */
  Go_t eqNat_goConst_buf;
  assign eqNat_goConst_r = (! eqNat_goConst_buf[0]);
  assign eqNat_initBufi_d = (eqNat_goConst_buf[0] ? eqNat_goConst_buf :
                             eqNat_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_goConst_buf <= 1'd0;
    else
      if ((eqNat_initBufi_r && eqNat_goConst_buf[0]))
        eqNat_goConst_buf <= 1'd0;
      else if (((! eqNat_initBufi_r) && (! eqNat_goConst_buf[0])))
        eqNat_goConst_buf <= eqNat_goConst_d;
  
  /* mergectrl (Ty C2,Ty Go) : [(eqNat_goMux1,Go),
                           (lizzieLet18_4Succ_3Succ_1_argbuf,Go)] > (go_9_goMux_choice,C2) (go_9_goMux_data,Go) */
  logic [1:0] eqNat_goMux1_select_d;
  assign eqNat_goMux1_select_d = ((| eqNat_goMux1_select_q) ? eqNat_goMux1_select_q :
                                  (eqNat_goMux1_d[0] ? 2'd1 :
                                   (lizzieLet18_4Succ_3Succ_1_argbuf_d[0] ? 2'd2 :
                                    2'd0)));
  logic [1:0] eqNat_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_goMux1_select_q <= 2'd0;
    else
      eqNat_goMux1_select_q <= (eqNat_goMux1_done ? 2'd0 :
                                eqNat_goMux1_select_d);
  logic [1:0] eqNat_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_goMux1_emit_q <= 2'd0;
    else
      eqNat_goMux1_emit_q <= (eqNat_goMux1_done ? 2'd0 :
                              eqNat_goMux1_emit_d);
  logic [1:0] eqNat_goMux1_emit_d;
  assign eqNat_goMux1_emit_d = (eqNat_goMux1_emit_q | ({go_9_goMux_choice_d[0],
                                                        go_9_goMux_data_d[0]} & {go_9_goMux_choice_r,
                                                                                 go_9_goMux_data_r}));
  logic eqNat_goMux1_done;
  assign eqNat_goMux1_done = (& eqNat_goMux1_emit_d);
  assign {lizzieLet18_4Succ_3Succ_1_argbuf_r,
          eqNat_goMux1_r} = (eqNat_goMux1_done ? eqNat_goMux1_select_d :
                             2'd0);
  assign go_9_goMux_data_d = ((eqNat_goMux1_select_d[0] && (! eqNat_goMux1_emit_q[0])) ? eqNat_goMux1_d :
                              ((eqNat_goMux1_select_d[1] && (! eqNat_goMux1_emit_q[0])) ? lizzieLet18_4Succ_3Succ_1_argbuf_d :
                               1'd0));
  assign go_9_goMux_choice_d = ((eqNat_goMux1_select_d[0] && (! eqNat_goMux1_emit_q[1])) ? C1_2_dc(1'd1) :
                                ((eqNat_goMux1_select_d[1] && (! eqNat_goMux1_emit_q[1])) ? C2_2_dc(1'd1) :
                                 {1'd0, 1'd0}));
  
  /* fork (Ty Go) : (eqNat_initBuf,Go) > [(eqNat_unlockFork1,Go),
                                     (eqNat_unlockFork2,Go),
                                     (eqNat_unlockFork3,Go)] */
  logic [2:0] eqNat_initBuf_emitted;
  logic [2:0] eqNat_initBuf_done;
  assign eqNat_unlockFork1_d = (eqNat_initBuf_d[0] && (! eqNat_initBuf_emitted[0]));
  assign eqNat_unlockFork2_d = (eqNat_initBuf_d[0] && (! eqNat_initBuf_emitted[1]));
  assign eqNat_unlockFork3_d = (eqNat_initBuf_d[0] && (! eqNat_initBuf_emitted[2]));
  assign eqNat_initBuf_done = (eqNat_initBuf_emitted | ({eqNat_unlockFork3_d[0],
                                                         eqNat_unlockFork2_d[0],
                                                         eqNat_unlockFork1_d[0]} & {eqNat_unlockFork3_r,
                                                                                    eqNat_unlockFork2_r,
                                                                                    eqNat_unlockFork1_r}));
  assign eqNat_initBuf_r = (& eqNat_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_initBuf_emitted <= 3'd0;
    else
      eqNat_initBuf_emitted <= (eqNat_initBuf_r ? 3'd0 :
                                eqNat_initBuf_done);
  
  /* initbuf (Ty Go,Dcon Go) : (eqNat_initBufi,Go) > (eqNat_initBuf,Go) */
  assign eqNat_initBufi_r = ((! eqNat_initBuf_d[0]) || eqNat_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) eqNat_initBuf_d <= Go_dc(1'd1);
    else if (eqNat_initBufi_r) eqNat_initBuf_d <= eqNat_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (eqNat_unlockFork1,Go) [(eqNatTupGo___Pointer_Nat___Pointer_Natgo_9,Go)] > (eqNat_goMux1,Go) */
  assign eqNat_goMux1_d = (eqNat_unlockFork1_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d[0]);
  assign eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_r = (eqNat_goMux1_r && (eqNat_unlockFork1_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d[0]));
  assign eqNat_unlockFork1_r = (eqNat_goMux1_r && (eqNat_unlockFork1_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natgo_9_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_Nat) : (eqNat_unlockFork2,Go) [(eqNatTupGo___Pointer_Nat___Pointer_Natxadg,Pointer_Nat)] > (eqNat_goMux2,Pointer_Nat) */
  assign eqNat_goMux2_d = {eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d[16:1],
                           (eqNat_unlockFork2_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d[0])};
  assign eqNatTupGo___Pointer_Nat___Pointer_Natxadg_r = (eqNat_goMux2_r && (eqNat_unlockFork2_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d[0]));
  assign eqNat_unlockFork2_r = (eqNat_goMux2_r && (eqNat_unlockFork2_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natxadg_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_Nat) : (eqNat_unlockFork3,Go) [(eqNatTupGo___Pointer_Nat___Pointer_Natyadh,Pointer_Nat)] > (eqNat_goMux3,Pointer_Nat) */
  assign eqNat_goMux3_d = {eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d[16:1],
                           (eqNat_unlockFork3_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d[0])};
  assign eqNatTupGo___Pointer_Nat___Pointer_Natyadh_r = (eqNat_goMux3_r && (eqNat_unlockFork3_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d[0]));
  assign eqNat_unlockFork3_r = (eqNat_goMux3_r && (eqNat_unlockFork3_d[0] && eqNatTupGo___Pointer_Nat___Pointer_Natyadh_d[0]));
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_1_1,MyBool) (lizzieLet6_4QVal_Bool_3,Go) > [(es_0_1_1MyFalse,Go),
                                                                  (es_0_1_1MyTrue,Go)] */
  logic [1:0] lizzieLet6_4QVal_Bool_3_onehotd;
  always_comb
    if ((es_0_1_1_d[0] && lizzieLet6_4QVal_Bool_3_d[0]))
      unique case (es_0_1_1_d[1:1])
        1'd0: lizzieLet6_4QVal_Bool_3_onehotd = 2'd1;
        1'd1: lizzieLet6_4QVal_Bool_3_onehotd = 2'd2;
        default: lizzieLet6_4QVal_Bool_3_onehotd = 2'd0;
      endcase
    else lizzieLet6_4QVal_Bool_3_onehotd = 2'd0;
  assign es_0_1_1MyFalse_d = lizzieLet6_4QVal_Bool_3_onehotd[0];
  assign es_0_1_1MyTrue_d = lizzieLet6_4QVal_Bool_3_onehotd[1];
  assign lizzieLet6_4QVal_Bool_3_r = (| (lizzieLet6_4QVal_Bool_3_onehotd & {es_0_1_1MyTrue_r,
                                                                            es_0_1_1MyFalse_r}));
  assign es_0_1_1_r = lizzieLet6_4QVal_Bool_3_r;
  
  /* buf (Ty Go) : (es_0_1_1MyFalse,Go) > (es_0_1_1MyFalse_1_argbuf,Go) */
  Go_t es_0_1_1MyFalse_bufchan_d;
  logic es_0_1_1MyFalse_bufchan_r;
  assign es_0_1_1MyFalse_r = ((! es_0_1_1MyFalse_bufchan_d[0]) || es_0_1_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_1_1MyFalse_r)
        es_0_1_1MyFalse_bufchan_d <= es_0_1_1MyFalse_d;
  Go_t es_0_1_1MyFalse_bufchan_buf;
  assign es_0_1_1MyFalse_bufchan_r = (! es_0_1_1MyFalse_bufchan_buf[0]);
  assign es_0_1_1MyFalse_1_argbuf_d = (es_0_1_1MyFalse_bufchan_buf[0] ? es_0_1_1MyFalse_bufchan_buf :
                                       es_0_1_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_1_1MyFalse_1_argbuf_r && es_0_1_1MyFalse_bufchan_buf[0]))
        es_0_1_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_1_1MyFalse_1_argbuf_r) && (! es_0_1_1MyFalse_bufchan_buf[0])))
        es_0_1_1MyFalse_bufchan_buf <= es_0_1_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_1_1MyTrue,Go) > [(es_0_1_1MyTrue_1,Go),
                                      (es_0_1_1MyTrue_2,Go)] */
  logic [1:0] es_0_1_1MyTrue_emitted;
  logic [1:0] es_0_1_1MyTrue_done;
  assign es_0_1_1MyTrue_1_d = (es_0_1_1MyTrue_d[0] && (! es_0_1_1MyTrue_emitted[0]));
  assign es_0_1_1MyTrue_2_d = (es_0_1_1MyTrue_d[0] && (! es_0_1_1MyTrue_emitted[1]));
  assign es_0_1_1MyTrue_done = (es_0_1_1MyTrue_emitted | ({es_0_1_1MyTrue_2_d[0],
                                                           es_0_1_1MyTrue_1_d[0]} & {es_0_1_1MyTrue_2_r,
                                                                                     es_0_1_1MyTrue_1_r}));
  assign es_0_1_1MyTrue_r = (& es_0_1_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_emitted <= 2'd0;
    else
      es_0_1_1MyTrue_emitted <= (es_0_1_1MyTrue_r ? 2'd0 :
                                 es_0_1_1MyTrue_done);
  
  /* dcon (Ty QTree_Nat,
      Dcon QNone_Nat) : [(es_0_1_1MyTrue_1,Go)] > (es_0_1_1MyTrue_1QNone_Nat,QTree_Nat) */
  assign es_0_1_1MyTrue_1QNone_Nat_d = QNone_Nat_dc((& {es_0_1_1MyTrue_1_d[0]}), es_0_1_1MyTrue_1_d);
  assign {es_0_1_1MyTrue_1_r} = {1 {(es_0_1_1MyTrue_1QNone_Nat_r && es_0_1_1MyTrue_1QNone_Nat_d[0])}};
  
  /* buf (Ty QTree_Nat) : (es_0_1_1MyTrue_1QNone_Nat,QTree_Nat) > (lizzieLet9_1_argbuf,QTree_Nat) */
  QTree_Nat_t es_0_1_1MyTrue_1QNone_Nat_bufchan_d;
  logic es_0_1_1MyTrue_1QNone_Nat_bufchan_r;
  assign es_0_1_1MyTrue_1QNone_Nat_r = ((! es_0_1_1MyTrue_1QNone_Nat_bufchan_d[0]) || es_0_1_1MyTrue_1QNone_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1MyTrue_1QNone_Nat_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_1MyTrue_1QNone_Nat_r)
        es_0_1_1MyTrue_1QNone_Nat_bufchan_d <= es_0_1_1MyTrue_1QNone_Nat_d;
  QTree_Nat_t es_0_1_1MyTrue_1QNone_Nat_bufchan_buf;
  assign es_0_1_1MyTrue_1QNone_Nat_bufchan_r = (! es_0_1_1MyTrue_1QNone_Nat_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (es_0_1_1MyTrue_1QNone_Nat_bufchan_buf[0] ? es_0_1_1MyTrue_1QNone_Nat_bufchan_buf :
                                  es_0_1_1MyTrue_1QNone_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_1MyTrue_1QNone_Nat_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && es_0_1_1MyTrue_1QNone_Nat_bufchan_buf[0]))
        es_0_1_1MyTrue_1QNone_Nat_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! es_0_1_1MyTrue_1QNone_Nat_bufchan_buf[0])))
        es_0_1_1MyTrue_1QNone_Nat_bufchan_buf <= es_0_1_1MyTrue_1QNone_Nat_bufchan_d;
  
  /* buf (Ty Go) : (es_0_1_1MyTrue_2,Go) > (es_0_1_1MyTrue_2_argbuf,Go) */
  Go_t es_0_1_1MyTrue_2_bufchan_d;
  logic es_0_1_1MyTrue_2_bufchan_r;
  assign es_0_1_1MyTrue_2_r = ((! es_0_1_1MyTrue_2_bufchan_d[0]) || es_0_1_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_1_1MyTrue_2_r)
        es_0_1_1MyTrue_2_bufchan_d <= es_0_1_1MyTrue_2_d;
  Go_t es_0_1_1MyTrue_2_bufchan_buf;
  assign es_0_1_1MyTrue_2_bufchan_r = (! es_0_1_1MyTrue_2_bufchan_buf[0]);
  assign es_0_1_1MyTrue_2_argbuf_d = (es_0_1_1MyTrue_2_bufchan_buf[0] ? es_0_1_1MyTrue_2_bufchan_buf :
                                      es_0_1_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_1_1MyTrue_2_argbuf_r && es_0_1_1MyTrue_2_bufchan_buf[0]))
        es_0_1_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_1_1MyTrue_2_argbuf_r) && (! es_0_1_1MyTrue_2_bufchan_buf[0])))
        es_0_1_1MyTrue_2_bufchan_buf <= es_0_1_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmain_map'_Bool_Nat) : (es_0_1_2,MyBool) (lizzieLet6_6QVal_Bool,Pointer_CTmain_map'_Bool_Nat) > [(es_0_1_2MyFalse,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                    (es_0_1_2MyTrue,Pointer_CTmain_map'_Bool_Nat)] */
  logic [1:0] lizzieLet6_6QVal_Bool_onehotd;
  always_comb
    if ((es_0_1_2_d[0] && lizzieLet6_6QVal_Bool_d[0]))
      unique case (es_0_1_2_d[1:1])
        1'd0: lizzieLet6_6QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet6_6QVal_Bool_onehotd = 2'd2;
        default: lizzieLet6_6QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet6_6QVal_Bool_onehotd = 2'd0;
  assign es_0_1_2MyFalse_d = {lizzieLet6_6QVal_Bool_d[16:1],
                              lizzieLet6_6QVal_Bool_onehotd[0]};
  assign es_0_1_2MyTrue_d = {lizzieLet6_6QVal_Bool_d[16:1],
                             lizzieLet6_6QVal_Bool_onehotd[1]};
  assign lizzieLet6_6QVal_Bool_r = (| (lizzieLet6_6QVal_Bool_onehotd & {es_0_1_2MyTrue_r,
                                                                        es_0_1_2MyFalse_r}));
  assign es_0_1_2_r = lizzieLet6_6QVal_Bool_r;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (es_0_1_2MyFalse,Pointer_CTmain_map'_Bool_Nat) > (es_0_1_2MyFalse_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyFalse_bufchan_d;
  logic es_0_1_2MyFalse_bufchan_r;
  assign es_0_1_2MyFalse_r = ((! es_0_1_2MyFalse_bufchan_d[0]) || es_0_1_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_1_2MyFalse_r)
        es_0_1_2MyFalse_bufchan_d <= es_0_1_2MyFalse_d;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyFalse_bufchan_buf;
  assign es_0_1_2MyFalse_bufchan_r = (! es_0_1_2MyFalse_bufchan_buf[0]);
  assign es_0_1_2MyFalse_1_argbuf_d = (es_0_1_2MyFalse_bufchan_buf[0] ? es_0_1_2MyFalse_bufchan_buf :
                                       es_0_1_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_2MyFalse_1_argbuf_r && es_0_1_2MyFalse_bufchan_buf[0]))
        es_0_1_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_2MyFalse_1_argbuf_r) && (! es_0_1_2MyFalse_bufchan_buf[0])))
        es_0_1_2MyFalse_bufchan_buf <= es_0_1_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (es_0_1_2MyTrue,Pointer_CTmain_map'_Bool_Nat) > (es_0_1_2MyTrue_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyTrue_bufchan_d;
  logic es_0_1_2MyTrue_bufchan_r;
  assign es_0_1_2MyTrue_r = ((! es_0_1_2MyTrue_bufchan_d[0]) || es_0_1_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_1_2MyTrue_r) es_0_1_2MyTrue_bufchan_d <= es_0_1_2MyTrue_d;
  \Pointer_CTmain_map'_Bool_Nat_t  es_0_1_2MyTrue_bufchan_buf;
  assign es_0_1_2MyTrue_bufchan_r = (! es_0_1_2MyTrue_bufchan_buf[0]);
  assign es_0_1_2MyTrue_1_argbuf_d = (es_0_1_2MyTrue_bufchan_buf[0] ? es_0_1_2MyTrue_bufchan_buf :
                                      es_0_1_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_2MyTrue_1_argbuf_r && es_0_1_2MyTrue_bufchan_buf[0]))
        es_0_1_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_2MyTrue_1_argbuf_r) && (! es_0_1_2MyTrue_bufchan_buf[0])))
        es_0_1_2MyTrue_bufchan_buf <= es_0_1_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_Nat) : (es_0_1_3,MyBool) (xacw_2,Pointer_Nat) > [(es_0_1_3MyFalse,Pointer_Nat),
                                                                   (_32,Pointer_Nat)] */
  logic [1:0] xacw_2_onehotd;
  always_comb
    if ((es_0_1_3_d[0] && xacw_2_d[0]))
      unique case (es_0_1_3_d[1:1])
        1'd0: xacw_2_onehotd = 2'd1;
        1'd1: xacw_2_onehotd = 2'd2;
        default: xacw_2_onehotd = 2'd0;
      endcase
    else xacw_2_onehotd = 2'd0;
  assign es_0_1_3MyFalse_d = {xacw_2_d[16:1], xacw_2_onehotd[0]};
  assign _32_d = {xacw_2_d[16:1], xacw_2_onehotd[1]};
  assign xacw_2_r = (| (xacw_2_onehotd & {_32_r,
                                          es_0_1_3MyFalse_r}));
  assign es_0_1_3_r = xacw_2_r;
  
  /* dcon (Ty QTree_Nat,
      Dcon QVal_Nat) : [(es_0_1_3MyFalse,Pointer_Nat)] > (es_0_1_3MyFalse_1QVal_Nat,QTree_Nat) */
  assign es_0_1_3MyFalse_1QVal_Nat_d = QVal_Nat_dc((& {es_0_1_3MyFalse_d[0]}), es_0_1_3MyFalse_d);
  assign {es_0_1_3MyFalse_r} = {1 {(es_0_1_3MyFalse_1QVal_Nat_r && es_0_1_3MyFalse_1QVal_Nat_d[0])}};
  
  /* buf (Ty QTree_Nat) : (es_0_1_3MyFalse_1QVal_Nat,QTree_Nat) > (lizzieLet8_1_argbuf,QTree_Nat) */
  QTree_Nat_t es_0_1_3MyFalse_1QVal_Nat_bufchan_d;
  logic es_0_1_3MyFalse_1QVal_Nat_bufchan_r;
  assign es_0_1_3MyFalse_1QVal_Nat_r = ((! es_0_1_3MyFalse_1QVal_Nat_bufchan_d[0]) || es_0_1_3MyFalse_1QVal_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_3MyFalse_1QVal_Nat_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_1_3MyFalse_1QVal_Nat_r)
        es_0_1_3MyFalse_1QVal_Nat_bufchan_d <= es_0_1_3MyFalse_1QVal_Nat_d;
  QTree_Nat_t es_0_1_3MyFalse_1QVal_Nat_bufchan_buf;
  assign es_0_1_3MyFalse_1QVal_Nat_bufchan_r = (! es_0_1_3MyFalse_1QVal_Nat_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (es_0_1_3MyFalse_1QVal_Nat_bufchan_buf[0] ? es_0_1_3MyFalse_1QVal_Nat_bufchan_buf :
                                  es_0_1_3MyFalse_1QVal_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_1_3MyFalse_1QVal_Nat_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && es_0_1_3MyFalse_1QVal_Nat_bufchan_buf[0]))
        es_0_1_3MyFalse_1QVal_Nat_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! es_0_1_3MyFalse_1QVal_Nat_bufchan_buf[0])))
        es_0_1_3MyFalse_1QVal_Nat_bufchan_buf <= es_0_1_3MyFalse_1QVal_Nat_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_0_2_1,MyBool) (lizzieLet12_1_4QVal_Bool_3,Go) > [(es_0_2_1MyFalse,Go),
                                                                     (es_0_2_1MyTrue,Go)] */
  logic [1:0] lizzieLet12_1_4QVal_Bool_3_onehotd;
  always_comb
    if ((es_0_2_1_d[0] && lizzieLet12_1_4QVal_Bool_3_d[0]))
      unique case (es_0_2_1_d[1:1])
        1'd0: lizzieLet12_1_4QVal_Bool_3_onehotd = 2'd1;
        1'd1: lizzieLet12_1_4QVal_Bool_3_onehotd = 2'd2;
        default: lizzieLet12_1_4QVal_Bool_3_onehotd = 2'd0;
      endcase
    else lizzieLet12_1_4QVal_Bool_3_onehotd = 2'd0;
  assign es_0_2_1MyFalse_d = lizzieLet12_1_4QVal_Bool_3_onehotd[0];
  assign es_0_2_1MyTrue_d = lizzieLet12_1_4QVal_Bool_3_onehotd[1];
  assign lizzieLet12_1_4QVal_Bool_3_r = (| (lizzieLet12_1_4QVal_Bool_3_onehotd & {es_0_2_1MyTrue_r,
                                                                                  es_0_2_1MyFalse_r}));
  assign es_0_2_1_r = lizzieLet12_1_4QVal_Bool_3_r;
  
  /* buf (Ty Go) : (es_0_2_1MyFalse,Go) > (es_0_2_1MyFalse_1_argbuf,Go) */
  Go_t es_0_2_1MyFalse_bufchan_d;
  logic es_0_2_1MyFalse_bufchan_r;
  assign es_0_2_1MyFalse_r = ((! es_0_2_1MyFalse_bufchan_d[0]) || es_0_2_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_0_2_1MyFalse_r)
        es_0_2_1MyFalse_bufchan_d <= es_0_2_1MyFalse_d;
  Go_t es_0_2_1MyFalse_bufchan_buf;
  assign es_0_2_1MyFalse_bufchan_r = (! es_0_2_1MyFalse_bufchan_buf[0]);
  assign es_0_2_1MyFalse_1_argbuf_d = (es_0_2_1MyFalse_bufchan_buf[0] ? es_0_2_1MyFalse_bufchan_buf :
                                       es_0_2_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_0_2_1MyFalse_1_argbuf_r && es_0_2_1MyFalse_bufchan_buf[0]))
        es_0_2_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_0_2_1MyFalse_1_argbuf_r) && (! es_0_2_1MyFalse_bufchan_buf[0])))
        es_0_2_1MyFalse_bufchan_buf <= es_0_2_1MyFalse_bufchan_d;
  
  /* fork (Ty Go) : (es_0_2_1MyTrue,Go) > [(es_0_2_1MyTrue_1,Go),
                                      (es_0_2_1MyTrue_2,Go)] */
  logic [1:0] es_0_2_1MyTrue_emitted;
  logic [1:0] es_0_2_1MyTrue_done;
  assign es_0_2_1MyTrue_1_d = (es_0_2_1MyTrue_d[0] && (! es_0_2_1MyTrue_emitted[0]));
  assign es_0_2_1MyTrue_2_d = (es_0_2_1MyTrue_d[0] && (! es_0_2_1MyTrue_emitted[1]));
  assign es_0_2_1MyTrue_done = (es_0_2_1MyTrue_emitted | ({es_0_2_1MyTrue_2_d[0],
                                                           es_0_2_1MyTrue_1_d[0]} & {es_0_2_1MyTrue_2_r,
                                                                                     es_0_2_1MyTrue_1_r}));
  assign es_0_2_1MyTrue_r = (& es_0_2_1MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_emitted <= 2'd0;
    else
      es_0_2_1MyTrue_emitted <= (es_0_2_1MyTrue_r ? 2'd0 :
                                 es_0_2_1MyTrue_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(es_0_2_1MyTrue_1,Go)] > (es_0_2_1MyTrue_1QNone_Bool,QTree_Bool) */
  assign es_0_2_1MyTrue_1QNone_Bool_d = QNone_Bool_dc((& {es_0_2_1MyTrue_1_d[0]}), es_0_2_1MyTrue_1_d);
  assign {es_0_2_1MyTrue_1_r} = {1 {(es_0_2_1MyTrue_1QNone_Bool_r && es_0_2_1MyTrue_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_2_1MyTrue_1QNone_Bool,QTree_Bool) > (lizzieLet15_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_2_1MyTrue_1QNone_Bool_bufchan_d;
  logic es_0_2_1MyTrue_1QNone_Bool_bufchan_r;
  assign es_0_2_1MyTrue_1QNone_Bool_r = ((! es_0_2_1MyTrue_1QNone_Bool_bufchan_d[0]) || es_0_2_1MyTrue_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1MyTrue_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_2_1MyTrue_1QNone_Bool_r)
        es_0_2_1MyTrue_1QNone_Bool_bufchan_d <= es_0_2_1MyTrue_1QNone_Bool_d;
  QTree_Bool_t es_0_2_1MyTrue_1QNone_Bool_bufchan_buf;
  assign es_0_2_1MyTrue_1QNone_Bool_bufchan_r = (! es_0_2_1MyTrue_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (es_0_2_1MyTrue_1QNone_Bool_bufchan_buf[0] ? es_0_2_1MyTrue_1QNone_Bool_bufchan_buf :
                                   es_0_2_1MyTrue_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && es_0_2_1MyTrue_1QNone_Bool_bufchan_buf[0]))
        es_0_2_1MyTrue_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! es_0_2_1MyTrue_1QNone_Bool_bufchan_buf[0])))
        es_0_2_1MyTrue_1QNone_Bool_bufchan_buf <= es_0_2_1MyTrue_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (es_0_2_1MyTrue_2,Go) > (es_0_2_1MyTrue_2_argbuf,Go) */
  Go_t es_0_2_1MyTrue_2_bufchan_d;
  logic es_0_2_1MyTrue_2_bufchan_r;
  assign es_0_2_1MyTrue_2_r = ((! es_0_2_1MyTrue_2_bufchan_d[0]) || es_0_2_1MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_0_2_1MyTrue_2_r)
        es_0_2_1MyTrue_2_bufchan_d <= es_0_2_1MyTrue_2_d;
  Go_t es_0_2_1MyTrue_2_bufchan_buf;
  assign es_0_2_1MyTrue_2_bufchan_r = (! es_0_2_1MyTrue_2_bufchan_buf[0]);
  assign es_0_2_1MyTrue_2_argbuf_d = (es_0_2_1MyTrue_2_bufchan_buf[0] ? es_0_2_1MyTrue_2_bufchan_buf :
                                      es_0_2_1MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_1MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_0_2_1MyTrue_2_argbuf_r && es_0_2_1MyTrue_2_bufchan_buf[0]))
        es_0_2_1MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_0_2_1MyTrue_2_argbuf_r) && (! es_0_2_1MyTrue_2_bufchan_buf[0])))
        es_0_2_1MyTrue_2_bufchan_buf <= es_0_2_1MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_2_2,MyBool) (lizzieLet12_1_6QVal_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(es_0_2_2MyFalse,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (es_0_2_2MyTrue,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [1:0] lizzieLet12_1_6QVal_Bool_onehotd;
  always_comb
    if ((es_0_2_2_d[0] && lizzieLet12_1_6QVal_Bool_d[0]))
      unique case (es_0_2_2_d[1:1])
        1'd0: lizzieLet12_1_6QVal_Bool_onehotd = 2'd1;
        1'd1: lizzieLet12_1_6QVal_Bool_onehotd = 2'd2;
        default: lizzieLet12_1_6QVal_Bool_onehotd = 2'd0;
      endcase
    else lizzieLet12_1_6QVal_Bool_onehotd = 2'd0;
  assign es_0_2_2MyFalse_d = {lizzieLet12_1_6QVal_Bool_d[16:1],
                              lizzieLet12_1_6QVal_Bool_onehotd[0]};
  assign es_0_2_2MyTrue_d = {lizzieLet12_1_6QVal_Bool_d[16:1],
                             lizzieLet12_1_6QVal_Bool_onehotd[1]};
  assign lizzieLet12_1_6QVal_Bool_r = (| (lizzieLet12_1_6QVal_Bool_onehotd & {es_0_2_2MyTrue_r,
                                                                              es_0_2_2MyFalse_r}));
  assign es_0_2_2_r = lizzieLet12_1_6QVal_Bool_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_2_2MyFalse,Pointer_CTmap''_map''_Bool_Bool_Bool) > (es_0_2_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyFalse_bufchan_d;
  logic es_0_2_2MyFalse_bufchan_r;
  assign es_0_2_2MyFalse_r = ((! es_0_2_2MyFalse_bufchan_d[0]) || es_0_2_2MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_2_2MyFalse_r)
        es_0_2_2MyFalse_bufchan_d <= es_0_2_2MyFalse_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyFalse_bufchan_buf;
  assign es_0_2_2MyFalse_bufchan_r = (! es_0_2_2MyFalse_bufchan_buf[0]);
  assign es_0_2_2MyFalse_1_argbuf_d = (es_0_2_2MyFalse_bufchan_buf[0] ? es_0_2_2MyFalse_bufchan_buf :
                                       es_0_2_2MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_2_2MyFalse_1_argbuf_r && es_0_2_2MyFalse_bufchan_buf[0]))
        es_0_2_2MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_2_2MyFalse_1_argbuf_r) && (! es_0_2_2MyFalse_bufchan_buf[0])))
        es_0_2_2MyFalse_bufchan_buf <= es_0_2_2MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (es_0_2_2MyTrue,Pointer_CTmap''_map''_Bool_Bool_Bool) > (es_0_2_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyTrue_bufchan_d;
  logic es_0_2_2MyTrue_bufchan_r;
  assign es_0_2_2MyTrue_r = ((! es_0_2_2MyTrue_bufchan_d[0]) || es_0_2_2MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_0_2_2MyTrue_r) es_0_2_2MyTrue_bufchan_d <= es_0_2_2MyTrue_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  es_0_2_2MyTrue_bufchan_buf;
  assign es_0_2_2MyTrue_bufchan_r = (! es_0_2_2MyTrue_bufchan_buf[0]);
  assign es_0_2_2MyTrue_1_argbuf_d = (es_0_2_2MyTrue_bufchan_buf[0] ? es_0_2_2MyTrue_bufchan_buf :
                                      es_0_2_2MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_0_2_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_2_2MyTrue_1_argbuf_r && es_0_2_2MyTrue_bufchan_buf[0]))
        es_0_2_2MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_2_2MyTrue_1_argbuf_r) && (! es_0_2_2MyTrue_bufchan_buf[0])))
        es_0_2_2MyTrue_bufchan_buf <= es_0_2_2MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyBool) : (es_0_2_3,MyBool) (xacw_1_2,MyBool) > [(es_0_2_3MyFalse,MyBool),
                                                           (_31,MyBool)] */
  logic [1:0] xacw_1_2_onehotd;
  always_comb
    if ((es_0_2_3_d[0] && xacw_1_2_d[0]))
      unique case (es_0_2_3_d[1:1])
        1'd0: xacw_1_2_onehotd = 2'd1;
        1'd1: xacw_1_2_onehotd = 2'd2;
        default: xacw_1_2_onehotd = 2'd0;
      endcase
    else xacw_1_2_onehotd = 2'd0;
  assign es_0_2_3MyFalse_d = {xacw_1_2_d[1:1], xacw_1_2_onehotd[0]};
  assign _31_d = {xacw_1_2_d[1:1], xacw_1_2_onehotd[1]};
  assign xacw_1_2_r = (| (xacw_1_2_onehotd & {_31_r,
                                              es_0_2_3MyFalse_r}));
  assign es_0_2_3_r = xacw_1_2_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QVal_Bool) : [(es_0_2_3MyFalse,MyBool)] > (es_0_2_3MyFalse_1QVal_Bool,QTree_Bool) */
  assign es_0_2_3MyFalse_1QVal_Bool_d = QVal_Bool_dc((& {es_0_2_3MyFalse_d[0]}), es_0_2_3MyFalse_d);
  assign {es_0_2_3MyFalse_r} = {1 {(es_0_2_3MyFalse_1QVal_Bool_r && es_0_2_3MyFalse_1QVal_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (es_0_2_3MyFalse_1QVal_Bool,QTree_Bool) > (lizzieLet14_1_argbuf,QTree_Bool) */
  QTree_Bool_t es_0_2_3MyFalse_1QVal_Bool_bufchan_d;
  logic es_0_2_3MyFalse_1QVal_Bool_bufchan_r;
  assign es_0_2_3MyFalse_1QVal_Bool_r = ((! es_0_2_3MyFalse_1QVal_Bool_bufchan_d[0]) || es_0_2_3MyFalse_1QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_3MyFalse_1QVal_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_0_2_3MyFalse_1QVal_Bool_r)
        es_0_2_3MyFalse_1QVal_Bool_bufchan_d <= es_0_2_3MyFalse_1QVal_Bool_d;
  QTree_Bool_t es_0_2_3MyFalse_1QVal_Bool_bufchan_buf;
  assign es_0_2_3MyFalse_1QVal_Bool_bufchan_r = (! es_0_2_3MyFalse_1QVal_Bool_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (es_0_2_3MyFalse_1QVal_Bool_bufchan_buf[0] ? es_0_2_3MyFalse_1QVal_Bool_bufchan_buf :
                                   es_0_2_3MyFalse_1QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_0_2_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && es_0_2_3MyFalse_1QVal_Bool_bufchan_buf[0]))
        es_0_2_3MyFalse_1QVal_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! es_0_2_3MyFalse_1QVal_Bool_bufchan_buf[0])))
        es_0_2_3MyFalse_1QVal_Bool_bufchan_buf <= es_0_2_3MyFalse_1QVal_Bool_bufchan_d;
  
  /* buf (Ty MyDTBool_Nat) : (gacR_2_2,MyDTBool_Nat) > (gacR_2_2_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t gacR_2_2_bufchan_d;
  logic gacR_2_2_bufchan_r;
  assign gacR_2_2_r = ((! gacR_2_2_bufchan_d[0]) || gacR_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_2_2_bufchan_d <= 1'd0;
    else if (gacR_2_2_r) gacR_2_2_bufchan_d <= gacR_2_2_d;
  MyDTBool_Nat_t gacR_2_2_bufchan_buf;
  assign gacR_2_2_bufchan_r = (! gacR_2_2_bufchan_buf[0]);
  assign gacR_2_2_argbuf_d = (gacR_2_2_bufchan_buf[0] ? gacR_2_2_bufchan_buf :
                              gacR_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacR_2_2_argbuf_r && gacR_2_2_bufchan_buf[0]))
        gacR_2_2_bufchan_buf <= 1'd0;
      else if (((! gacR_2_2_argbuf_r) && (! gacR_2_2_bufchan_buf[0])))
        gacR_2_2_bufchan_buf <= gacR_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Nat) : (gacR_2_destruct,MyDTBool_Nat) > [(gacR_2_1,MyDTBool_Nat),
                                                           (gacR_2_2,MyDTBool_Nat)] */
  logic [1:0] gacR_2_destruct_emitted;
  logic [1:0] gacR_2_destruct_done;
  assign gacR_2_1_d = (gacR_2_destruct_d[0] && (! gacR_2_destruct_emitted[0]));
  assign gacR_2_2_d = (gacR_2_destruct_d[0] && (! gacR_2_destruct_emitted[1]));
  assign gacR_2_destruct_done = (gacR_2_destruct_emitted | ({gacR_2_2_d[0],
                                                             gacR_2_1_d[0]} & {gacR_2_2_r,
                                                                               gacR_2_1_r}));
  assign gacR_2_destruct_r = (& gacR_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_2_destruct_emitted <= 2'd0;
    else
      gacR_2_destruct_emitted <= (gacR_2_destruct_r ? 2'd0 :
                                  gacR_2_destruct_done);
  
  /* buf (Ty MyDTBool_Nat) : (gacR_3_2,MyDTBool_Nat) > (gacR_3_2_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t gacR_3_2_bufchan_d;
  logic gacR_3_2_bufchan_r;
  assign gacR_3_2_r = ((! gacR_3_2_bufchan_d[0]) || gacR_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_3_2_bufchan_d <= 1'd0;
    else if (gacR_3_2_r) gacR_3_2_bufchan_d <= gacR_3_2_d;
  MyDTBool_Nat_t gacR_3_2_bufchan_buf;
  assign gacR_3_2_bufchan_r = (! gacR_3_2_bufchan_buf[0]);
  assign gacR_3_2_argbuf_d = (gacR_3_2_bufchan_buf[0] ? gacR_3_2_bufchan_buf :
                              gacR_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacR_3_2_argbuf_r && gacR_3_2_bufchan_buf[0]))
        gacR_3_2_bufchan_buf <= 1'd0;
      else if (((! gacR_3_2_argbuf_r) && (! gacR_3_2_bufchan_buf[0])))
        gacR_3_2_bufchan_buf <= gacR_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Nat) : (gacR_3_destruct,MyDTBool_Nat) > [(gacR_3_1,MyDTBool_Nat),
                                                           (gacR_3_2,MyDTBool_Nat)] */
  logic [1:0] gacR_3_destruct_emitted;
  logic [1:0] gacR_3_destruct_done;
  assign gacR_3_1_d = (gacR_3_destruct_d[0] && (! gacR_3_destruct_emitted[0]));
  assign gacR_3_2_d = (gacR_3_destruct_d[0] && (! gacR_3_destruct_emitted[1]));
  assign gacR_3_destruct_done = (gacR_3_destruct_emitted | ({gacR_3_2_d[0],
                                                             gacR_3_1_d[0]} & {gacR_3_2_r,
                                                                               gacR_3_1_r}));
  assign gacR_3_destruct_r = (& gacR_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_3_destruct_emitted <= 2'd0;
    else
      gacR_3_destruct_emitted <= (gacR_3_destruct_r ? 2'd0 :
                                  gacR_3_destruct_done);
  
  /* buf (Ty MyDTBool_Nat) : (gacR_4_destruct,MyDTBool_Nat) > (gacR_4_1_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t gacR_4_destruct_bufchan_d;
  logic gacR_4_destruct_bufchan_r;
  assign gacR_4_destruct_r = ((! gacR_4_destruct_bufchan_d[0]) || gacR_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacR_4_destruct_r)
        gacR_4_destruct_bufchan_d <= gacR_4_destruct_d;
  MyDTBool_Nat_t gacR_4_destruct_bufchan_buf;
  assign gacR_4_destruct_bufchan_r = (! gacR_4_destruct_bufchan_buf[0]);
  assign gacR_4_1_argbuf_d = (gacR_4_destruct_bufchan_buf[0] ? gacR_4_destruct_bufchan_buf :
                              gacR_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacR_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacR_4_1_argbuf_r && gacR_4_destruct_bufchan_buf[0]))
        gacR_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacR_4_1_argbuf_r) && (! gacR_4_destruct_bufchan_buf[0])))
        gacR_4_destruct_bufchan_buf <= gacR_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacZ_2_2,MyDTBool_Bool_Bool) > (gacZ_2_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacZ_2_2_bufchan_d;
  logic gacZ_2_2_bufchan_r;
  assign gacZ_2_2_r = ((! gacZ_2_2_bufchan_d[0]) || gacZ_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_2_2_bufchan_d <= 1'd0;
    else if (gacZ_2_2_r) gacZ_2_2_bufchan_d <= gacZ_2_2_d;
  MyDTBool_Bool_Bool_t gacZ_2_2_bufchan_buf;
  assign gacZ_2_2_bufchan_r = (! gacZ_2_2_bufchan_buf[0]);
  assign gacZ_2_2_argbuf_d = (gacZ_2_2_bufchan_buf[0] ? gacZ_2_2_bufchan_buf :
                              gacZ_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_2_2_bufchan_buf <= 1'd0;
    else
      if ((gacZ_2_2_argbuf_r && gacZ_2_2_bufchan_buf[0]))
        gacZ_2_2_bufchan_buf <= 1'd0;
      else if (((! gacZ_2_2_argbuf_r) && (! gacZ_2_2_bufchan_buf[0])))
        gacZ_2_2_bufchan_buf <= gacZ_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacZ_2_destruct,MyDTBool_Bool_Bool) > [(gacZ_2_1,MyDTBool_Bool_Bool),
                                                                       (gacZ_2_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacZ_2_destruct_emitted;
  logic [1:0] gacZ_2_destruct_done;
  assign gacZ_2_1_d = (gacZ_2_destruct_d[0] && (! gacZ_2_destruct_emitted[0]));
  assign gacZ_2_2_d = (gacZ_2_destruct_d[0] && (! gacZ_2_destruct_emitted[1]));
  assign gacZ_2_destruct_done = (gacZ_2_destruct_emitted | ({gacZ_2_2_d[0],
                                                             gacZ_2_1_d[0]} & {gacZ_2_2_r,
                                                                               gacZ_2_1_r}));
  assign gacZ_2_destruct_r = (& gacZ_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_2_destruct_emitted <= 2'd0;
    else
      gacZ_2_destruct_emitted <= (gacZ_2_destruct_r ? 2'd0 :
                                  gacZ_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacZ_3_2,MyDTBool_Bool_Bool) > (gacZ_3_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacZ_3_2_bufchan_d;
  logic gacZ_3_2_bufchan_r;
  assign gacZ_3_2_r = ((! gacZ_3_2_bufchan_d[0]) || gacZ_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_3_2_bufchan_d <= 1'd0;
    else if (gacZ_3_2_r) gacZ_3_2_bufchan_d <= gacZ_3_2_d;
  MyDTBool_Bool_Bool_t gacZ_3_2_bufchan_buf;
  assign gacZ_3_2_bufchan_r = (! gacZ_3_2_bufchan_buf[0]);
  assign gacZ_3_2_argbuf_d = (gacZ_3_2_bufchan_buf[0] ? gacZ_3_2_bufchan_buf :
                              gacZ_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_3_2_bufchan_buf <= 1'd0;
    else
      if ((gacZ_3_2_argbuf_r && gacZ_3_2_bufchan_buf[0]))
        gacZ_3_2_bufchan_buf <= 1'd0;
      else if (((! gacZ_3_2_argbuf_r) && (! gacZ_3_2_bufchan_buf[0])))
        gacZ_3_2_bufchan_buf <= gacZ_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gacZ_3_destruct,MyDTBool_Bool_Bool) > [(gacZ_3_1,MyDTBool_Bool_Bool),
                                                                       (gacZ_3_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gacZ_3_destruct_emitted;
  logic [1:0] gacZ_3_destruct_done;
  assign gacZ_3_1_d = (gacZ_3_destruct_d[0] && (! gacZ_3_destruct_emitted[0]));
  assign gacZ_3_2_d = (gacZ_3_destruct_d[0] && (! gacZ_3_destruct_emitted[1]));
  assign gacZ_3_destruct_done = (gacZ_3_destruct_emitted | ({gacZ_3_2_d[0],
                                                             gacZ_3_1_d[0]} & {gacZ_3_2_r,
                                                                               gacZ_3_1_r}));
  assign gacZ_3_destruct_r = (& gacZ_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_3_destruct_emitted <= 2'd0;
    else
      gacZ_3_destruct_emitted <= (gacZ_3_destruct_r ? 2'd0 :
                                  gacZ_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gacZ_4_destruct,MyDTBool_Bool_Bool) > (gacZ_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gacZ_4_destruct_bufchan_d;
  logic gacZ_4_destruct_bufchan_r;
  assign gacZ_4_destruct_r = ((! gacZ_4_destruct_bufchan_d[0]) || gacZ_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_4_destruct_bufchan_d <= 1'd0;
    else
      if (gacZ_4_destruct_r)
        gacZ_4_destruct_bufchan_d <= gacZ_4_destruct_d;
  MyDTBool_Bool_Bool_t gacZ_4_destruct_bufchan_buf;
  assign gacZ_4_destruct_bufchan_r = (! gacZ_4_destruct_bufchan_buf[0]);
  assign gacZ_4_1_argbuf_d = (gacZ_4_destruct_bufchan_buf[0] ? gacZ_4_destruct_bufchan_buf :
                              gacZ_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gacZ_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gacZ_4_1_argbuf_r && gacZ_4_destruct_bufchan_buf[0]))
        gacZ_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gacZ_4_1_argbuf_r) && (! gacZ_4_destruct_bufchan_buf[0])))
        gacZ_4_destruct_bufchan_buf <= gacZ_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gad8_2_2,MyDTBool_Bool_Bool) > (gad8_2_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gad8_2_2_bufchan_d;
  logic gad8_2_2_bufchan_r;
  assign gad8_2_2_r = ((! gad8_2_2_bufchan_d[0]) || gad8_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_2_2_bufchan_d <= 1'd0;
    else if (gad8_2_2_r) gad8_2_2_bufchan_d <= gad8_2_2_d;
  MyDTBool_Bool_Bool_t gad8_2_2_bufchan_buf;
  assign gad8_2_2_bufchan_r = (! gad8_2_2_bufchan_buf[0]);
  assign gad8_2_2_argbuf_d = (gad8_2_2_bufchan_buf[0] ? gad8_2_2_bufchan_buf :
                              gad8_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_2_2_bufchan_buf <= 1'd0;
    else
      if ((gad8_2_2_argbuf_r && gad8_2_2_bufchan_buf[0]))
        gad8_2_2_bufchan_buf <= 1'd0;
      else if (((! gad8_2_2_argbuf_r) && (! gad8_2_2_bufchan_buf[0])))
        gad8_2_2_bufchan_buf <= gad8_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gad8_2_destruct,MyDTBool_Bool_Bool) > [(gad8_2_1,MyDTBool_Bool_Bool),
                                                                       (gad8_2_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gad8_2_destruct_emitted;
  logic [1:0] gad8_2_destruct_done;
  assign gad8_2_1_d = (gad8_2_destruct_d[0] && (! gad8_2_destruct_emitted[0]));
  assign gad8_2_2_d = (gad8_2_destruct_d[0] && (! gad8_2_destruct_emitted[1]));
  assign gad8_2_destruct_done = (gad8_2_destruct_emitted | ({gad8_2_2_d[0],
                                                             gad8_2_1_d[0]} & {gad8_2_2_r,
                                                                               gad8_2_1_r}));
  assign gad8_2_destruct_r = (& gad8_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_2_destruct_emitted <= 2'd0;
    else
      gad8_2_destruct_emitted <= (gad8_2_destruct_r ? 2'd0 :
                                  gad8_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gad8_3_2,MyDTBool_Bool_Bool) > (gad8_3_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gad8_3_2_bufchan_d;
  logic gad8_3_2_bufchan_r;
  assign gad8_3_2_r = ((! gad8_3_2_bufchan_d[0]) || gad8_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_3_2_bufchan_d <= 1'd0;
    else if (gad8_3_2_r) gad8_3_2_bufchan_d <= gad8_3_2_d;
  MyDTBool_Bool_Bool_t gad8_3_2_bufchan_buf;
  assign gad8_3_2_bufchan_r = (! gad8_3_2_bufchan_buf[0]);
  assign gad8_3_2_argbuf_d = (gad8_3_2_bufchan_buf[0] ? gad8_3_2_bufchan_buf :
                              gad8_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_3_2_bufchan_buf <= 1'd0;
    else
      if ((gad8_3_2_argbuf_r && gad8_3_2_bufchan_buf[0]))
        gad8_3_2_bufchan_buf <= 1'd0;
      else if (((! gad8_3_2_argbuf_r) && (! gad8_3_2_bufchan_buf[0])))
        gad8_3_2_bufchan_buf <= gad8_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (gad8_3_destruct,MyDTBool_Bool_Bool) > [(gad8_3_1,MyDTBool_Bool_Bool),
                                                                       (gad8_3_2,MyDTBool_Bool_Bool)] */
  logic [1:0] gad8_3_destruct_emitted;
  logic [1:0] gad8_3_destruct_done;
  assign gad8_3_1_d = (gad8_3_destruct_d[0] && (! gad8_3_destruct_emitted[0]));
  assign gad8_3_2_d = (gad8_3_destruct_d[0] && (! gad8_3_destruct_emitted[1]));
  assign gad8_3_destruct_done = (gad8_3_destruct_emitted | ({gad8_3_2_d[0],
                                                             gad8_3_1_d[0]} & {gad8_3_2_r,
                                                                               gad8_3_1_r}));
  assign gad8_3_destruct_r = (& gad8_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_3_destruct_emitted <= 2'd0;
    else
      gad8_3_destruct_emitted <= (gad8_3_destruct_r ? 2'd0 :
                                  gad8_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (gad8_4_destruct,MyDTBool_Bool_Bool) > (gad8_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t gad8_4_destruct_bufchan_d;
  logic gad8_4_destruct_bufchan_r;
  assign gad8_4_destruct_r = ((! gad8_4_destruct_bufchan_d[0]) || gad8_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_4_destruct_bufchan_d <= 1'd0;
    else
      if (gad8_4_destruct_r)
        gad8_4_destruct_bufchan_d <= gad8_4_destruct_d;
  MyDTBool_Bool_Bool_t gad8_4_destruct_bufchan_buf;
  assign gad8_4_destruct_bufchan_r = (! gad8_4_destruct_bufchan_buf[0]);
  assign gad8_4_1_argbuf_d = (gad8_4_destruct_bufchan_buf[0] ? gad8_4_destruct_bufchan_buf :
                              gad8_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) gad8_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((gad8_4_1_argbuf_r && gad8_4_destruct_bufchan_buf[0]))
        gad8_4_destruct_bufchan_buf <= 1'd0;
      else if (((! gad8_4_1_argbuf_r) && (! gad8_4_destruct_bufchan_buf[0])))
        gad8_4_destruct_bufchan_buf <= gad8_4_destruct_bufchan_d;
  
  /* dcon (Ty MyDTBool_Nat,
      Dcon Dcon_to_nat) : [(go_1,Go)] > (go_1Dcon_to_nat,MyDTBool_Nat) */
  assign go_1Dcon_to_nat_d = Dcon_to_nat_dc((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(go_1Dcon_to_nat_r && go_1Dcon_to_nat_d[0])}};
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lkron_kron_Bool_Bool_Boolsbos) : [(go_10_1,Go)] > (go_10_1Lkron_kron_Bool_Bool_Boolsbos,CTkron_kron_Bool_Bool_Bool) */
  assign go_10_1Lkron_kron_Bool_Bool_Boolsbos_d = Lkron_kron_Bool_Bool_Boolsbos_dc((& {go_10_1_d[0]}), go_10_1_d);
  assign {go_10_1_r} = {1 {(go_10_1Lkron_kron_Bool_Bool_Boolsbos_r && go_10_1Lkron_kron_Bool_Bool_Boolsbos_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (go_10_1Lkron_kron_Bool_Bool_Boolsbos,CTkron_kron_Bool_Bool_Bool) > (lizzieLet21_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d;
  logic go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r;
  assign go_10_1Lkron_kron_Bool_Bool_Boolsbos_r = ((! go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d[0]) || go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d <= {83'd0, 1'd0};
    else
      if (go_10_1Lkron_kron_Bool_Bool_Boolsbos_r)
        go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d <= go_10_1Lkron_kron_Bool_Bool_Boolsbos_d;
  CTkron_kron_Bool_Bool_Bool_t go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf;
  assign go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_r = (! go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0] ? go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf :
                                   go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= {83'd0, 1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0]))
        go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= {83'd0, 1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf[0])))
        go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_buf <= go_10_1Lkron_kron_Bool_Bool_Boolsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_10_2,Go) > (go_10_2_argbuf,Go) */
  Go_t go_10_2_bufchan_d;
  logic go_10_2_bufchan_r;
  assign go_10_2_r = ((! go_10_2_bufchan_d[0]) || go_10_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_2_bufchan_d <= 1'd0;
    else if (go_10_2_r) go_10_2_bufchan_d <= go_10_2_d;
  Go_t go_10_2_bufchan_buf;
  assign go_10_2_bufchan_r = (! go_10_2_bufchan_buf[0]);
  assign go_10_2_argbuf_d = (go_10_2_bufchan_buf[0] ? go_10_2_bufchan_buf :
                             go_10_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_2_bufchan_buf <= 1'd0;
    else
      if ((go_10_2_argbuf_r && go_10_2_bufchan_buf[0]))
        go_10_2_bufchan_buf <= 1'd0;
      else if (((! go_10_2_argbuf_r) && (! go_10_2_bufchan_buf[0])))
        go_10_2_bufchan_buf <= go_10_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) : [(go_10_2_argbuf,Go),
                                                                                                                                         (isZad7_1_1_argbuf,MyDTBool_Bool),
                                                                                                                                         (gad8_1_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                                                         (m1ad9_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                                         (m2ada_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                                         (lizzieLet14_1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool) */
  assign call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_dc((& {go_10_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       isZad7_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       gad8_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       m1ad9_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       m2ada_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                       lizzieLet14_1_1_argbuf_d[0]}), go_10_2_argbuf_d, isZad7_1_1_argbuf_d, gad8_1_1_argbuf_d, m1ad9_1_1_argbuf_d, m2ada_1_1_argbuf_d, lizzieLet14_1_1_argbuf_d);
  assign {go_10_2_argbuf_r,
          isZad7_1_1_argbuf_r,
          gad8_1_1_argbuf_r,
          m1ad9_1_1_argbuf_r,
          m2ada_1_1_argbuf_r,
          lizzieLet14_1_1_argbuf_r} = {6 {(call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_r && call_kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTkron_kron_Bool_Bool_Bool_1_d[0])}};
  
  /* dcon (Ty CTmain_map'_Bool_Nat,
      Dcon Lmain_map'_Bool_Natsbos) : [(go_11_1,Go)] > (go_11_1Lmain_map'_Bool_Natsbos,CTmain_map'_Bool_Nat) */
  assign \go_11_1Lmain_map'_Bool_Natsbos_d  = \Lmain_map'_Bool_Natsbos_dc ((& {go_11_1_d[0]}), go_11_1_d);
  assign {go_11_1_r} = {1 {(\go_11_1Lmain_map'_Bool_Natsbos_r  && \go_11_1Lmain_map'_Bool_Natsbos_d [0])}};
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (go_11_1Lmain_map'_Bool_Natsbos,CTmain_map'_Bool_Nat) > (lizzieLet22_1_argbuf,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d ;
  logic \go_11_1Lmain_map'_Bool_Natsbos_bufchan_r ;
  assign \go_11_1Lmain_map'_Bool_Natsbos_r  = ((! \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d [0]) || \go_11_1Lmain_map'_Bool_Natsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d  <= {67'd0, 1'd0};
    else
      if (\go_11_1Lmain_map'_Bool_Natsbos_r )
        \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d  <= \go_11_1Lmain_map'_Bool_Natsbos_d ;
  \CTmain_map'_Bool_Nat_t  \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf ;
  assign \go_11_1Lmain_map'_Bool_Natsbos_bufchan_r  = (! \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf [0]);
  assign lizzieLet22_1_argbuf_d = (\go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf [0] ? \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf  :
                                   \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf  <= {67'd0, 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf [0]))
        \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf  <= {67'd0, 1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf [0])))
        \go_11_1Lmain_map'_Bool_Natsbos_bufchan_buf  <= \go_11_1Lmain_map'_Bool_Natsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_11_2,Go) > (go_11_2_argbuf,Go) */
  Go_t go_11_2_bufchan_d;
  logic go_11_2_bufchan_r;
  assign go_11_2_r = ((! go_11_2_bufchan_d[0]) || go_11_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_2_bufchan_d <= 1'd0;
    else if (go_11_2_r) go_11_2_bufchan_d <= go_11_2_d;
  Go_t go_11_2_bufchan_buf;
  assign go_11_2_bufchan_r = (! go_11_2_bufchan_buf[0]);
  assign go_11_2_argbuf_d = (go_11_2_bufchan_buf[0] ? go_11_2_bufchan_buf :
                             go_11_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_2_bufchan_buf <= 1'd0;
    else
      if ((go_11_2_argbuf_r && go_11_2_bufchan_buf[0]))
        go_11_2_bufchan_buf <= 1'd0;
      else if (((! go_11_2_argbuf_r) && (! go_11_2_bufchan_buf[0])))
        go_11_2_bufchan_buf <= go_11_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat,
      Dcon TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat) : [(go_11_2_argbuf,Go),
                                                                                                       (isZacQ_1_1_argbuf,MyDTNat_Bool),
                                                                                                       (gacR_1_1_argbuf,MyDTBool_Nat),
                                                                                                       (macS_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                       (lizzieLet5_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat)] > (call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1,TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat) */
  assign \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d  = \TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_dc ((& {go_11_2_argbuf_d[0],
                                                                                                                                                                                                                                 isZacQ_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 gacR_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 macS_1_1_argbuf_d[0],
                                                                                                                                                                                                                                 lizzieLet5_1_1_argbuf_d[0]}), go_11_2_argbuf_d, isZacQ_1_1_argbuf_d, gacR_1_1_argbuf_d, macS_1_1_argbuf_d, lizzieLet5_1_1_argbuf_d);
  assign {go_11_2_argbuf_r,
          isZacQ_1_1_argbuf_r,
          gacR_1_1_argbuf_r,
          macS_1_1_argbuf_r,
          lizzieLet5_1_1_argbuf_r} = {5 {(\call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_r  && \call_main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool___Pointer_CTmain_map'_Bool_Nat_1_d [0])}};
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lmap''_map''_Bool_Bool_Boolsbos) : [(go_12_1,Go)] > (go_12_1Lmap''_map''_Bool_Bool_Boolsbos,CTmap''_map''_Bool_Bool_Bool) */
  assign \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_d  = \Lmap''_map''_Bool_Bool_Boolsbos_dc ((& {go_12_1_d[0]}), go_12_1_d);
  assign {go_12_1_r} = {1 {(\go_12_1Lmap''_map''_Bool_Bool_Boolsbos_r  && \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (go_12_1Lmap''_map''_Bool_Bool_Boolsbos,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet23_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d ;
  logic \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r ;
  assign \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_r  = ((! \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d [0]) || \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d  <= {68'd0,
                                                             1'd0};
    else
      if (\go_12_1Lmap''_map''_Bool_Bool_Boolsbos_r )
        \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d  <= \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf ;
  assign \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_r  = (! \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0]);
  assign lizzieLet23_1_argbuf_d = (\go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0] ? \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  :
                                   \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= {68'd0,
                                                               1'd0};
    else
      if ((lizzieLet23_1_argbuf_r && \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0]))
        \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= {68'd0,
                                                                 1'd0};
      else if (((! lizzieLet23_1_argbuf_r) && (! \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf [0])))
        \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_buf  <= \go_12_1Lmap''_map''_Bool_Bool_Boolsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_12_2,Go) > (go_12_2_argbuf,Go) */
  Go_t go_12_2_bufchan_d;
  logic go_12_2_bufchan_r;
  assign go_12_2_r = ((! go_12_2_bufchan_d[0]) || go_12_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_d <= 1'd0;
    else if (go_12_2_r) go_12_2_bufchan_d <= go_12_2_d;
  Go_t go_12_2_bufchan_buf;
  assign go_12_2_bufchan_r = (! go_12_2_bufchan_buf[0]);
  assign go_12_2_argbuf_d = (go_12_2_bufchan_buf[0] ? go_12_2_bufchan_buf :
                             go_12_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_2_bufchan_buf <= 1'd0;
    else
      if ((go_12_2_argbuf_r && go_12_2_bufchan_buf[0]))
        go_12_2_bufchan_buf <= 1'd0;
      else if (((! go_12_2_argbuf_r) && (! go_12_2_bufchan_buf[0])))
        go_12_2_bufchan_buf <= go_12_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) : [(go_12_2_argbuf,Go),
                                                                                                                               (isZacY_1_1_argbuf,MyDTBool_Bool),
                                                                                                                               (gacZ_1_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                                               (v'ad0_1_1_argbuf,MyBool),
                                                                                                                               (mad1_1_1_argbuf,Pointer_QTree_Bool),
                                                                                                                               (lizzieLet10_1_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool) */
  assign \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d  = \TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_dc ((& {go_12_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                         isZacY_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         gacZ_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         \v'ad0_1_1_argbuf_d [0],
                                                                                                                                                                                                                                                                                         mad1_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                         lizzieLet10_1_1_argbuf_d[0]}), go_12_2_argbuf_d, isZacY_1_1_argbuf_d, gacZ_1_1_argbuf_d, \v'ad0_1_1_argbuf_d , mad1_1_1_argbuf_d, lizzieLet10_1_1_argbuf_d);
  assign {go_12_2_argbuf_r,
          isZacY_1_1_argbuf_r,
          gacZ_1_1_argbuf_r,
          \v'ad0_1_1_argbuf_r ,
          mad1_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = {6 {(\call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_r  && \call_map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool___Pointer_CTmap''_map''_Bool_Bool_Bool_1_d [0])}};
  
  /* fork (Ty C4) : (go_13_goMux_choice,C4) > [(go_13_goMux_choice_1,C4),
                                          (go_13_goMux_choice_2,C4)] */
  logic [1:0] go_13_goMux_choice_emitted;
  logic [1:0] go_13_goMux_choice_done;
  assign go_13_goMux_choice_1_d = {go_13_goMux_choice_d[2:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[0]))};
  assign go_13_goMux_choice_2_d = {go_13_goMux_choice_d[2:1],
                                   (go_13_goMux_choice_d[0] && (! go_13_goMux_choice_emitted[1]))};
  assign go_13_goMux_choice_done = (go_13_goMux_choice_emitted | ({go_13_goMux_choice_2_d[0],
                                                                   go_13_goMux_choice_1_d[0]} & {go_13_goMux_choice_2_r,
                                                                                                 go_13_goMux_choice_1_r}));
  assign go_13_goMux_choice_r = (& go_13_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_goMux_choice_emitted <= 2'd0;
    else
      go_13_goMux_choice_emitted <= (go_13_goMux_choice_r ? 2'd0 :
                                     go_13_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Pointer_QTree_Bool) : (go_13_goMux_choice_1,C4) [(lizzieLet11_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet12_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet13_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet11_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet12_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet13_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[16:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_13_goMux_choice_1_d[0])};
  assign go_13_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet13_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (go_13_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (go_13_goMux_choice_2,C4) [(lizzieLet2_7QNone_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (sc_0_6_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (lizzieLet2_7QVal_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                         (lizzieLet2_7QError_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (scfarg_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_13_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet2_7QNone_Bool_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet2_7QVal_Bool_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet2_7QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_13_goMux_choice_2_d[0])};
  assign go_13_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet2_7QError_Bool_1_argbuf_r,
          lizzieLet2_7QVal_Bool_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet2_7QNone_Bool_1_argbuf_r} = (go_13_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                                4'd0);
  
  /* fork (Ty C5) : (go_14_goMux_choice,C5) > [(go_14_goMux_choice_1,C5),
                                          (go_14_goMux_choice_2,C5)] */
  logic [1:0] go_14_goMux_choice_emitted;
  logic [1:0] go_14_goMux_choice_done;
  assign go_14_goMux_choice_1_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[0]))};
  assign go_14_goMux_choice_2_d = {go_14_goMux_choice_d[3:1],
                                   (go_14_goMux_choice_d[0] && (! go_14_goMux_choice_emitted[1]))};
  assign go_14_goMux_choice_done = (go_14_goMux_choice_emitted | ({go_14_goMux_choice_2_d[0],
                                                                   go_14_goMux_choice_1_d[0]} & {go_14_goMux_choice_2_r,
                                                                                                 go_14_goMux_choice_1_r}));
  assign go_14_goMux_choice_r = (& go_14_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_goMux_choice_emitted <= 2'd0;
    else
      go_14_goMux_choice_emitted <= (go_14_goMux_choice_r ? 2'd0 :
                                     go_14_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Nat) : (go_14_goMux_choice_1,C5) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Nat),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Nat),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Nat),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Nat),
                                                        (lizzieLet4_1_1_argbuf,Pointer_QTree_Nat)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Nat) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [4:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet3_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet4_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_14_goMux_choice_1_d[0])};
  assign go_14_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet4_1_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_14_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Bool_Nat) : (go_14_goMux_choice_2,C5) [(lizzieLet6_6QNone_Bool_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                   (sc_0_10_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                   (es_0_1_2MyFalse_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                   (es_0_1_2MyTrue_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                   (lizzieLet6_6QError_Bool_1_argbuf,Pointer_CTmain_map'_Bool_Nat)] > (scfarg_0_1_goMux_mux,Pointer_CTmain_map'_Bool_Nat) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [4:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_14_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet6_6QNone_Bool_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd2,
                                                                   sc_0_10_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd4,
                                                                   es_0_1_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd8,
                                                                   es_0_1_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet6_6QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_14_goMux_choice_2_d[0])};
  assign go_14_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_6QError_Bool_1_argbuf_r,
          es_0_1_2MyTrue_1_argbuf_r,
          es_0_1_2MyFalse_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet6_6QNone_Bool_1_argbuf_r} = (go_14_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                                5'd0);
  
  /* fork (Ty C5) : (go_15_goMux_choice,C5) > [(go_15_goMux_choice_1,C5),
                                          (go_15_goMux_choice_2,C5)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[3:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[3:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_15_goMux_choice_1,C5) [(lizzieLet6_1_1_argbuf,Pointer_QTree_Bool),
                                                         (contRet_0_2_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool),
                                                         (lizzieLet9_1_1_argbuf,Pointer_QTree_Bool)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [4:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet6_1_1_argbuf_d};
      3'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   contRet_0_2_1_argbuf_d};
      3'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   lizzieLet7_1_1_argbuf_d};
      3'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   lizzieLet8_1_1_argbuf_d};
      3'd4:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet9_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (go_15_goMux_choice_2,C5) [(lizzieLet12_1_6QNone_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (sc_0_14_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (es_0_2_2MyFalse_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (es_0_2_2MyTrue_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                           (lizzieLet12_1_6QError_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (scfarg_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [4:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd1,
                                                                   lizzieLet12_1_6QNone_Bool_1_argbuf_d};
      3'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd2,
                                                                   sc_0_14_1_argbuf_d};
      3'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd4,
                                                                   es_0_2_2MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd8,
                                                                   es_0_2_2MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet12_1_6QError_Bool_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {5'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet12_1_6QError_Bool_1_argbuf_r,
          es_0_2_2MyTrue_1_argbuf_r,
          es_0_2_2MyFalse_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet12_1_6QNone_Bool_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                   5'd0);
  
  /* buf (Ty Nat) : (go_16_1Zero,Nat) > (lizzieLet39_1_argbuf,Nat) */
  Nat_t go_16_1Zero_bufchan_d;
  logic go_16_1Zero_bufchan_r;
  assign go_16_1Zero_r = ((! go_16_1Zero_bufchan_d[0]) || go_16_1Zero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_1Zero_bufchan_d <= {17'd0, 1'd0};
    else if (go_16_1Zero_r) go_16_1Zero_bufchan_d <= go_16_1Zero_d;
  Nat_t go_16_1Zero_bufchan_buf;
  assign go_16_1Zero_bufchan_r = (! go_16_1Zero_bufchan_buf[0]);
  assign lizzieLet39_1_argbuf_d = (go_16_1Zero_bufchan_buf[0] ? go_16_1Zero_bufchan_buf :
                                   go_16_1Zero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_1Zero_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((lizzieLet39_1_argbuf_r && go_16_1Zero_bufchan_buf[0]))
        go_16_1Zero_bufchan_buf <= {17'd0, 1'd0};
      else if (((! lizzieLet39_1_argbuf_r) && (! go_16_1Zero_bufchan_buf[0])))
        go_16_1Zero_bufchan_buf <= go_16_1Zero_bufchan_d;
  
  /* buf (Ty MyDTBool_Nat) : (go_1Dcon_to_nat,MyDTBool_Nat) > (es_1_1_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t go_1Dcon_to_nat_bufchan_d;
  logic go_1Dcon_to_nat_bufchan_r;
  assign go_1Dcon_to_nat_r = ((! go_1Dcon_to_nat_bufchan_d[0]) || go_1Dcon_to_nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1Dcon_to_nat_bufchan_d <= 1'd0;
    else
      if (go_1Dcon_to_nat_r)
        go_1Dcon_to_nat_bufchan_d <= go_1Dcon_to_nat_d;
  MyDTBool_Nat_t go_1Dcon_to_nat_bufchan_buf;
  assign go_1Dcon_to_nat_bufchan_r = (! go_1Dcon_to_nat_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (go_1Dcon_to_nat_bufchan_buf[0] ? go_1Dcon_to_nat_bufchan_buf :
                            go_1Dcon_to_nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1Dcon_to_nat_bufchan_buf <= 1'd0;
    else
      if ((es_1_1_argbuf_r && go_1Dcon_to_nat_bufchan_buf[0]))
        go_1Dcon_to_nat_bufchan_buf <= 1'd0;
      else if (((! es_1_1_argbuf_r) && (! go_1Dcon_to_nat_bufchan_buf[0])))
        go_1Dcon_to_nat_bufchan_buf <= go_1Dcon_to_nat_bufchan_d;
  
  /* dcon (Ty MyDTNat_Bool,
      Dcon Dcon_is_z_nut) : [(go_2,Go)] > (go_2Dcon_is_z_nut,MyDTNat_Bool) */
  assign go_2Dcon_is_z_nut_d = Dcon_is_z_nut_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_is_z_nut_r && go_2Dcon_is_z_nut_d[0])}};
  
  /* buf (Ty MyDTNat_Bool) : (go_2Dcon_is_z_nut,MyDTNat_Bool) > (es_0_1_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t go_2Dcon_is_z_nut_bufchan_d;
  logic go_2Dcon_is_z_nut_bufchan_r;
  assign go_2Dcon_is_z_nut_r = ((! go_2Dcon_is_z_nut_bufchan_d[0]) || go_2Dcon_is_z_nut_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_is_z_nut_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_is_z_nut_r)
        go_2Dcon_is_z_nut_bufchan_d <= go_2Dcon_is_z_nut_d;
  MyDTNat_Bool_t go_2Dcon_is_z_nut_bufchan_buf;
  assign go_2Dcon_is_z_nut_bufchan_r = (! go_2Dcon_is_z_nut_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (go_2Dcon_is_z_nut_bufchan_buf[0] ? go_2Dcon_is_z_nut_bufchan_buf :
                            go_2Dcon_is_z_nut_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_is_z_nut_bufchan_buf <= 1'd0;
    else
      if ((es_0_1_argbuf_r && go_2Dcon_is_z_nut_bufchan_buf[0]))
        go_2Dcon_is_z_nut_bufchan_buf <= 1'd0;
      else if (((! es_0_1_argbuf_r) && (! go_2Dcon_is_z_nut_bufchan_buf[0])))
        go_2Dcon_is_z_nut_bufchan_buf <= go_2Dcon_is_z_nut_bufchan_d;
  
  /* dcon (Ty MyDTBool_Bool_Bool,
      Dcon Dcon_&&) : [(go_3,Go)] > (go_3Dcon_&&,MyDTBool_Bool_Bool) */
  assign \go_3Dcon_&&_d  = \Dcon_&&_dc ((& {go_3_d[0]}), go_3_d);
  assign {go_3_r} = {1 {(\go_3Dcon_&&_r  && \go_3Dcon_&&_d [0])}};
  
  /* buf (Ty MyDTBool_Bool_Bool) : (go_3Dcon_&&,MyDTBool_Bool_Bool) > (es_4_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \go_3Dcon_&&_bufchan_d ;
  logic \go_3Dcon_&&_bufchan_r ;
  assign \go_3Dcon_&&_r  = ((! \go_3Dcon_&&_bufchan_d [0]) || \go_3Dcon_&&_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_3Dcon_&&_bufchan_d  <= 1'd0;
    else
      if (\go_3Dcon_&&_r ) \go_3Dcon_&&_bufchan_d  <= \go_3Dcon_&&_d ;
  MyDTBool_Bool_Bool_t \go_3Dcon_&&_bufchan_buf ;
  assign \go_3Dcon_&&_bufchan_r  = (! \go_3Dcon_&&_bufchan_buf [0]);
  assign es_4_1_argbuf_d = (\go_3Dcon_&&_bufchan_buf [0] ? \go_3Dcon_&&_bufchan_buf  :
                            \go_3Dcon_&&_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_3Dcon_&&_bufchan_buf  <= 1'd0;
    else
      if ((es_4_1_argbuf_r && \go_3Dcon_&&_bufchan_buf [0]))
        \go_3Dcon_&&_bufchan_buf  <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! \go_3Dcon_&&_bufchan_buf [0])))
        \go_3Dcon_&&_bufchan_buf  <= \go_3Dcon_&&_bufchan_d ;
  
  /* dcon (Ty MyDTBool_Bool,
      Dcon Dcon_main1) : [(go_4,Go)] > (go_4Dcon_main1,MyDTBool_Bool) */
  assign go_4Dcon_main1_d = Dcon_main1_dc((& {go_4_d[0]}), go_4_d);
  assign {go_4_r} = {1 {(go_4Dcon_main1_r && go_4Dcon_main1_d[0])}};
  
  /* buf (Ty MyDTBool_Bool) : (go_4Dcon_main1,MyDTBool_Bool) > (es_3_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t go_4Dcon_main1_bufchan_d;
  logic go_4Dcon_main1_bufchan_r;
  assign go_4Dcon_main1_r = ((! go_4Dcon_main1_bufchan_d[0]) || go_4Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_4Dcon_main1_r) go_4Dcon_main1_bufchan_d <= go_4Dcon_main1_d;
  MyDTBool_Bool_t go_4Dcon_main1_bufchan_buf;
  assign go_4Dcon_main1_bufchan_r = (! go_4Dcon_main1_bufchan_buf[0]);
  assign es_3_1_argbuf_d = (go_4Dcon_main1_bufchan_buf[0] ? go_4Dcon_main1_bufchan_buf :
                            go_4Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_3_1_argbuf_r && go_4Dcon_main1_bufchan_buf[0]))
        go_4Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! go_4Dcon_main1_bufchan_buf[0])))
        go_4Dcon_main1_bufchan_buf <= go_4Dcon_main1_bufchan_d;
  
  /* buf (Ty Go) : (go_5,Go) > (go_5_argbuf,Go) */
  Go_t go_5_bufchan_d;
  logic go_5_bufchan_r;
  assign go_5_r = ((! go_5_bufchan_d[0]) || go_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_d <= 1'd0;
    else if (go_5_r) go_5_bufchan_d <= go_5_d;
  Go_t go_5_bufchan_buf;
  assign go_5_bufchan_r = (! go_5_bufchan_buf[0]);
  assign go_5_argbuf_d = (go_5_bufchan_buf[0] ? go_5_bufchan_buf :
                          go_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_buf <= 1'd0;
    else
      if ((go_5_argbuf_r && go_5_bufchan_buf[0]))
        go_5_bufchan_buf <= 1'd0;
      else if (((! go_5_argbuf_r) && (! go_5_bufchan_buf[0])))
        go_5_bufchan_buf <= go_5_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : [(go_5_argbuf,Go),
                                                                                                    (es_3_1_argbuf,MyDTBool_Bool),
                                                                                                    (es_4_1_argbuf,MyDTBool_Bool_Bool),
                                                                                                    (m1adn_0,Pointer_QTree_Bool),
                                                                                                    (m2ado_1,Pointer_QTree_Bool)] > (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) */
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_dc((& {go_5_argbuf_d[0],
                                                                                                                                                                                                                        es_3_1_argbuf_d[0],
                                                                                                                                                                                                                        es_4_1_argbuf_d[0],
                                                                                                                                                                                                                        m1adn_0_d[0],
                                                                                                                                                                                                                        m2ado_1_d[0]}), go_5_argbuf_d, es_3_1_argbuf_d, es_4_1_argbuf_d, m1adn_0_d, m2ado_1_d);
  assign {go_5_argbuf_r,
          es_3_1_argbuf_r,
          es_4_1_argbuf_r,
          m1adn_0_r,
          m2ado_1_r} = {5 {(kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0])}};
  
  /* buf (Ty Go) : (go_6,Go) > (go_6_argbuf,Go) */
  Go_t go_6_bufchan_d;
  logic go_6_bufchan_r;
  assign go_6_r = ((! go_6_bufchan_d[0]) || go_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_d <= 1'd0;
    else if (go_6_r) go_6_bufchan_d <= go_6_d;
  Go_t go_6_bufchan_buf;
  assign go_6_bufchan_r = (! go_6_bufchan_buf[0]);
  assign go_6_argbuf_d = (go_6_bufchan_buf[0] ? go_6_bufchan_buf :
                          go_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_buf <= 1'd0;
    else
      if ((go_6_argbuf_r && go_6_bufchan_buf[0]))
        go_6_bufchan_buf <= 1'd0;
      else if (((! go_6_argbuf_r) && (! go_6_bufchan_buf[0])))
        go_6_bufchan_buf <= go_6_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool,
      Dcon TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool) : [(go_6_argbuf,Go),
                                                                        (es_0_1_argbuf,MyDTNat_Bool),
                                                                        (es_1_1_argbuf,MyDTBool_Nat),
                                                                        (es_2_1_argbuf,Pointer_QTree_Bool)] > (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1,TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool) */
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d  = TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_dc((& {go_6_argbuf_d[0],
                                                                                                                                                            es_0_1_argbuf_d[0],
                                                                                                                                                            es_1_1_argbuf_d[0],
                                                                                                                                                            es_2_1_argbuf_d[0]}), go_6_argbuf_d, es_0_1_argbuf_d, es_1_1_argbuf_d, es_2_1_argbuf_d);
  assign {go_6_argbuf_r,
          es_0_1_argbuf_r,
          es_1_1_argbuf_r,
          es_2_1_argbuf_r} = {4 {(\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_r  && \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [0])}};
  
  /* fork (Ty C5) : (go_6_goMux_choice,C5) > [(go_6_goMux_choice_1,C5),
                                         (go_6_goMux_choice_2,C5),
                                         (go_6_goMux_choice_3,C5),
                                         (go_6_goMux_choice_4,C5),
                                         (go_6_goMux_choice_5,C5)] */
  logic [4:0] go_6_goMux_choice_emitted;
  logic [4:0] go_6_goMux_choice_done;
  assign go_6_goMux_choice_1_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[0]))};
  assign go_6_goMux_choice_2_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[1]))};
  assign go_6_goMux_choice_3_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[2]))};
  assign go_6_goMux_choice_4_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[3]))};
  assign go_6_goMux_choice_5_d = {go_6_goMux_choice_d[3:1],
                                  (go_6_goMux_choice_d[0] && (! go_6_goMux_choice_emitted[4]))};
  assign go_6_goMux_choice_done = (go_6_goMux_choice_emitted | ({go_6_goMux_choice_5_d[0],
                                                                 go_6_goMux_choice_4_d[0],
                                                                 go_6_goMux_choice_3_d[0],
                                                                 go_6_goMux_choice_2_d[0],
                                                                 go_6_goMux_choice_1_d[0]} & {go_6_goMux_choice_5_r,
                                                                                              go_6_goMux_choice_4_r,
                                                                                              go_6_goMux_choice_3_r,
                                                                                              go_6_goMux_choice_2_r,
                                                                                              go_6_goMux_choice_1_r}));
  assign go_6_goMux_choice_r = (& go_6_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_goMux_choice_emitted <= 5'd0;
    else
      go_6_goMux_choice_emitted <= (go_6_goMux_choice_r ? 5'd0 :
                                    go_6_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool) : (go_6_goMux_choice_1,C5) [(call_kron_kron_Bool_Bool_Bool_goMux2,MyDTBool_Bool),
                                                   (isZad7_2_2_argbuf,MyDTBool_Bool),
                                                   (isZad7_3_2_argbuf,MyDTBool_Bool),
                                                   (isZad7_4_1_argbuf,MyDTBool_Bool),
                                                   (lizzieLet2_5QNode_Bool_2_argbuf,MyDTBool_Bool)] > (isZad7_goMux_mux,MyDTBool_Bool) */
  logic [0:0] isZad7_goMux_mux_mux;
  logic [4:0] isZad7_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_1_d[3:1])
      3'd0:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd1,
                                                           call_kron_kron_Bool_Bool_Bool_goMux2_d};
      3'd1:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd2,
                                                           isZad7_2_2_argbuf_d};
      3'd2:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd4,
                                                           isZad7_3_2_argbuf_d};
      3'd3:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd8,
                                                           isZad7_4_1_argbuf_d};
      3'd4:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd16,
                                                           lizzieLet2_5QNode_Bool_2_argbuf_d};
      default:
        {isZad7_goMux_mux_onehot, isZad7_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZad7_goMux_mux_d = (isZad7_goMux_mux_mux[0] && go_6_goMux_choice_1_d[0]);
  assign go_6_goMux_choice_1_r = (isZad7_goMux_mux_d[0] && isZad7_goMux_mux_r);
  assign {lizzieLet2_5QNode_Bool_2_argbuf_r,
          isZad7_4_1_argbuf_r,
          isZad7_3_2_argbuf_r,
          isZad7_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux2_r} = (go_6_goMux_choice_1_r ? isZad7_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool_Bool) : (go_6_goMux_choice_2,C5) [(call_kron_kron_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool),
                                                        (gad8_2_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gad8_3_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gad8_4_1_argbuf,MyDTBool_Bool_Bool),
                                                        (lizzieLet2_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool)] > (gad8_goMux_mux,MyDTBool_Bool_Bool) */
  logic [0:0] gad8_goMux_mux_mux;
  logic [4:0] gad8_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_2_d[3:1])
      3'd0:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Bool_Bool_Bool_goMux3_d};
      3'd1:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd2,
                                                       gad8_2_2_argbuf_d};
      3'd2:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd4,
                                                       gad8_3_2_argbuf_d};
      3'd3:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd8,
                                                       gad8_4_1_argbuf_d};
      3'd4:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd16,
                                                       lizzieLet2_3QNode_Bool_2_argbuf_d};
      default:
        {gad8_goMux_mux_onehot, gad8_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gad8_goMux_mux_d = (gad8_goMux_mux_mux[0] && go_6_goMux_choice_2_d[0]);
  assign go_6_goMux_choice_2_r = (gad8_goMux_mux_d[0] && gad8_goMux_mux_r);
  assign {lizzieLet2_3QNode_Bool_2_argbuf_r,
          gad8_4_1_argbuf_r,
          gad8_3_2_argbuf_r,
          gad8_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux3_r} = (go_6_goMux_choice_2_r ? gad8_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_6_goMux_choice_3,C5) [(call_kron_kron_Bool_Bool_Bool_goMux4,Pointer_QTree_Bool),
                                                        (q3ade_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2add_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1adc_3_1_argbuf,Pointer_QTree_Bool),
                                                        (q4adf_1_argbuf,Pointer_QTree_Bool)] > (m1ad9_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m1ad9_goMux_mux_mux;
  logic [4:0] m1ad9_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_3_d[3:1])
      3'd0:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Bool_Bool_Bool_goMux4_d};
      3'd1:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd2,
                                                         q3ade_1_1_argbuf_d};
      3'd2:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd4,
                                                         q2add_2_1_argbuf_d};
      3'd3:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd8,
                                                         q1adc_3_1_argbuf_d};
      3'd4:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd16,
                                                         q4adf_1_argbuf_d};
      default:
        {m1ad9_goMux_mux_onehot, m1ad9_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1ad9_goMux_mux_d = {m1ad9_goMux_mux_mux[16:1],
                              (m1ad9_goMux_mux_mux[0] && go_6_goMux_choice_3_d[0])};
  assign go_6_goMux_choice_3_r = (m1ad9_goMux_mux_d[0] && m1ad9_goMux_mux_r);
  assign {q4adf_1_argbuf_r,
          q1adc_3_1_argbuf_r,
          q2add_2_1_argbuf_r,
          q3ade_1_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux4_r} = (go_6_goMux_choice_3_r ? m1ad9_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_6_goMux_choice_4,C5) [(call_kron_kron_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool),
                                                        (m2ada_2_2_argbuf,Pointer_QTree_Bool),
                                                        (m2ada_3_2_argbuf,Pointer_QTree_Bool),
                                                        (m2ada_4_1_argbuf,Pointer_QTree_Bool),
                                                        (lizzieLet2_6QNode_Bool_2_argbuf,Pointer_QTree_Bool)] > (m2ada_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] m2ada_goMux_mux_mux;
  logic [4:0] m2ada_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_4_d[3:1])
      3'd0:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd1,
                                                         call_kron_kron_Bool_Bool_Bool_goMux5_d};
      3'd1:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd2,
                                                         m2ada_2_2_argbuf_d};
      3'd2:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd4,
                                                         m2ada_3_2_argbuf_d};
      3'd3:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd8,
                                                         m2ada_4_1_argbuf_d};
      3'd4:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd16,
                                                         lizzieLet2_6QNode_Bool_2_argbuf_d};
      default:
        {m2ada_goMux_mux_onehot, m2ada_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ada_goMux_mux_d = {m2ada_goMux_mux_mux[16:1],
                              (m2ada_goMux_mux_mux[0] && go_6_goMux_choice_4_d[0])};
  assign go_6_goMux_choice_4_r = (m2ada_goMux_mux_d[0] && m2ada_goMux_mux_r);
  assign {lizzieLet2_6QNode_Bool_2_argbuf_r,
          m2ada_4_1_argbuf_r,
          m2ada_3_2_argbuf_r,
          m2ada_2_2_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux5_r} = (go_6_goMux_choice_4_r ? m2ada_goMux_mux_onehot :
                                                     5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (go_6_goMux_choice_5,C5) [(call_kron_kron_Bool_Bool_Bool_goMux6,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                        (sca3_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool)] > (sc_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_6_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_kron_kron_Bool_Bool_Bool_goMux6_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_6_goMux_choice_5_d[0])};
  assign go_6_goMux_choice_5_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_kron_kron_Bool_Bool_Bool_goMux6_r} = (go_6_goMux_choice_5_r ? sc_0_goMux_mux_onehot :
                                                     5'd0);
  
  /* fork (Ty C5) : (go_7_goMux_choice,C5) > [(go_7_goMux_choice_1,C5),
                                         (go_7_goMux_choice_2,C5),
                                         (go_7_goMux_choice_3,C5),
                                         (go_7_goMux_choice_4,C5)] */
  logic [3:0] go_7_goMux_choice_emitted;
  logic [3:0] go_7_goMux_choice_done;
  assign go_7_goMux_choice_1_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[0]))};
  assign go_7_goMux_choice_2_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[1]))};
  assign go_7_goMux_choice_3_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[2]))};
  assign go_7_goMux_choice_4_d = {go_7_goMux_choice_d[3:1],
                                  (go_7_goMux_choice_d[0] && (! go_7_goMux_choice_emitted[3]))};
  assign go_7_goMux_choice_done = (go_7_goMux_choice_emitted | ({go_7_goMux_choice_4_d[0],
                                                                 go_7_goMux_choice_3_d[0],
                                                                 go_7_goMux_choice_2_d[0],
                                                                 go_7_goMux_choice_1_d[0]} & {go_7_goMux_choice_4_r,
                                                                                              go_7_goMux_choice_3_r,
                                                                                              go_7_goMux_choice_2_r,
                                                                                              go_7_goMux_choice_1_r}));
  assign go_7_goMux_choice_r = (& go_7_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_goMux_choice_emitted <= 4'd0;
    else
      go_7_goMux_choice_emitted <= (go_7_goMux_choice_r ? 4'd0 :
                                    go_7_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTNat_Bool) : (go_7_goMux_choice_1,C5) [(call_main_map'_Bool_Nat_goMux2,MyDTNat_Bool),
                                                  (isZacQ_2_2_argbuf,MyDTNat_Bool),
                                                  (isZacQ_3_2_argbuf,MyDTNat_Bool),
                                                  (isZacQ_4_1_argbuf,MyDTNat_Bool),
                                                  (lizzieLet6_5QNode_Bool_2_argbuf,MyDTNat_Bool)] > (isZacQ_goMux_mux,MyDTNat_Bool) */
  logic [0:0] isZacQ_goMux_mux_mux;
  logic [4:0] isZacQ_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_1_d[3:1])
      3'd0:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Bool_Nat_goMux2_d };
      3'd1:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd2,
                                                           isZacQ_2_2_argbuf_d};
      3'd2:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd4,
                                                           isZacQ_3_2_argbuf_d};
      3'd3:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd8,
                                                           isZacQ_4_1_argbuf_d};
      3'd4:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd16,
                                                           lizzieLet6_5QNode_Bool_2_argbuf_d};
      default:
        {isZacQ_goMux_mux_onehot, isZacQ_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacQ_goMux_mux_d = (isZacQ_goMux_mux_mux[0] && go_7_goMux_choice_1_d[0]);
  assign go_7_goMux_choice_1_r = (isZacQ_goMux_mux_d[0] && isZacQ_goMux_mux_r);
  assign {lizzieLet6_5QNode_Bool_2_argbuf_r,
          isZacQ_4_1_argbuf_r,
          isZacQ_3_2_argbuf_r,
          isZacQ_2_2_argbuf_r,
          \call_main_map'_Bool_Nat_goMux2_r } = (go_7_goMux_choice_1_r ? isZacQ_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty MyDTBool_Nat) : (go_7_goMux_choice_2,C5) [(call_main_map'_Bool_Nat_goMux3,MyDTBool_Nat),
                                                  (gacR_2_2_argbuf,MyDTBool_Nat),
                                                  (gacR_3_2_argbuf,MyDTBool_Nat),
                                                  (gacR_4_1_argbuf,MyDTBool_Nat),
                                                  (lizzieLet6_3QNode_Bool_2_argbuf,MyDTBool_Nat)] > (gacR_goMux_mux,MyDTBool_Nat) */
  logic [0:0] gacR_goMux_mux_mux;
  logic [4:0] gacR_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_2_d[3:1])
      3'd0:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Bool_Nat_goMux3_d };
      3'd1:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd2,
                                                       gacR_2_2_argbuf_d};
      3'd2:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd4,
                                                       gacR_3_2_argbuf_d};
      3'd3:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd8,
                                                       gacR_4_1_argbuf_d};
      3'd4:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd16,
                                                       lizzieLet6_3QNode_Bool_2_argbuf_d};
      default:
        {gacR_goMux_mux_onehot, gacR_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacR_goMux_mux_d = (gacR_goMux_mux_mux[0] && go_7_goMux_choice_2_d[0]);
  assign go_7_goMux_choice_2_r = (gacR_goMux_mux_d[0] && gacR_goMux_mux_r);
  assign {lizzieLet6_3QNode_Bool_2_argbuf_r,
          gacR_4_1_argbuf_r,
          gacR_3_2_argbuf_r,
          gacR_2_2_argbuf_r,
          \call_main_map'_Bool_Nat_goMux3_r } = (go_7_goMux_choice_2_r ? gacR_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_7_goMux_choice_3,C5) [(call_main_map'_Bool_Nat_goMux4,Pointer_QTree_Bool),
                                                        (q3acW_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2acV_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1acU_3_1_argbuf,Pointer_QTree_Bool),
                                                        (q4acX_1_argbuf,Pointer_QTree_Bool)] > (macS_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] macS_goMux_mux_mux;
  logic [4:0] macS_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_3_d[3:1])
      3'd0:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd1,
                                                       \call_main_map'_Bool_Nat_goMux4_d };
      3'd1:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd2,
                                                       q3acW_1_1_argbuf_d};
      3'd2:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd4,
                                                       q2acV_2_1_argbuf_d};
      3'd3:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd8,
                                                       q1acU_3_1_argbuf_d};
      3'd4:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd16,
                                                       q4acX_1_argbuf_d};
      default:
        {macS_goMux_mux_onehot, macS_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign macS_goMux_mux_d = {macS_goMux_mux_mux[16:1],
                             (macS_goMux_mux_mux[0] && go_7_goMux_choice_3_d[0])};
  assign go_7_goMux_choice_3_r = (macS_goMux_mux_d[0] && macS_goMux_mux_r);
  assign {q4acX_1_argbuf_r,
          q1acU_3_1_argbuf_r,
          q2acV_2_1_argbuf_r,
          q3acW_1_1_argbuf_r,
          \call_main_map'_Bool_Nat_goMux4_r } = (go_7_goMux_choice_3_r ? macS_goMux_mux_onehot :
                                                 5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmain_map'_Bool_Nat) : (go_7_goMux_choice_4,C5) [(call_main_map'_Bool_Nat_goMux5,Pointer_CTmain_map'_Bool_Nat),
                                                                  (sca2_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                  (sca1_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                  (sca0_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat),
                                                                  (sca3_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat)] > (sc_0_1_goMux_mux,Pointer_CTmain_map'_Bool_Nat) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_7_goMux_choice_4_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_main_map'_Bool_Nat_goMux5_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_7_goMux_choice_4_d[0])};
  assign go_7_goMux_choice_4_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_main_map'_Bool_Nat_goMux5_r } = (go_7_goMux_choice_4_r ? sc_0_1_goMux_mux_onehot :
                                                 5'd0);
  
  /* fork (Ty C5) : (go_8_goMux_choice,C5) > [(go_8_goMux_choice_1,C5),
                                         (go_8_goMux_choice_2,C5),
                                         (go_8_goMux_choice_3,C5),
                                         (go_8_goMux_choice_4,C5),
                                         (go_8_goMux_choice_5,C5)] */
  logic [4:0] go_8_goMux_choice_emitted;
  logic [4:0] go_8_goMux_choice_done;
  assign go_8_goMux_choice_1_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[0]))};
  assign go_8_goMux_choice_2_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[1]))};
  assign go_8_goMux_choice_3_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[2]))};
  assign go_8_goMux_choice_4_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[3]))};
  assign go_8_goMux_choice_5_d = {go_8_goMux_choice_d[3:1],
                                  (go_8_goMux_choice_d[0] && (! go_8_goMux_choice_emitted[4]))};
  assign go_8_goMux_choice_done = (go_8_goMux_choice_emitted | ({go_8_goMux_choice_5_d[0],
                                                                 go_8_goMux_choice_4_d[0],
                                                                 go_8_goMux_choice_3_d[0],
                                                                 go_8_goMux_choice_2_d[0],
                                                                 go_8_goMux_choice_1_d[0]} & {go_8_goMux_choice_5_r,
                                                                                              go_8_goMux_choice_4_r,
                                                                                              go_8_goMux_choice_3_r,
                                                                                              go_8_goMux_choice_2_r,
                                                                                              go_8_goMux_choice_1_r}));
  assign go_8_goMux_choice_r = (& go_8_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_8_goMux_choice_emitted <= 5'd0;
    else
      go_8_goMux_choice_emitted <= (go_8_goMux_choice_r ? 5'd0 :
                                    go_8_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool) : (go_8_goMux_choice_1,C5) [(call_map''_map''_Bool_Bool_Bool_goMux2,MyDTBool_Bool),
                                                   (isZacY_2_2_argbuf,MyDTBool_Bool),
                                                   (isZacY_3_2_argbuf,MyDTBool_Bool),
                                                   (isZacY_4_1_argbuf,MyDTBool_Bool),
                                                   (lizzieLet12_1_5QNode_Bool_2_argbuf,MyDTBool_Bool)] > (isZacY_goMux_mux,MyDTBool_Bool) */
  logic [0:0] isZacY_goMux_mux_mux;
  logic [4:0] isZacY_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_1_d[3:1])
      3'd0:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Bool_Bool_Bool_goMux2_d };
      3'd1:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd2,
                                                           isZacY_2_2_argbuf_d};
      3'd2:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd4,
                                                           isZacY_3_2_argbuf_d};
      3'd3:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd8,
                                                           isZacY_4_1_argbuf_d};
      3'd4:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd16,
                                                           lizzieLet12_1_5QNode_Bool_2_argbuf_d};
      default:
        {isZacY_goMux_mux_onehot, isZacY_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign isZacY_goMux_mux_d = (isZacY_goMux_mux_mux[0] && go_8_goMux_choice_1_d[0]);
  assign go_8_goMux_choice_1_r = (isZacY_goMux_mux_d[0] && isZacY_goMux_mux_r);
  assign {lizzieLet12_1_5QNode_Bool_2_argbuf_r,
          isZacY_4_1_argbuf_r,
          isZacY_3_2_argbuf_r,
          isZacY_2_2_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux2_r } = (go_8_goMux_choice_1_r ? isZacY_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty MyDTBool_Bool_Bool) : (go_8_goMux_choice_2,C5) [(call_map''_map''_Bool_Bool_Bool_goMux3,MyDTBool_Bool_Bool),
                                                        (gacZ_2_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacZ_3_2_argbuf,MyDTBool_Bool_Bool),
                                                        (gacZ_4_1_argbuf,MyDTBool_Bool_Bool),
                                                        (lizzieLet12_1_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool)] > (gacZ_goMux_mux,MyDTBool_Bool_Bool) */
  logic [0:0] gacZ_goMux_mux_mux;
  logic [4:0] gacZ_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_2_d[3:1])
      3'd0:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Bool_Bool_Bool_goMux3_d };
      3'd1:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd2,
                                                       gacZ_2_2_argbuf_d};
      3'd2:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd4,
                                                       gacZ_3_2_argbuf_d};
      3'd3:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd8,
                                                       gacZ_4_1_argbuf_d};
      3'd4:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd16,
                                                       lizzieLet12_1_3QNode_Bool_2_argbuf_d};
      default:
        {gacZ_goMux_mux_onehot, gacZ_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign gacZ_goMux_mux_d = (gacZ_goMux_mux_mux[0] && go_8_goMux_choice_2_d[0]);
  assign go_8_goMux_choice_2_r = (gacZ_goMux_mux_d[0] && gacZ_goMux_mux_r);
  assign {lizzieLet12_1_3QNode_Bool_2_argbuf_r,
          gacZ_4_1_argbuf_r,
          gacZ_3_2_argbuf_r,
          gacZ_2_2_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux3_r } = (go_8_goMux_choice_2_r ? gacZ_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty MyBool) : (go_8_goMux_choice_3,C5) [(call_map''_map''_Bool_Bool_Bool_goMux4,MyBool),
                                            (v'ad0_2_2_argbuf,MyBool),
                                            (v'ad0_3_2_argbuf,MyBool),
                                            (v'ad0_4_1_argbuf,MyBool),
                                            (lizzieLet12_1_7QNode_Bool_2_argbuf,MyBool)] > (v'ad0_goMux_mux,MyBool) */
  logic [1:0] \v'ad0_goMux_mux_mux ;
  logic [4:0] \v'ad0_goMux_mux_onehot ;
  always_comb
    unique case (go_8_goMux_choice_3_d[3:1])
      3'd0:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd1,
                                                             \call_map''_map''_Bool_Bool_Bool_goMux4_d };
      3'd1:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd2,
                                                             \v'ad0_2_2_argbuf_d };
      3'd2:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd4,
                                                             \v'ad0_3_2_argbuf_d };
      3'd3:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd8,
                                                             \v'ad0_4_1_argbuf_d };
      3'd4:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd16,
                                                             lizzieLet12_1_7QNode_Bool_2_argbuf_d};
      default:
        {\v'ad0_goMux_mux_onehot , \v'ad0_goMux_mux_mux } = {5'd0,
                                                             {1'd0, 1'd0}};
    endcase
  assign \v'ad0_goMux_mux_d  = {\v'ad0_goMux_mux_mux [1:1],
                                (\v'ad0_goMux_mux_mux [0] && go_8_goMux_choice_3_d[0])};
  assign go_8_goMux_choice_3_r = (\v'ad0_goMux_mux_d [0] && \v'ad0_goMux_mux_r );
  assign {lizzieLet12_1_7QNode_Bool_2_argbuf_r,
          \v'ad0_4_1_argbuf_r ,
          \v'ad0_3_2_argbuf_r ,
          \v'ad0_2_2_argbuf_r ,
          \call_map''_map''_Bool_Bool_Bool_goMux4_r } = (go_8_goMux_choice_3_r ? \v'ad0_goMux_mux_onehot  :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Bool) : (go_8_goMux_choice_4,C5) [(call_map''_map''_Bool_Bool_Bool_goMux5,Pointer_QTree_Bool),
                                                        (q3ad5_1_1_argbuf,Pointer_QTree_Bool),
                                                        (q2ad4_2_1_argbuf,Pointer_QTree_Bool),
                                                        (q1ad3_3_1_argbuf,Pointer_QTree_Bool),
                                                        (q4ad6_1_argbuf,Pointer_QTree_Bool)] > (mad1_goMux_mux,Pointer_QTree_Bool) */
  logic [16:0] mad1_goMux_mux_mux;
  logic [4:0] mad1_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_4_d[3:1])
      3'd0:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd1,
                                                       \call_map''_map''_Bool_Bool_Bool_goMux5_d };
      3'd1:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd2,
                                                       q3ad5_1_1_argbuf_d};
      3'd2:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd4,
                                                       q2ad4_2_1_argbuf_d};
      3'd3:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd8,
                                                       q1ad3_3_1_argbuf_d};
      3'd4:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd16,
                                                       q4ad6_1_argbuf_d};
      default:
        {mad1_goMux_mux_onehot, mad1_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign mad1_goMux_mux_d = {mad1_goMux_mux_mux[16:1],
                             (mad1_goMux_mux_mux[0] && go_8_goMux_choice_4_d[0])};
  assign go_8_goMux_choice_4_r = (mad1_goMux_mux_d[0] && mad1_goMux_mux_r);
  assign {q4ad6_1_argbuf_r,
          q1ad3_3_1_argbuf_r,
          q2ad4_2_1_argbuf_r,
          q3ad5_1_1_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux5_r } = (go_8_goMux_choice_4_r ? mad1_goMux_mux_onehot :
                                                         5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (go_8_goMux_choice_5,C5) [(call_map''_map''_Bool_Bool_Bool_goMux6,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca2_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca1_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                          (sca3_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (sc_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_8_goMux_choice_5_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           \call_map''_map''_Bool_Bool_Bool_goMux6_d };
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_8_goMux_choice_5_d[0])};
  assign go_8_goMux_choice_5_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          \call_map''_map''_Bool_Bool_Bool_goMux6_r } = (go_8_goMux_choice_5_r ? sc_0_2_goMux_mux_onehot :
                                                         5'd0);
  
  /* fork (Ty C2) : (go_9_goMux_choice,C2) > [(go_9_goMux_choice_1,C2),
                                         (go_9_goMux_choice_2,C2)] */
  logic [1:0] go_9_goMux_choice_emitted;
  logic [1:0] go_9_goMux_choice_done;
  assign go_9_goMux_choice_1_d = {go_9_goMux_choice_d[1:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[0]))};
  assign go_9_goMux_choice_2_d = {go_9_goMux_choice_d[1:1],
                                  (go_9_goMux_choice_d[0] && (! go_9_goMux_choice_emitted[1]))};
  assign go_9_goMux_choice_done = (go_9_goMux_choice_emitted | ({go_9_goMux_choice_2_d[0],
                                                                 go_9_goMux_choice_1_d[0]} & {go_9_goMux_choice_2_r,
                                                                                              go_9_goMux_choice_1_r}));
  assign go_9_goMux_choice_r = (& go_9_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_9_goMux_choice_emitted <= 2'd0;
    else
      go_9_goMux_choice_emitted <= (go_9_goMux_choice_r ? 2'd0 :
                                    go_9_goMux_choice_done);
  
  /* mux (Ty C2,
     Ty Pointer_Nat) : (go_9_goMux_choice_1,C2) [(eqNat_goMux2,Pointer_Nat),
                                                 (lizzieLet18_4Succ_4Succ_1_argbuf,Pointer_Nat)] > (xadg_goMux_mux,Pointer_Nat) */
  logic [16:0] xadg_goMux_mux_mux;
  logic [1:0] xadg_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_1_d[1:1])
      1'd0:
        {xadg_goMux_mux_onehot, xadg_goMux_mux_mux} = {2'd1,
                                                       eqNat_goMux2_d};
      1'd1:
        {xadg_goMux_mux_onehot, xadg_goMux_mux_mux} = {2'd2,
                                                       lizzieLet18_4Succ_4Succ_1_argbuf_d};
      default:
        {xadg_goMux_mux_onehot, xadg_goMux_mux_mux} = {2'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign xadg_goMux_mux_d = {xadg_goMux_mux_mux[16:1],
                             (xadg_goMux_mux_mux[0] && go_9_goMux_choice_1_d[0])};
  assign go_9_goMux_choice_1_r = (xadg_goMux_mux_d[0] && xadg_goMux_mux_r);
  assign {lizzieLet18_4Succ_4Succ_1_argbuf_r,
          eqNat_goMux2_r} = (go_9_goMux_choice_1_r ? xadg_goMux_mux_onehot :
                             2'd0);
  
  /* mux (Ty C2,
     Ty Pointer_Nat) : (go_9_goMux_choice_2,C2) [(eqNat_goMux3,Pointer_Nat),
                                                 (y1adk_1_argbuf,Pointer_Nat)] > (yadh_goMux_mux,Pointer_Nat) */
  logic [16:0] yadh_goMux_mux_mux;
  logic [1:0] yadh_goMux_mux_onehot;
  always_comb
    unique case (go_9_goMux_choice_2_d[1:1])
      1'd0:
        {yadh_goMux_mux_onehot, yadh_goMux_mux_mux} = {2'd1,
                                                       eqNat_goMux3_d};
      1'd1:
        {yadh_goMux_mux_onehot, yadh_goMux_mux_mux} = {2'd2,
                                                       y1adk_1_argbuf_d};
      default:
        {yadh_goMux_mux_onehot, yadh_goMux_mux_mux} = {2'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign yadh_goMux_mux_d = {yadh_goMux_mux_mux[16:1],
                             (yadh_goMux_mux_mux[0] && go_9_goMux_choice_2_d[0])};
  assign go_9_goMux_choice_2_r = (yadh_goMux_mux_d[0] && yadh_goMux_mux_r);
  assign {y1adk_1_argbuf_r,
          eqNat_goMux3_r} = (go_9_goMux_choice_2_r ? yadh_goMux_mux_onehot :
                             2'd0);
  
  /* buf (Ty MyDTNat_Bool) : (isZacQ_2_2,MyDTNat_Bool) > (isZacQ_2_2_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t isZacQ_2_2_bufchan_d;
  logic isZacQ_2_2_bufchan_r;
  assign isZacQ_2_2_r = ((! isZacQ_2_2_bufchan_d[0]) || isZacQ_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_2_2_bufchan_d <= 1'd0;
    else if (isZacQ_2_2_r) isZacQ_2_2_bufchan_d <= isZacQ_2_2_d;
  MyDTNat_Bool_t isZacQ_2_2_bufchan_buf;
  assign isZacQ_2_2_bufchan_r = (! isZacQ_2_2_bufchan_buf[0]);
  assign isZacQ_2_2_argbuf_d = (isZacQ_2_2_bufchan_buf[0] ? isZacQ_2_2_bufchan_buf :
                                isZacQ_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacQ_2_2_argbuf_r && isZacQ_2_2_bufchan_buf[0]))
        isZacQ_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacQ_2_2_argbuf_r) && (! isZacQ_2_2_bufchan_buf[0])))
        isZacQ_2_2_bufchan_buf <= isZacQ_2_2_bufchan_d;
  
  /* fork (Ty MyDTNat_Bool) : (isZacQ_2_destruct,MyDTNat_Bool) > [(isZacQ_2_1,MyDTNat_Bool),
                                                             (isZacQ_2_2,MyDTNat_Bool)] */
  logic [1:0] isZacQ_2_destruct_emitted;
  logic [1:0] isZacQ_2_destruct_done;
  assign isZacQ_2_1_d = (isZacQ_2_destruct_d[0] && (! isZacQ_2_destruct_emitted[0]));
  assign isZacQ_2_2_d = (isZacQ_2_destruct_d[0] && (! isZacQ_2_destruct_emitted[1]));
  assign isZacQ_2_destruct_done = (isZacQ_2_destruct_emitted | ({isZacQ_2_2_d[0],
                                                                 isZacQ_2_1_d[0]} & {isZacQ_2_2_r,
                                                                                     isZacQ_2_1_r}));
  assign isZacQ_2_destruct_r = (& isZacQ_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_2_destruct_emitted <= 2'd0;
    else
      isZacQ_2_destruct_emitted <= (isZacQ_2_destruct_r ? 2'd0 :
                                    isZacQ_2_destruct_done);
  
  /* buf (Ty MyDTNat_Bool) : (isZacQ_3_2,MyDTNat_Bool) > (isZacQ_3_2_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t isZacQ_3_2_bufchan_d;
  logic isZacQ_3_2_bufchan_r;
  assign isZacQ_3_2_r = ((! isZacQ_3_2_bufchan_d[0]) || isZacQ_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_3_2_bufchan_d <= 1'd0;
    else if (isZacQ_3_2_r) isZacQ_3_2_bufchan_d <= isZacQ_3_2_d;
  MyDTNat_Bool_t isZacQ_3_2_bufchan_buf;
  assign isZacQ_3_2_bufchan_r = (! isZacQ_3_2_bufchan_buf[0]);
  assign isZacQ_3_2_argbuf_d = (isZacQ_3_2_bufchan_buf[0] ? isZacQ_3_2_bufchan_buf :
                                isZacQ_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacQ_3_2_argbuf_r && isZacQ_3_2_bufchan_buf[0]))
        isZacQ_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacQ_3_2_argbuf_r) && (! isZacQ_3_2_bufchan_buf[0])))
        isZacQ_3_2_bufchan_buf <= isZacQ_3_2_bufchan_d;
  
  /* fork (Ty MyDTNat_Bool) : (isZacQ_3_destruct,MyDTNat_Bool) > [(isZacQ_3_1,MyDTNat_Bool),
                                                             (isZacQ_3_2,MyDTNat_Bool)] */
  logic [1:0] isZacQ_3_destruct_emitted;
  logic [1:0] isZacQ_3_destruct_done;
  assign isZacQ_3_1_d = (isZacQ_3_destruct_d[0] && (! isZacQ_3_destruct_emitted[0]));
  assign isZacQ_3_2_d = (isZacQ_3_destruct_d[0] && (! isZacQ_3_destruct_emitted[1]));
  assign isZacQ_3_destruct_done = (isZacQ_3_destruct_emitted | ({isZacQ_3_2_d[0],
                                                                 isZacQ_3_1_d[0]} & {isZacQ_3_2_r,
                                                                                     isZacQ_3_1_r}));
  assign isZacQ_3_destruct_r = (& isZacQ_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_3_destruct_emitted <= 2'd0;
    else
      isZacQ_3_destruct_emitted <= (isZacQ_3_destruct_r ? 2'd0 :
                                    isZacQ_3_destruct_done);
  
  /* buf (Ty MyDTNat_Bool) : (isZacQ_4_destruct,MyDTNat_Bool) > (isZacQ_4_1_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t isZacQ_4_destruct_bufchan_d;
  logic isZacQ_4_destruct_bufchan_r;
  assign isZacQ_4_destruct_r = ((! isZacQ_4_destruct_bufchan_d[0]) || isZacQ_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacQ_4_destruct_r)
        isZacQ_4_destruct_bufchan_d <= isZacQ_4_destruct_d;
  MyDTNat_Bool_t isZacQ_4_destruct_bufchan_buf;
  assign isZacQ_4_destruct_bufchan_r = (! isZacQ_4_destruct_bufchan_buf[0]);
  assign isZacQ_4_1_argbuf_d = (isZacQ_4_destruct_bufchan_buf[0] ? isZacQ_4_destruct_bufchan_buf :
                                isZacQ_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacQ_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacQ_4_1_argbuf_r && isZacQ_4_destruct_bufchan_buf[0]))
        isZacQ_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacQ_4_1_argbuf_r) && (! isZacQ_4_destruct_bufchan_buf[0])))
        isZacQ_4_destruct_bufchan_buf <= isZacQ_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (isZacY_2_2,MyDTBool_Bool) > (isZacY_2_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacY_2_2_bufchan_d;
  logic isZacY_2_2_bufchan_r;
  assign isZacY_2_2_r = ((! isZacY_2_2_bufchan_d[0]) || isZacY_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_2_2_bufchan_d <= 1'd0;
    else if (isZacY_2_2_r) isZacY_2_2_bufchan_d <= isZacY_2_2_d;
  MyDTBool_Bool_t isZacY_2_2_bufchan_buf;
  assign isZacY_2_2_bufchan_r = (! isZacY_2_2_bufchan_buf[0]);
  assign isZacY_2_2_argbuf_d = (isZacY_2_2_bufchan_buf[0] ? isZacY_2_2_bufchan_buf :
                                isZacY_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZacY_2_2_argbuf_r && isZacY_2_2_bufchan_buf[0]))
        isZacY_2_2_bufchan_buf <= 1'd0;
      else if (((! isZacY_2_2_argbuf_r) && (! isZacY_2_2_bufchan_buf[0])))
        isZacY_2_2_bufchan_buf <= isZacY_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacY_2_destruct,MyDTBool_Bool) > [(isZacY_2_1,MyDTBool_Bool),
                                                               (isZacY_2_2,MyDTBool_Bool)] */
  logic [1:0] isZacY_2_destruct_emitted;
  logic [1:0] isZacY_2_destruct_done;
  assign isZacY_2_1_d = (isZacY_2_destruct_d[0] && (! isZacY_2_destruct_emitted[0]));
  assign isZacY_2_2_d = (isZacY_2_destruct_d[0] && (! isZacY_2_destruct_emitted[1]));
  assign isZacY_2_destruct_done = (isZacY_2_destruct_emitted | ({isZacY_2_2_d[0],
                                                                 isZacY_2_1_d[0]} & {isZacY_2_2_r,
                                                                                     isZacY_2_1_r}));
  assign isZacY_2_destruct_r = (& isZacY_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_2_destruct_emitted <= 2'd0;
    else
      isZacY_2_destruct_emitted <= (isZacY_2_destruct_r ? 2'd0 :
                                    isZacY_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacY_3_2,MyDTBool_Bool) > (isZacY_3_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacY_3_2_bufchan_d;
  logic isZacY_3_2_bufchan_r;
  assign isZacY_3_2_r = ((! isZacY_3_2_bufchan_d[0]) || isZacY_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_3_2_bufchan_d <= 1'd0;
    else if (isZacY_3_2_r) isZacY_3_2_bufchan_d <= isZacY_3_2_d;
  MyDTBool_Bool_t isZacY_3_2_bufchan_buf;
  assign isZacY_3_2_bufchan_r = (! isZacY_3_2_bufchan_buf[0]);
  assign isZacY_3_2_argbuf_d = (isZacY_3_2_bufchan_buf[0] ? isZacY_3_2_bufchan_buf :
                                isZacY_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZacY_3_2_argbuf_r && isZacY_3_2_bufchan_buf[0]))
        isZacY_3_2_bufchan_buf <= 1'd0;
      else if (((! isZacY_3_2_argbuf_r) && (! isZacY_3_2_bufchan_buf[0])))
        isZacY_3_2_bufchan_buf <= isZacY_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZacY_3_destruct,MyDTBool_Bool) > [(isZacY_3_1,MyDTBool_Bool),
                                                               (isZacY_3_2,MyDTBool_Bool)] */
  logic [1:0] isZacY_3_destruct_emitted;
  logic [1:0] isZacY_3_destruct_done;
  assign isZacY_3_1_d = (isZacY_3_destruct_d[0] && (! isZacY_3_destruct_emitted[0]));
  assign isZacY_3_2_d = (isZacY_3_destruct_d[0] && (! isZacY_3_destruct_emitted[1]));
  assign isZacY_3_destruct_done = (isZacY_3_destruct_emitted | ({isZacY_3_2_d[0],
                                                                 isZacY_3_1_d[0]} & {isZacY_3_2_r,
                                                                                     isZacY_3_1_r}));
  assign isZacY_3_destruct_r = (& isZacY_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_3_destruct_emitted <= 2'd0;
    else
      isZacY_3_destruct_emitted <= (isZacY_3_destruct_r ? 2'd0 :
                                    isZacY_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZacY_4_destruct,MyDTBool_Bool) > (isZacY_4_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZacY_4_destruct_bufchan_d;
  logic isZacY_4_destruct_bufchan_r;
  assign isZacY_4_destruct_r = ((! isZacY_4_destruct_bufchan_d[0]) || isZacY_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZacY_4_destruct_r)
        isZacY_4_destruct_bufchan_d <= isZacY_4_destruct_d;
  MyDTBool_Bool_t isZacY_4_destruct_bufchan_buf;
  assign isZacY_4_destruct_bufchan_r = (! isZacY_4_destruct_bufchan_buf[0]);
  assign isZacY_4_1_argbuf_d = (isZacY_4_destruct_bufchan_buf[0] ? isZacY_4_destruct_bufchan_buf :
                                isZacY_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZacY_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZacY_4_1_argbuf_r && isZacY_4_destruct_bufchan_buf[0]))
        isZacY_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZacY_4_1_argbuf_r) && (! isZacY_4_destruct_bufchan_buf[0])))
        isZacY_4_destruct_bufchan_buf <= isZacY_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (isZad7_2_2,MyDTBool_Bool) > (isZad7_2_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZad7_2_2_bufchan_d;
  logic isZad7_2_2_bufchan_r;
  assign isZad7_2_2_r = ((! isZad7_2_2_bufchan_d[0]) || isZad7_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_2_2_bufchan_d <= 1'd0;
    else if (isZad7_2_2_r) isZad7_2_2_bufchan_d <= isZad7_2_2_d;
  MyDTBool_Bool_t isZad7_2_2_bufchan_buf;
  assign isZad7_2_2_bufchan_r = (! isZad7_2_2_bufchan_buf[0]);
  assign isZad7_2_2_argbuf_d = (isZad7_2_2_bufchan_buf[0] ? isZad7_2_2_bufchan_buf :
                                isZad7_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_2_2_bufchan_buf <= 1'd0;
    else
      if ((isZad7_2_2_argbuf_r && isZad7_2_2_bufchan_buf[0]))
        isZad7_2_2_bufchan_buf <= 1'd0;
      else if (((! isZad7_2_2_argbuf_r) && (! isZad7_2_2_bufchan_buf[0])))
        isZad7_2_2_bufchan_buf <= isZad7_2_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZad7_2_destruct,MyDTBool_Bool) > [(isZad7_2_1,MyDTBool_Bool),
                                                               (isZad7_2_2,MyDTBool_Bool)] */
  logic [1:0] isZad7_2_destruct_emitted;
  logic [1:0] isZad7_2_destruct_done;
  assign isZad7_2_1_d = (isZad7_2_destruct_d[0] && (! isZad7_2_destruct_emitted[0]));
  assign isZad7_2_2_d = (isZad7_2_destruct_d[0] && (! isZad7_2_destruct_emitted[1]));
  assign isZad7_2_destruct_done = (isZad7_2_destruct_emitted | ({isZad7_2_2_d[0],
                                                                 isZad7_2_1_d[0]} & {isZad7_2_2_r,
                                                                                     isZad7_2_1_r}));
  assign isZad7_2_destruct_r = (& isZad7_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_2_destruct_emitted <= 2'd0;
    else
      isZad7_2_destruct_emitted <= (isZad7_2_destruct_r ? 2'd0 :
                                    isZad7_2_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZad7_3_2,MyDTBool_Bool) > (isZad7_3_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZad7_3_2_bufchan_d;
  logic isZad7_3_2_bufchan_r;
  assign isZad7_3_2_r = ((! isZad7_3_2_bufchan_d[0]) || isZad7_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_3_2_bufchan_d <= 1'd0;
    else if (isZad7_3_2_r) isZad7_3_2_bufchan_d <= isZad7_3_2_d;
  MyDTBool_Bool_t isZad7_3_2_bufchan_buf;
  assign isZad7_3_2_bufchan_r = (! isZad7_3_2_bufchan_buf[0]);
  assign isZad7_3_2_argbuf_d = (isZad7_3_2_bufchan_buf[0] ? isZad7_3_2_bufchan_buf :
                                isZad7_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_3_2_bufchan_buf <= 1'd0;
    else
      if ((isZad7_3_2_argbuf_r && isZad7_3_2_bufchan_buf[0]))
        isZad7_3_2_bufchan_buf <= 1'd0;
      else if (((! isZad7_3_2_argbuf_r) && (! isZad7_3_2_bufchan_buf[0])))
        isZad7_3_2_bufchan_buf <= isZad7_3_2_bufchan_d;
  
  /* fork (Ty MyDTBool_Bool) : (isZad7_3_destruct,MyDTBool_Bool) > [(isZad7_3_1,MyDTBool_Bool),
                                                               (isZad7_3_2,MyDTBool_Bool)] */
  logic [1:0] isZad7_3_destruct_emitted;
  logic [1:0] isZad7_3_destruct_done;
  assign isZad7_3_1_d = (isZad7_3_destruct_d[0] && (! isZad7_3_destruct_emitted[0]));
  assign isZad7_3_2_d = (isZad7_3_destruct_d[0] && (! isZad7_3_destruct_emitted[1]));
  assign isZad7_3_destruct_done = (isZad7_3_destruct_emitted | ({isZad7_3_2_d[0],
                                                                 isZad7_3_1_d[0]} & {isZad7_3_2_r,
                                                                                     isZad7_3_1_r}));
  assign isZad7_3_destruct_r = (& isZad7_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_3_destruct_emitted <= 2'd0;
    else
      isZad7_3_destruct_emitted <= (isZad7_3_destruct_r ? 2'd0 :
                                    isZad7_3_destruct_done);
  
  /* buf (Ty MyDTBool_Bool) : (isZad7_4_destruct,MyDTBool_Bool) > (isZad7_4_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t isZad7_4_destruct_bufchan_d;
  logic isZad7_4_destruct_bufchan_r;
  assign isZad7_4_destruct_r = ((! isZad7_4_destruct_bufchan_d[0]) || isZad7_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_4_destruct_bufchan_d <= 1'd0;
    else
      if (isZad7_4_destruct_r)
        isZad7_4_destruct_bufchan_d <= isZad7_4_destruct_d;
  MyDTBool_Bool_t isZad7_4_destruct_bufchan_buf;
  assign isZad7_4_destruct_bufchan_r = (! isZad7_4_destruct_bufchan_buf[0]);
  assign isZad7_4_1_argbuf_d = (isZad7_4_destruct_bufchan_buf[0] ? isZad7_4_destruct_bufchan_buf :
                                isZad7_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) isZad7_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((isZad7_4_1_argbuf_r && isZad7_4_destruct_bufchan_buf[0]))
        isZad7_4_destruct_bufchan_buf <= 1'd0;
      else if (((! isZad7_4_1_argbuf_r) && (! isZad7_4_destruct_bufchan_buf[0])))
        isZad7_4_destruct_bufchan_buf <= isZad7_4_destruct_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool) > [(kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10,Go),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1,MyDTBool_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1,Pointer_QTree_Bool),
                                                                                                                                                                                                                                                                                                                (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1,Pointer_QTree_Bool)] */
  logic [4:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted;
  logic [4:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[0]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[1]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[2]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_d = {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[16:1],
                                                                                                                                  (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[3]))};
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_d = {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[32:17],
                                                                                                                                  (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted[4]))};
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted | ({kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_d[0],
                                                                                                                                                                                                                                                           kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_d[0]} & {kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_r,
                                                                                                                                                                                                                                                                                                                                                                                      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_r,
                                                                                                                                                                                                                                                                                                                                                                                      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_r,
                                                                                                                                                                                                                                                                                                                                                                                      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_r,
                                                                                                                                                                                                                                                                                                                                                                                      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_r}));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r = (& kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= 5'd0;
    else
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_emitted <= (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_r ? 5'd0 :
                                                                                                                                 kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Bool_1_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1,MyDTBool_Bool_Bool) > (gad8_1_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_d;
  MyDTBool_Bool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf[0]);
  assign gad8_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf :
                              kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf <= 1'd0;
    else
      if ((gad8_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf <= 1'd0;
      else if (((! gad8_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgad8_1_bufchan_d;
  
  /* fork (Ty Go) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10,Go) > [(go_10_1,Go),
                                                                                                                                         (go_10_2,Go)] */
  logic [1:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted;
  logic [1:0] kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_done;
  assign go_10_1_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted[0]));
  assign go_10_2_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_d[0] && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted[1]));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_done = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted | ({go_10_2_d[0],
                                                                                                                                                                                                                                                                 go_10_1_d[0]} & {go_10_2_r,
                                                                                                                                                                                                                                                                                  go_10_1_r}));
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_r = (& kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted <= 2'd0;
    else
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_emitted <= (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_r ? 2'd0 :
                                                                                                                                    kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolgo_10_done);
  
  /* buf (Ty MyDTBool_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1,MyDTBool_Bool) > (isZad7_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d <= 1'd0;
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_d;
  MyDTBool_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf[0]);
  assign isZad7_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf :
                                kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf <= 1'd0;
    else
      if ((isZad7_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf <= 1'd0;
      else if (((! isZad7_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_BoolisZad7_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1,Pointer_QTree_Bool) > (m1ad9_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d <= {16'd0,
                                                                                                                                        1'd0};
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf[0]);
  assign m1ad9_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf :
                               kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf <= {16'd0,
                                                                                                                                          1'd0};
    else
      if ((m1ad9_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf <= {16'd0,
                                                                                                                                            1'd0};
      else if (((! m1ad9_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm1ad9_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1,Pointer_QTree_Bool) > (m2ada_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d;
  logic kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_r;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_r = ((! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d[0]) || kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d <= {16'd0,
                                                                                                                                        1'd0};
    else
      if (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_r)
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf;
  assign kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_r = (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf[0]);
  assign m2ada_1_1_argbuf_d = (kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf[0] ? kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf :
                               kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf <= {16'd0,
                                                                                                                                          1'd0};
    else
      if ((m2ada_1_1_argbuf_r && kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf[0]))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf <= {16'd0,
                                                                                                                                            1'd0};
      else if (((! m2ada_1_1_argbuf_r) && (! kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf[0])))
        kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_buf <= kron_kron_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___Pointer_QTree_Bool___Pointer_QTree_Boolm2ada_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (kron_kron_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) > (es_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_bufchan_d;
  logic kron_kron_Bool_Bool_Bool_resbuf_bufchan_r;
  assign kron_kron_Bool_Bool_Bool_resbuf_r = ((! kron_kron_Bool_Bool_Bool_resbuf_bufchan_d[0]) || kron_kron_Bool_Bool_Bool_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_Bool_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (kron_kron_Bool_Bool_Bool_resbuf_r)
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_d <= kron_kron_Bool_Bool_Bool_resbuf_d;
  Pointer_QTree_Bool_t kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf;
  assign kron_kron_Bool_Bool_Bool_resbuf_bufchan_r = (! kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0]);
  assign es_2_1_argbuf_d = (kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0] ? kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf :
                            kron_kron_Bool_Bool_Bool_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_1_argbuf_r && kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0]))
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_1_argbuf_r) && (! kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf[0])))
        kron_kron_Bool_Bool_Bool_resbuf_bufchan_buf <= kron_kron_Bool_Bool_Bool_resbuf_bufchan_d;
  
  /* buf (Ty Nat) : (lizzieLet0_1_1Succ,Nat) > (lizzieLet40_1_argbuf,Nat) */
  Nat_t lizzieLet0_1_1Succ_bufchan_d;
  logic lizzieLet0_1_1Succ_bufchan_r;
  assign lizzieLet0_1_1Succ_r = ((! lizzieLet0_1_1Succ_bufchan_d[0]) || lizzieLet0_1_1Succ_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_1Succ_bufchan_d <= {17'd0, 1'd0};
    else
      if (lizzieLet0_1_1Succ_r)
        lizzieLet0_1_1Succ_bufchan_d <= lizzieLet0_1_1Succ_d;
  Nat_t lizzieLet0_1_1Succ_bufchan_buf;
  assign lizzieLet0_1_1Succ_bufchan_r = (! lizzieLet0_1_1Succ_bufchan_buf[0]);
  assign lizzieLet40_1_argbuf_d = (lizzieLet0_1_1Succ_bufchan_buf[0] ? lizzieLet0_1_1Succ_bufchan_buf :
                                   lizzieLet0_1_1Succ_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet0_1_1Succ_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((lizzieLet40_1_argbuf_r && lizzieLet0_1_1Succ_bufchan_buf[0]))
        lizzieLet0_1_1Succ_bufchan_buf <= {17'd0, 1'd0};
      else if (((! lizzieLet40_1_argbuf_r) && (! lizzieLet0_1_1Succ_bufchan_buf[0])))
        lizzieLet0_1_1Succ_bufchan_buf <= lizzieLet0_1_1Succ_bufchan_d;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet12_1_1QNode_Bool,QTree_Bool) > [(q1ad3_destruct,Pointer_QTree_Bool),
                                                                       (q2ad4_destruct,Pointer_QTree_Bool),
                                                                       (q3ad5_destruct,Pointer_QTree_Bool),
                                                                       (q4ad6_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet12_1_1QNode_Bool_emitted;
  logic [3:0] lizzieLet12_1_1QNode_Bool_done;
  assign q1ad3_destruct_d = {lizzieLet12_1_1QNode_Bool_d[18:3],
                             (lizzieLet12_1_1QNode_Bool_d[0] && (! lizzieLet12_1_1QNode_Bool_emitted[0]))};
  assign q2ad4_destruct_d = {lizzieLet12_1_1QNode_Bool_d[34:19],
                             (lizzieLet12_1_1QNode_Bool_d[0] && (! lizzieLet12_1_1QNode_Bool_emitted[1]))};
  assign q3ad5_destruct_d = {lizzieLet12_1_1QNode_Bool_d[50:35],
                             (lizzieLet12_1_1QNode_Bool_d[0] && (! lizzieLet12_1_1QNode_Bool_emitted[2]))};
  assign q4ad6_destruct_d = {lizzieLet12_1_1QNode_Bool_d[66:51],
                             (lizzieLet12_1_1QNode_Bool_d[0] && (! lizzieLet12_1_1QNode_Bool_emitted[3]))};
  assign lizzieLet12_1_1QNode_Bool_done = (lizzieLet12_1_1QNode_Bool_emitted | ({q4ad6_destruct_d[0],
                                                                                 q3ad5_destruct_d[0],
                                                                                 q2ad4_destruct_d[0],
                                                                                 q1ad3_destruct_d[0]} & {q4ad6_destruct_r,
                                                                                                         q3ad5_destruct_r,
                                                                                                         q2ad4_destruct_r,
                                                                                                         q1ad3_destruct_r}));
  assign lizzieLet12_1_1QNode_Bool_r = (& lizzieLet12_1_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet12_1_1QNode_Bool_emitted <= (lizzieLet12_1_1QNode_Bool_r ? 4'd0 :
                                            lizzieLet12_1_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet12_1_1QVal_Bool,QTree_Bool) > [(vad2_destruct,MyBool)] */
  assign vad2_destruct_d = {lizzieLet12_1_1QVal_Bool_d[3:3],
                            lizzieLet12_1_1QVal_Bool_d[0]};
  assign lizzieLet12_1_1QVal_Bool_r = vad2_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet12_1_2,QTree_Bool) (lizzieLet12_1_1,QTree_Bool) > [(_30,QTree_Bool),
                                                                                     (lizzieLet12_1_1QVal_Bool,QTree_Bool),
                                                                                     (lizzieLet12_1_1QNode_Bool,QTree_Bool),
                                                                                     (_29,QTree_Bool)] */
  logic [3:0] lizzieLet12_1_1_onehotd;
  always_comb
    if ((lizzieLet12_1_2_d[0] && lizzieLet12_1_1_d[0]))
      unique case (lizzieLet12_1_2_d[2:1])
        2'd0: lizzieLet12_1_1_onehotd = 4'd1;
        2'd1: lizzieLet12_1_1_onehotd = 4'd2;
        2'd2: lizzieLet12_1_1_onehotd = 4'd4;
        2'd3: lizzieLet12_1_1_onehotd = 4'd8;
        default: lizzieLet12_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet12_1_1_onehotd = 4'd0;
  assign _30_d = {lizzieLet12_1_1_d[66:1],
                  lizzieLet12_1_1_onehotd[0]};
  assign lizzieLet12_1_1QVal_Bool_d = {lizzieLet12_1_1_d[66:1],
                                       lizzieLet12_1_1_onehotd[1]};
  assign lizzieLet12_1_1QNode_Bool_d = {lizzieLet12_1_1_d[66:1],
                                        lizzieLet12_1_1_onehotd[2]};
  assign _29_d = {lizzieLet12_1_1_d[66:1],
                  lizzieLet12_1_1_onehotd[3]};
  assign lizzieLet12_1_1_r = (| (lizzieLet12_1_1_onehotd & {_29_r,
                                                            lizzieLet12_1_1QNode_Bool_r,
                                                            lizzieLet12_1_1QVal_Bool_r,
                                                            _30_r}));
  assign lizzieLet12_1_2_r = lizzieLet12_1_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet12_1_3,QTree_Bool) (gacZ_goMux_mux,MyDTBool_Bool_Bool) > [(_28,MyDTBool_Bool_Bool),
                                                                                                    (lizzieLet12_1_3QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                    (lizzieLet12_1_3QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                    (_27,MyDTBool_Bool_Bool)] */
  logic [3:0] gacZ_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_1_3_d[0] && gacZ_goMux_mux_d[0]))
      unique case (lizzieLet12_1_3_d[2:1])
        2'd0: gacZ_goMux_mux_onehotd = 4'd1;
        2'd1: gacZ_goMux_mux_onehotd = 4'd2;
        2'd2: gacZ_goMux_mux_onehotd = 4'd4;
        2'd3: gacZ_goMux_mux_onehotd = 4'd8;
        default: gacZ_goMux_mux_onehotd = 4'd0;
      endcase
    else gacZ_goMux_mux_onehotd = 4'd0;
  assign _28_d = gacZ_goMux_mux_onehotd[0];
  assign lizzieLet12_1_3QVal_Bool_d = gacZ_goMux_mux_onehotd[1];
  assign lizzieLet12_1_3QNode_Bool_d = gacZ_goMux_mux_onehotd[2];
  assign _27_d = gacZ_goMux_mux_onehotd[3];
  assign gacZ_goMux_mux_r = (| (gacZ_goMux_mux_onehotd & {_27_r,
                                                          lizzieLet12_1_3QNode_Bool_r,
                                                          lizzieLet12_1_3QVal_Bool_r,
                                                          _28_r}));
  assign lizzieLet12_1_3_r = gacZ_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (lizzieLet12_1_3QNode_Bool,MyDTBool_Bool_Bool) > [(lizzieLet12_1_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                                                 (lizzieLet12_1_3QNode_Bool_2,MyDTBool_Bool_Bool)] */
  logic [1:0] lizzieLet12_1_3QNode_Bool_emitted;
  logic [1:0] lizzieLet12_1_3QNode_Bool_done;
  assign lizzieLet12_1_3QNode_Bool_1_d = (lizzieLet12_1_3QNode_Bool_d[0] && (! lizzieLet12_1_3QNode_Bool_emitted[0]));
  assign lizzieLet12_1_3QNode_Bool_2_d = (lizzieLet12_1_3QNode_Bool_d[0] && (! lizzieLet12_1_3QNode_Bool_emitted[1]));
  assign lizzieLet12_1_3QNode_Bool_done = (lizzieLet12_1_3QNode_Bool_emitted | ({lizzieLet12_1_3QNode_Bool_2_d[0],
                                                                                 lizzieLet12_1_3QNode_Bool_1_d[0]} & {lizzieLet12_1_3QNode_Bool_2_r,
                                                                                                                      lizzieLet12_1_3QNode_Bool_1_r}));
  assign lizzieLet12_1_3QNode_Bool_r = (& lizzieLet12_1_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet12_1_3QNode_Bool_emitted <= (lizzieLet12_1_3QNode_Bool_r ? 2'd0 :
                                            lizzieLet12_1_3QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet12_1_3QNode_Bool_2,MyDTBool_Bool_Bool) > (lizzieLet12_1_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_2_bufchan_d;
  logic lizzieLet12_1_3QNode_Bool_2_bufchan_r;
  assign lizzieLet12_1_3QNode_Bool_2_r = ((! lizzieLet12_1_3QNode_Bool_2_bufchan_d[0]) || lizzieLet12_1_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QNode_Bool_2_r)
        lizzieLet12_1_3QNode_Bool_2_bufchan_d <= lizzieLet12_1_3QNode_Bool_2_d;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet12_1_3QNode_Bool_2_bufchan_r = (! lizzieLet12_1_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_3QNode_Bool_2_argbuf_d = (lizzieLet12_1_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet12_1_3QNode_Bool_2_bufchan_buf :
                                                 lizzieLet12_1_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QNode_Bool_2_argbuf_r && lizzieLet12_1_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QNode_Bool_2_argbuf_r) && (! lizzieLet12_1_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_3QNode_Bool_2_bufchan_buf <= lizzieLet12_1_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet12_1_3QVal_Bool,MyDTBool_Bool_Bool) > (lizzieLet12_1_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QVal_Bool_bufchan_d;
  logic lizzieLet12_1_3QVal_Bool_bufchan_r;
  assign lizzieLet12_1_3QVal_Bool_r = ((! lizzieLet12_1_3QVal_Bool_bufchan_d[0]) || lizzieLet12_1_3QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_3QVal_Bool_r)
        lizzieLet12_1_3QVal_Bool_bufchan_d <= lizzieLet12_1_3QVal_Bool_d;
  MyDTBool_Bool_Bool_t lizzieLet12_1_3QVal_Bool_bufchan_buf;
  assign lizzieLet12_1_3QVal_Bool_bufchan_r = (! lizzieLet12_1_3QVal_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_3QVal_Bool_1_argbuf_d = (lizzieLet12_1_3QVal_Bool_bufchan_buf[0] ? lizzieLet12_1_3QVal_Bool_bufchan_buf :
                                                lizzieLet12_1_3QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_3QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_3QVal_Bool_1_argbuf_r && lizzieLet12_1_3QVal_Bool_bufchan_buf[0]))
        lizzieLet12_1_3QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_3QVal_Bool_1_argbuf_r) && (! lizzieLet12_1_3QVal_Bool_bufchan_buf[0])))
        lizzieLet12_1_3QVal_Bool_bufchan_buf <= lizzieLet12_1_3QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet12_1_4,QTree_Bool) (go_8_goMux_data,Go) > [(lizzieLet12_1_4QNone_Bool,Go),
                                                                     (lizzieLet12_1_4QVal_Bool,Go),
                                                                     (lizzieLet12_1_4QNode_Bool,Go),
                                                                     (lizzieLet12_1_4QError_Bool,Go)] */
  logic [3:0] go_8_goMux_data_onehotd;
  always_comb
    if ((lizzieLet12_1_4_d[0] && go_8_goMux_data_d[0]))
      unique case (lizzieLet12_1_4_d[2:1])
        2'd0: go_8_goMux_data_onehotd = 4'd1;
        2'd1: go_8_goMux_data_onehotd = 4'd2;
        2'd2: go_8_goMux_data_onehotd = 4'd4;
        2'd3: go_8_goMux_data_onehotd = 4'd8;
        default: go_8_goMux_data_onehotd = 4'd0;
      endcase
    else go_8_goMux_data_onehotd = 4'd0;
  assign lizzieLet12_1_4QNone_Bool_d = go_8_goMux_data_onehotd[0];
  assign lizzieLet12_1_4QVal_Bool_d = go_8_goMux_data_onehotd[1];
  assign lizzieLet12_1_4QNode_Bool_d = go_8_goMux_data_onehotd[2];
  assign lizzieLet12_1_4QError_Bool_d = go_8_goMux_data_onehotd[3];
  assign go_8_goMux_data_r = (| (go_8_goMux_data_onehotd & {lizzieLet12_1_4QError_Bool_r,
                                                            lizzieLet12_1_4QNode_Bool_r,
                                                            lizzieLet12_1_4QVal_Bool_r,
                                                            lizzieLet12_1_4QNone_Bool_r}));
  assign lizzieLet12_1_4_r = go_8_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet12_1_4QError_Bool,Go) > [(lizzieLet12_1_4QError_Bool_1,Go),
                                                  (lizzieLet12_1_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet12_1_4QError_Bool_emitted;
  logic [1:0] lizzieLet12_1_4QError_Bool_done;
  assign lizzieLet12_1_4QError_Bool_1_d = (lizzieLet12_1_4QError_Bool_d[0] && (! lizzieLet12_1_4QError_Bool_emitted[0]));
  assign lizzieLet12_1_4QError_Bool_2_d = (lizzieLet12_1_4QError_Bool_d[0] && (! lizzieLet12_1_4QError_Bool_emitted[1]));
  assign lizzieLet12_1_4QError_Bool_done = (lizzieLet12_1_4QError_Bool_emitted | ({lizzieLet12_1_4QError_Bool_2_d[0],
                                                                                   lizzieLet12_1_4QError_Bool_1_d[0]} & {lizzieLet12_1_4QError_Bool_2_r,
                                                                                                                         lizzieLet12_1_4QError_Bool_1_r}));
  assign lizzieLet12_1_4QError_Bool_r = (& lizzieLet12_1_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet12_1_4QError_Bool_emitted <= (lizzieLet12_1_4QError_Bool_r ? 2'd0 :
                                             lizzieLet12_1_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet12_1_4QError_Bool_1,Go)] > (lizzieLet12_1_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet12_1_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet12_1_4QError_Bool_1_d[0]}), lizzieLet12_1_4QError_Bool_1_d);
  assign {lizzieLet12_1_4QError_Bool_1_r} = {1 {(lizzieLet12_1_4QError_Bool_1QError_Bool_r && lizzieLet12_1_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_1_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet17_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet12_1_4QError_Bool_1QError_Bool_r = ((! lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet12_1_4QError_Bool_1QError_Bool_r)
        lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet12_1_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet17_1_argbuf_d = (lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf :
                                   lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                              1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0,
                                                                1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet12_1_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_4QError_Bool_2,Go) > (lizzieLet12_1_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet12_1_4QError_Bool_2_bufchan_d;
  logic lizzieLet12_1_4QError_Bool_2_bufchan_r;
  assign lizzieLet12_1_4QError_Bool_2_r = ((! lizzieLet12_1_4QError_Bool_2_bufchan_d[0]) || lizzieLet12_1_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_4QError_Bool_2_r)
        lizzieLet12_1_4QError_Bool_2_bufchan_d <= lizzieLet12_1_4QError_Bool_2_d;
  Go_t lizzieLet12_1_4QError_Bool_2_bufchan_buf;
  assign lizzieLet12_1_4QError_Bool_2_bufchan_r = (! lizzieLet12_1_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_4QError_Bool_2_argbuf_d = (lizzieLet12_1_4QError_Bool_2_bufchan_buf[0] ? lizzieLet12_1_4QError_Bool_2_bufchan_buf :
                                                  lizzieLet12_1_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_4QError_Bool_2_argbuf_r && lizzieLet12_1_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_4QError_Bool_2_argbuf_r) && (! lizzieLet12_1_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_4QError_Bool_2_bufchan_buf <= lizzieLet12_1_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_4QNode_Bool,Go) > (lizzieLet12_1_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet12_1_4QNode_Bool_bufchan_d;
  logic lizzieLet12_1_4QNode_Bool_bufchan_r;
  assign lizzieLet12_1_4QNode_Bool_r = ((! lizzieLet12_1_4QNode_Bool_bufchan_d[0]) || lizzieLet12_1_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_4QNode_Bool_r)
        lizzieLet12_1_4QNode_Bool_bufchan_d <= lizzieLet12_1_4QNode_Bool_d;
  Go_t lizzieLet12_1_4QNode_Bool_bufchan_buf;
  assign lizzieLet12_1_4QNode_Bool_bufchan_r = (! lizzieLet12_1_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_4QNode_Bool_1_argbuf_d = (lizzieLet12_1_4QNode_Bool_bufchan_buf[0] ? lizzieLet12_1_4QNode_Bool_bufchan_buf :
                                                 lizzieLet12_1_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_4QNode_Bool_1_argbuf_r && lizzieLet12_1_4QNode_Bool_bufchan_buf[0]))
        lizzieLet12_1_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_4QNode_Bool_1_argbuf_r) && (! lizzieLet12_1_4QNode_Bool_bufchan_buf[0])))
        lizzieLet12_1_4QNode_Bool_bufchan_buf <= lizzieLet12_1_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet12_1_4QNone_Bool,Go) > [(lizzieLet12_1_4QNone_Bool_1,Go),
                                                 (lizzieLet12_1_4QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet12_1_4QNone_Bool_emitted;
  logic [1:0] lizzieLet12_1_4QNone_Bool_done;
  assign lizzieLet12_1_4QNone_Bool_1_d = (lizzieLet12_1_4QNone_Bool_d[0] && (! lizzieLet12_1_4QNone_Bool_emitted[0]));
  assign lizzieLet12_1_4QNone_Bool_2_d = (lizzieLet12_1_4QNone_Bool_d[0] && (! lizzieLet12_1_4QNone_Bool_emitted[1]));
  assign lizzieLet12_1_4QNone_Bool_done = (lizzieLet12_1_4QNone_Bool_emitted | ({lizzieLet12_1_4QNone_Bool_2_d[0],
                                                                                 lizzieLet12_1_4QNone_Bool_1_d[0]} & {lizzieLet12_1_4QNone_Bool_2_r,
                                                                                                                      lizzieLet12_1_4QNone_Bool_1_r}));
  assign lizzieLet12_1_4QNone_Bool_r = (& lizzieLet12_1_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet12_1_4QNone_Bool_emitted <= (lizzieLet12_1_4QNone_Bool_r ? 2'd0 :
                                            lizzieLet12_1_4QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet12_1_4QNone_Bool_1,Go)] > (lizzieLet12_1_4QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet12_1_4QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet12_1_4QNone_Bool_1_d[0]}), lizzieLet12_1_4QNone_Bool_1_d);
  assign {lizzieLet12_1_4QNone_Bool_1_r} = {1 {(lizzieLet12_1_4QNone_Bool_1QNone_Bool_r && lizzieLet12_1_4QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet12_1_4QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet13_1_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet12_1_4QNone_Bool_1QNone_Bool_r = ((! lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet12_1_4QNone_Bool_1QNone_Bool_r)
        lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet12_1_4QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet13_1_1_argbuf_d = (lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf :
                                     lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet13_1_1_argbuf_r && lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet13_1_1_argbuf_r) && (! lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet12_1_4QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet12_1_4QNone_Bool_2,Go) > (lizzieLet12_1_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet12_1_4QNone_Bool_2_bufchan_d;
  logic lizzieLet12_1_4QNone_Bool_2_bufchan_r;
  assign lizzieLet12_1_4QNone_Bool_2_r = ((! lizzieLet12_1_4QNone_Bool_2_bufchan_d[0]) || lizzieLet12_1_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_4QNone_Bool_2_r)
        lizzieLet12_1_4QNone_Bool_2_bufchan_d <= lizzieLet12_1_4QNone_Bool_2_d;
  Go_t lizzieLet12_1_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet12_1_4QNone_Bool_2_bufchan_r = (! lizzieLet12_1_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_4QNone_Bool_2_argbuf_d = (lizzieLet12_1_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet12_1_4QNone_Bool_2_bufchan_buf :
                                                 lizzieLet12_1_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_4QNone_Bool_2_argbuf_r && lizzieLet12_1_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_4QNone_Bool_2_argbuf_r) && (! lizzieLet12_1_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_4QNone_Bool_2_bufchan_buf <= lizzieLet12_1_4QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet12_1_4QNone_Bool_2_argbuf,Go),
                           (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf,Go),
                           (es_0_2_1MyFalse_1_argbuf,Go),
                           (es_0_2_1MyTrue_2_argbuf,Go),
                           (lizzieLet12_1_4QError_Bool_2_argbuf,Go)] > (go_15_goMux_choice,C5) (go_15_goMux_data,Go) */
  logic [4:0] lizzieLet12_1_4QNone_Bool_2_argbuf_select_d;
  assign lizzieLet12_1_4QNone_Bool_2_argbuf_select_d = ((| lizzieLet12_1_4QNone_Bool_2_argbuf_select_q) ? lizzieLet12_1_4QNone_Bool_2_argbuf_select_q :
                                                        (lizzieLet12_1_4QNone_Bool_2_argbuf_d[0] ? 5'd1 :
                                                         (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d [0] ? 5'd2 :
                                                          (es_0_2_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                           (es_0_2_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                            (lizzieLet12_1_4QError_Bool_2_argbuf_d[0] ? 5'd16 :
                                                             5'd0))))));
  logic [4:0] lizzieLet12_1_4QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Bool_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet12_1_4QNone_Bool_2_argbuf_select_q <= (lizzieLet12_1_4QNone_Bool_2_argbuf_done ? 5'd0 :
                                                      lizzieLet12_1_4QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q <= (lizzieLet12_1_4QNone_Bool_2_argbuf_done ? 2'd0 :
                                                    lizzieLet12_1_4QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet12_1_4QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet12_1_4QNone_Bool_2_argbuf_emit_d = (lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                                    go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                              go_15_goMux_data_r}));
  logic lizzieLet12_1_4QNone_Bool_2_argbuf_done;
  assign lizzieLet12_1_4QNone_Bool_2_argbuf_done = (& lizzieLet12_1_4QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet12_1_4QError_Bool_2_argbuf_r,
          es_0_2_1MyTrue_2_argbuf_r,
          es_0_2_1MyFalse_1_argbuf_r,
          \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ,
          lizzieLet12_1_4QNone_Bool_2_argbuf_r} = (lizzieLet12_1_4QNone_Bool_2_argbuf_done ? lizzieLet12_1_4QNone_Bool_2_argbuf_select_d :
                                                   5'd0);
  assign go_15_goMux_data_d = ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet12_1_4QNone_Bool_2_argbuf_d :
                               ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[0])) ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d  :
                                ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_2_1MyFalse_1_argbuf_d :
                                 ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_2_1MyTrue_2_argbuf_d :
                                  ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet12_1_4QError_Bool_2_argbuf_d :
                                   1'd0)))));
  assign go_15_goMux_choice_d = ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet12_1_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet12_1_4QNone_Bool_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet12_1_4QVal_Bool,Go) > [(lizzieLet12_1_4QVal_Bool_1,Go),
                                                (lizzieLet12_1_4QVal_Bool_2,Go),
                                                (lizzieLet12_1_4QVal_Bool_3,Go)] */
  logic [2:0] lizzieLet12_1_4QVal_Bool_emitted;
  logic [2:0] lizzieLet12_1_4QVal_Bool_done;
  assign lizzieLet12_1_4QVal_Bool_1_d = (lizzieLet12_1_4QVal_Bool_d[0] && (! lizzieLet12_1_4QVal_Bool_emitted[0]));
  assign lizzieLet12_1_4QVal_Bool_2_d = (lizzieLet12_1_4QVal_Bool_d[0] && (! lizzieLet12_1_4QVal_Bool_emitted[1]));
  assign lizzieLet12_1_4QVal_Bool_3_d = (lizzieLet12_1_4QVal_Bool_d[0] && (! lizzieLet12_1_4QVal_Bool_emitted[2]));
  assign lizzieLet12_1_4QVal_Bool_done = (lizzieLet12_1_4QVal_Bool_emitted | ({lizzieLet12_1_4QVal_Bool_3_d[0],
                                                                               lizzieLet12_1_4QVal_Bool_2_d[0],
                                                                               lizzieLet12_1_4QVal_Bool_1_d[0]} & {lizzieLet12_1_4QVal_Bool_3_r,
                                                                                                                   lizzieLet12_1_4QVal_Bool_2_r,
                                                                                                                   lizzieLet12_1_4QVal_Bool_1_r}));
  assign lizzieLet12_1_4QVal_Bool_r = (& lizzieLet12_1_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet12_1_4QVal_Bool_emitted <= (lizzieLet12_1_4QVal_Bool_r ? 3'd0 :
                                           lizzieLet12_1_4QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet12_1_4QVal_Bool_1,Go) > (lizzieLet12_1_4QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet12_1_4QVal_Bool_1_bufchan_d;
  logic lizzieLet12_1_4QVal_Bool_1_bufchan_r;
  assign lizzieLet12_1_4QVal_Bool_1_r = ((! lizzieLet12_1_4QVal_Bool_1_bufchan_d[0]) || lizzieLet12_1_4QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_4QVal_Bool_1_r)
        lizzieLet12_1_4QVal_Bool_1_bufchan_d <= lizzieLet12_1_4QVal_Bool_1_d;
  Go_t lizzieLet12_1_4QVal_Bool_1_bufchan_buf;
  assign lizzieLet12_1_4QVal_Bool_1_bufchan_r = (! lizzieLet12_1_4QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet12_1_4QVal_Bool_1_argbuf_d = (lizzieLet12_1_4QVal_Bool_1_bufchan_buf[0] ? lizzieLet12_1_4QVal_Bool_1_bufchan_buf :
                                                lizzieLet12_1_4QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_4QVal_Bool_1_argbuf_r && lizzieLet12_1_4QVal_Bool_1_bufchan_buf[0]))
        lizzieLet12_1_4QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_4QVal_Bool_1_argbuf_r) && (! lizzieLet12_1_4QVal_Bool_1_bufchan_buf[0])))
        lizzieLet12_1_4QVal_Bool_1_bufchan_buf <= lizzieLet12_1_4QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool_Bool___MyBool___MyBool,
      Dcon TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) : [(lizzieLet12_1_4QVal_Bool_1_argbuf,Go),
                                                            (lizzieLet12_1_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool),
                                                            (lizzieLet12_1_7QVal_Bool_1_argbuf,MyBool),
                                                            (vad2_1_argbuf,MyBool)] > (applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1,TupGo___MyDTBool_Bool_Bool___MyBool___MyBool) */
  assign applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d = TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_dc((& {lizzieLet12_1_4QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet12_1_3QVal_Bool_1_argbuf_d[0],
                                                                                                                                       lizzieLet12_1_7QVal_Bool_1_argbuf_d[0],
                                                                                                                                       vad2_1_argbuf_d[0]}), lizzieLet12_1_4QVal_Bool_1_argbuf_d, lizzieLet12_1_3QVal_Bool_1_argbuf_d, lizzieLet12_1_7QVal_Bool_1_argbuf_d, vad2_1_argbuf_d);
  assign {lizzieLet12_1_4QVal_Bool_1_argbuf_r,
          lizzieLet12_1_3QVal_Bool_1_argbuf_r,
          lizzieLet12_1_7QVal_Bool_1_argbuf_r,
          vad2_1_argbuf_r} = {4 {(applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_r && applyfnBool_Bool_Bool_5TupGo___MyDTBool_Bool_Bool___MyBool___MyBool_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet12_1_4QVal_Bool_2,Go) > (lizzieLet12_1_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet12_1_4QVal_Bool_2_bufchan_d;
  logic lizzieLet12_1_4QVal_Bool_2_bufchan_r;
  assign lizzieLet12_1_4QVal_Bool_2_r = ((! lizzieLet12_1_4QVal_Bool_2_bufchan_d[0]) || lizzieLet12_1_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_4QVal_Bool_2_r)
        lizzieLet12_1_4QVal_Bool_2_bufchan_d <= lizzieLet12_1_4QVal_Bool_2_d;
  Go_t lizzieLet12_1_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet12_1_4QVal_Bool_2_bufchan_r = (! lizzieLet12_1_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_4QVal_Bool_2_argbuf_d = (lizzieLet12_1_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet12_1_4QVal_Bool_2_bufchan_buf :
                                                lizzieLet12_1_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_4QVal_Bool_2_argbuf_r && lizzieLet12_1_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_4QVal_Bool_2_argbuf_r) && (! lizzieLet12_1_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_4QVal_Bool_2_bufchan_buf <= lizzieLet12_1_4QVal_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyBool,
      Dcon TupGo___MyDTBool_Bool___MyBool) : [(lizzieLet12_1_4QVal_Bool_2_argbuf,Go),
                                              (lizzieLet12_1_5QVal_Bool_1_argbuf,MyDTBool_Bool),
                                              (xacw_1_1_argbuf,MyBool)] > (applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1,TupGo___MyDTBool_Bool___MyBool) */
  assign applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d = TupGo___MyDTBool_Bool___MyBool_dc((& {lizzieLet12_1_4QVal_Bool_2_argbuf_d[0],
                                                                                                      lizzieLet12_1_5QVal_Bool_1_argbuf_d[0],
                                                                                                      xacw_1_1_argbuf_d[0]}), lizzieLet12_1_4QVal_Bool_2_argbuf_d, lizzieLet12_1_5QVal_Bool_1_argbuf_d, xacw_1_1_argbuf_d);
  assign {lizzieLet12_1_4QVal_Bool_2_argbuf_r,
          lizzieLet12_1_5QVal_Bool_1_argbuf_r,
          xacw_1_1_argbuf_r} = {3 {(applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_r && applyfnBool_Bool_5TupGo___MyDTBool_Bool___MyBool_1_d[0])}};
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool) : (lizzieLet12_1_5,QTree_Bool) (isZacY_goMux_mux,MyDTBool_Bool) > [(_26,MyDTBool_Bool),
                                                                                            (lizzieLet12_1_5QVal_Bool,MyDTBool_Bool),
                                                                                            (lizzieLet12_1_5QNode_Bool,MyDTBool_Bool),
                                                                                            (_25,MyDTBool_Bool)] */
  logic [3:0] isZacY_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_1_5_d[0] && isZacY_goMux_mux_d[0]))
      unique case (lizzieLet12_1_5_d[2:1])
        2'd0: isZacY_goMux_mux_onehotd = 4'd1;
        2'd1: isZacY_goMux_mux_onehotd = 4'd2;
        2'd2: isZacY_goMux_mux_onehotd = 4'd4;
        2'd3: isZacY_goMux_mux_onehotd = 4'd8;
        default: isZacY_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacY_goMux_mux_onehotd = 4'd0;
  assign _26_d = isZacY_goMux_mux_onehotd[0];
  assign lizzieLet12_1_5QVal_Bool_d = isZacY_goMux_mux_onehotd[1];
  assign lizzieLet12_1_5QNode_Bool_d = isZacY_goMux_mux_onehotd[2];
  assign _25_d = isZacY_goMux_mux_onehotd[3];
  assign isZacY_goMux_mux_r = (| (isZacY_goMux_mux_onehotd & {_25_r,
                                                              lizzieLet12_1_5QNode_Bool_r,
                                                              lizzieLet12_1_5QVal_Bool_r,
                                                              _26_r}));
  assign lizzieLet12_1_5_r = isZacY_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool) : (lizzieLet12_1_5QNode_Bool,MyDTBool_Bool) > [(lizzieLet12_1_5QNode_Bool_1,MyDTBool_Bool),
                                                                       (lizzieLet12_1_5QNode_Bool_2,MyDTBool_Bool)] */
  logic [1:0] lizzieLet12_1_5QNode_Bool_emitted;
  logic [1:0] lizzieLet12_1_5QNode_Bool_done;
  assign lizzieLet12_1_5QNode_Bool_1_d = (lizzieLet12_1_5QNode_Bool_d[0] && (! lizzieLet12_1_5QNode_Bool_emitted[0]));
  assign lizzieLet12_1_5QNode_Bool_2_d = (lizzieLet12_1_5QNode_Bool_d[0] && (! lizzieLet12_1_5QNode_Bool_emitted[1]));
  assign lizzieLet12_1_5QNode_Bool_done = (lizzieLet12_1_5QNode_Bool_emitted | ({lizzieLet12_1_5QNode_Bool_2_d[0],
                                                                                 lizzieLet12_1_5QNode_Bool_1_d[0]} & {lizzieLet12_1_5QNode_Bool_2_r,
                                                                                                                      lizzieLet12_1_5QNode_Bool_1_r}));
  assign lizzieLet12_1_5QNode_Bool_r = (& lizzieLet12_1_5QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_5QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet12_1_5QNode_Bool_emitted <= (lizzieLet12_1_5QNode_Bool_r ? 2'd0 :
                                            lizzieLet12_1_5QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet12_1_5QNode_Bool_2,MyDTBool_Bool) > (lizzieLet12_1_5QNode_Bool_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_2_bufchan_d;
  logic lizzieLet12_1_5QNode_Bool_2_bufchan_r;
  assign lizzieLet12_1_5QNode_Bool_2_r = ((! lizzieLet12_1_5QNode_Bool_2_bufchan_d[0]) || lizzieLet12_1_5QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_5QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_5QNode_Bool_2_r)
        lizzieLet12_1_5QNode_Bool_2_bufchan_d <= lizzieLet12_1_5QNode_Bool_2_d;
  MyDTBool_Bool_t lizzieLet12_1_5QNode_Bool_2_bufchan_buf;
  assign lizzieLet12_1_5QNode_Bool_2_bufchan_r = (! lizzieLet12_1_5QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_5QNode_Bool_2_argbuf_d = (lizzieLet12_1_5QNode_Bool_2_bufchan_buf[0] ? lizzieLet12_1_5QNode_Bool_2_bufchan_buf :
                                                 lizzieLet12_1_5QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_5QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_5QNode_Bool_2_argbuf_r && lizzieLet12_1_5QNode_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_5QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_5QNode_Bool_2_argbuf_r) && (! lizzieLet12_1_5QNode_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_5QNode_Bool_2_bufchan_buf <= lizzieLet12_1_5QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet12_1_5QVal_Bool,MyDTBool_Bool) > (lizzieLet12_1_5QVal_Bool_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet12_1_5QVal_Bool_bufchan_d;
  logic lizzieLet12_1_5QVal_Bool_bufchan_r;
  assign lizzieLet12_1_5QVal_Bool_r = ((! lizzieLet12_1_5QVal_Bool_bufchan_d[0]) || lizzieLet12_1_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_5QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet12_1_5QVal_Bool_r)
        lizzieLet12_1_5QVal_Bool_bufchan_d <= lizzieLet12_1_5QVal_Bool_d;
  MyDTBool_Bool_t lizzieLet12_1_5QVal_Bool_bufchan_buf;
  assign lizzieLet12_1_5QVal_Bool_bufchan_r = (! lizzieLet12_1_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_5QVal_Bool_1_argbuf_d = (lizzieLet12_1_5QVal_Bool_bufchan_buf[0] ? lizzieLet12_1_5QVal_Bool_bufchan_buf :
                                                lizzieLet12_1_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_5QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet12_1_5QVal_Bool_1_argbuf_r && lizzieLet12_1_5QVal_Bool_bufchan_buf[0]))
        lizzieLet12_1_5QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet12_1_5QVal_Bool_1_argbuf_r) && (! lizzieLet12_1_5QVal_Bool_bufchan_buf[0])))
        lizzieLet12_1_5QVal_Bool_bufchan_buf <= lizzieLet12_1_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet12_1_6,QTree_Bool) (sc_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) > [(lizzieLet12_1_6QNone_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet12_1_6QVal_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet12_1_6QNode_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                          (lizzieLet12_1_6QError_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet12_1_6_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet12_1_6_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet12_1_6QNone_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                        sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet12_1_6QVal_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                       sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet12_1_6QNode_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                        sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet12_1_6QError_Bool_d = {sc_0_2_goMux_mux_d[16:1],
                                         sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet12_1_6QError_Bool_r,
                                                              lizzieLet12_1_6QNode_Bool_r,
                                                              lizzieLet12_1_6QVal_Bool_r,
                                                              lizzieLet12_1_6QNone_Bool_r}));
  assign lizzieLet12_1_6_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet12_1_6QError_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet12_1_6QError_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QError_Bool_bufchan_d;
  logic lizzieLet12_1_6QError_Bool_bufchan_r;
  assign lizzieLet12_1_6QError_Bool_r = ((! lizzieLet12_1_6QError_Bool_bufchan_d[0]) || lizzieLet12_1_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_6QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_1_6QError_Bool_r)
        lizzieLet12_1_6QError_Bool_bufchan_d <= lizzieLet12_1_6QError_Bool_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QError_Bool_bufchan_buf;
  assign lizzieLet12_1_6QError_Bool_bufchan_r = (! lizzieLet12_1_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_6QError_Bool_1_argbuf_d = (lizzieLet12_1_6QError_Bool_bufchan_buf[0] ? lizzieLet12_1_6QError_Bool_bufchan_buf :
                                                  lizzieLet12_1_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_6QError_Bool_1_argbuf_r && lizzieLet12_1_6QError_Bool_bufchan_buf[0]))
        lizzieLet12_1_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_6QError_Bool_1_argbuf_r) && (! lizzieLet12_1_6QError_Bool_bufchan_buf[0])))
        lizzieLet12_1_6QError_Bool_bufchan_buf <= lizzieLet12_1_6QError_Bool_bufchan_d;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool3) : [(lizzieLet12_1_6QNode_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (lizzieLet12_1_5QNode_Bool_1,MyDTBool_Bool),
                                                 (lizzieLet12_1_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                 (lizzieLet12_1_7QNode_Bool_1,MyBool),
                                                 (q1ad3_destruct,Pointer_QTree_Bool),
                                                 (q2ad4_destruct,Pointer_QTree_Bool),
                                                 (q3ad5_destruct,Pointer_QTree_Bool)] > (lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_d  = \Lcall_map''_map''_Bool_Bool_Bool3_dc ((& {lizzieLet12_1_6QNode_Bool_d[0],
                                                                                                                                                                                                                             lizzieLet12_1_5QNode_Bool_1_d[0],
                                                                                                                                                                                                                             lizzieLet12_1_3QNode_Bool_1_d[0],
                                                                                                                                                                                                                             lizzieLet12_1_7QNode_Bool_1_d[0],
                                                                                                                                                                                                                             q1ad3_destruct_d[0],
                                                                                                                                                                                                                             q2ad4_destruct_d[0],
                                                                                                                                                                                                                             q3ad5_destruct_d[0]}), lizzieLet12_1_6QNode_Bool_d, lizzieLet12_1_5QNode_Bool_1_d, lizzieLet12_1_3QNode_Bool_1_d, lizzieLet12_1_7QNode_Bool_1_d, q1ad3_destruct_d, q2ad4_destruct_d, q3ad5_destruct_d);
  assign {lizzieLet12_1_6QNode_Bool_r,
          lizzieLet12_1_5QNode_Bool_1_r,
          lizzieLet12_1_3QNode_Bool_1_r,
          lizzieLet12_1_7QNode_Bool_1_r,
          q1ad3_destruct_r,
          q2ad4_destruct_r,
          q3ad5_destruct_r} = {7 {(\lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_r  && \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet16_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  logic \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r ;
  assign \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_r  = ((! \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d [0]) || \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= {68'd0,
                                                                                                                                                                                         1'd0};
    else
      if (\lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_r )
        \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf ;
  assign \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r  = (! \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]);
  assign lizzieLet16_1_argbuf_d = (\lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0] ? \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  :
                                   \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= {68'd0,
                                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]))
        \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= {68'd0,
                                                                                                                                                                                             1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0])))
        \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= \lizzieLet12_1_6QNode_Bool_1lizzieLet12_1_5QNode_Bool_1lizzieLet12_1_3QNode_Bool_1lizzieLet12_1_7QNode_Bool_1q1ad3_1q2ad4_1q3ad5_1Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (lizzieLet12_1_6QNone_Bool,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet12_1_6QNone_Bool_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QNone_Bool_bufchan_d;
  logic lizzieLet12_1_6QNone_Bool_bufchan_r;
  assign lizzieLet12_1_6QNone_Bool_r = ((! lizzieLet12_1_6QNone_Bool_bufchan_d[0]) || lizzieLet12_1_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet12_1_6QNone_Bool_r)
        lizzieLet12_1_6QNone_Bool_bufchan_d <= lizzieLet12_1_6QNone_Bool_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  lizzieLet12_1_6QNone_Bool_bufchan_buf;
  assign lizzieLet12_1_6QNone_Bool_bufchan_r = (! lizzieLet12_1_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_6QNone_Bool_1_argbuf_d = (lizzieLet12_1_6QNone_Bool_bufchan_buf[0] ? lizzieLet12_1_6QNone_Bool_bufchan_buf :
                                                 lizzieLet12_1_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_6QNone_Bool_1_argbuf_r && lizzieLet12_1_6QNone_Bool_bufchan_buf[0]))
        lizzieLet12_1_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_6QNone_Bool_1_argbuf_r) && (! lizzieLet12_1_6QNone_Bool_bufchan_buf[0])))
        lizzieLet12_1_6QNone_Bool_bufchan_buf <= lizzieLet12_1_6QNone_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyBool) : (lizzieLet12_1_7,QTree_Bool) (v'ad0_goMux_mux,MyBool) > [(_24,MyBool),
                                                                             (lizzieLet12_1_7QVal_Bool,MyBool),
                                                                             (lizzieLet12_1_7QNode_Bool,MyBool),
                                                                             (_23,MyBool)] */
  logic [3:0] \v'ad0_goMux_mux_onehotd ;
  always_comb
    if ((lizzieLet12_1_7_d[0] && \v'ad0_goMux_mux_d [0]))
      unique case (lizzieLet12_1_7_d[2:1])
        2'd0: \v'ad0_goMux_mux_onehotd  = 4'd1;
        2'd1: \v'ad0_goMux_mux_onehotd  = 4'd2;
        2'd2: \v'ad0_goMux_mux_onehotd  = 4'd4;
        2'd3: \v'ad0_goMux_mux_onehotd  = 4'd8;
        default: \v'ad0_goMux_mux_onehotd  = 4'd0;
      endcase
    else \v'ad0_goMux_mux_onehotd  = 4'd0;
  assign _24_d = {\v'ad0_goMux_mux_d [1:1],
                  \v'ad0_goMux_mux_onehotd [0]};
  assign lizzieLet12_1_7QVal_Bool_d = {\v'ad0_goMux_mux_d [1:1],
                                       \v'ad0_goMux_mux_onehotd [1]};
  assign lizzieLet12_1_7QNode_Bool_d = {\v'ad0_goMux_mux_d [1:1],
                                        \v'ad0_goMux_mux_onehotd [2]};
  assign _23_d = {\v'ad0_goMux_mux_d [1:1],
                  \v'ad0_goMux_mux_onehotd [3]};
  assign \v'ad0_goMux_mux_r  = (| (\v'ad0_goMux_mux_onehotd  & {_23_r,
                                                                lizzieLet12_1_7QNode_Bool_r,
                                                                lizzieLet12_1_7QVal_Bool_r,
                                                                _24_r}));
  assign lizzieLet12_1_7_r = \v'ad0_goMux_mux_r ;
  
  /* fork (Ty MyBool) : (lizzieLet12_1_7QNode_Bool,MyBool) > [(lizzieLet12_1_7QNode_Bool_1,MyBool),
                                                         (lizzieLet12_1_7QNode_Bool_2,MyBool)] */
  logic [1:0] lizzieLet12_1_7QNode_Bool_emitted;
  logic [1:0] lizzieLet12_1_7QNode_Bool_done;
  assign lizzieLet12_1_7QNode_Bool_1_d = {lizzieLet12_1_7QNode_Bool_d[1:1],
                                          (lizzieLet12_1_7QNode_Bool_d[0] && (! lizzieLet12_1_7QNode_Bool_emitted[0]))};
  assign lizzieLet12_1_7QNode_Bool_2_d = {lizzieLet12_1_7QNode_Bool_d[1:1],
                                          (lizzieLet12_1_7QNode_Bool_d[0] && (! lizzieLet12_1_7QNode_Bool_emitted[1]))};
  assign lizzieLet12_1_7QNode_Bool_done = (lizzieLet12_1_7QNode_Bool_emitted | ({lizzieLet12_1_7QNode_Bool_2_d[0],
                                                                                 lizzieLet12_1_7QNode_Bool_1_d[0]} & {lizzieLet12_1_7QNode_Bool_2_r,
                                                                                                                      lizzieLet12_1_7QNode_Bool_1_r}));
  assign lizzieLet12_1_7QNode_Bool_r = (& lizzieLet12_1_7QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet12_1_7QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet12_1_7QNode_Bool_emitted <= (lizzieLet12_1_7QNode_Bool_r ? 2'd0 :
                                            lizzieLet12_1_7QNode_Bool_done);
  
  /* buf (Ty MyBool) : (lizzieLet12_1_7QNode_Bool_2,MyBool) > (lizzieLet12_1_7QNode_Bool_2_argbuf,MyBool) */
  MyBool_t lizzieLet12_1_7QNode_Bool_2_bufchan_d;
  logic lizzieLet12_1_7QNode_Bool_2_bufchan_r;
  assign lizzieLet12_1_7QNode_Bool_2_r = ((! lizzieLet12_1_7QNode_Bool_2_bufchan_d[0]) || lizzieLet12_1_7QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_7QNode_Bool_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet12_1_7QNode_Bool_2_r)
        lizzieLet12_1_7QNode_Bool_2_bufchan_d <= lizzieLet12_1_7QNode_Bool_2_d;
  MyBool_t lizzieLet12_1_7QNode_Bool_2_bufchan_buf;
  assign lizzieLet12_1_7QNode_Bool_2_bufchan_r = (! lizzieLet12_1_7QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet12_1_7QNode_Bool_2_argbuf_d = (lizzieLet12_1_7QNode_Bool_2_bufchan_buf[0] ? lizzieLet12_1_7QNode_Bool_2_bufchan_buf :
                                                 lizzieLet12_1_7QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_7QNode_Bool_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet12_1_7QNode_Bool_2_argbuf_r && lizzieLet12_1_7QNode_Bool_2_bufchan_buf[0]))
        lizzieLet12_1_7QNode_Bool_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet12_1_7QNode_Bool_2_argbuf_r) && (! lizzieLet12_1_7QNode_Bool_2_bufchan_buf[0])))
        lizzieLet12_1_7QNode_Bool_2_bufchan_buf <= lizzieLet12_1_7QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyBool) : (lizzieLet12_1_7QVal_Bool,MyBool) > (lizzieLet12_1_7QVal_Bool_1_argbuf,MyBool) */
  MyBool_t lizzieLet12_1_7QVal_Bool_bufchan_d;
  logic lizzieLet12_1_7QVal_Bool_bufchan_r;
  assign lizzieLet12_1_7QVal_Bool_r = ((! lizzieLet12_1_7QVal_Bool_bufchan_d[0]) || lizzieLet12_1_7QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_7QVal_Bool_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet12_1_7QVal_Bool_r)
        lizzieLet12_1_7QVal_Bool_bufchan_d <= lizzieLet12_1_7QVal_Bool_d;
  MyBool_t lizzieLet12_1_7QVal_Bool_bufchan_buf;
  assign lizzieLet12_1_7QVal_Bool_bufchan_r = (! lizzieLet12_1_7QVal_Bool_bufchan_buf[0]);
  assign lizzieLet12_1_7QVal_Bool_1_argbuf_d = (lizzieLet12_1_7QVal_Bool_bufchan_buf[0] ? lizzieLet12_1_7QVal_Bool_bufchan_buf :
                                                lizzieLet12_1_7QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet12_1_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet12_1_7QVal_Bool_1_argbuf_r && lizzieLet12_1_7QVal_Bool_bufchan_buf[0]))
        lizzieLet12_1_7QVal_Bool_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet12_1_7QVal_Bool_1_argbuf_r) && (! lizzieLet12_1_7QVal_Bool_bufchan_buf[0])))
        lizzieLet12_1_7QVal_Bool_bufchan_buf <= lizzieLet12_1_7QVal_Bool_bufchan_d;
  
  /* destruct (Ty Nat,
          Dcon Succ) : (lizzieLet18_1Succ,Nat) > [(x1adj_destruct,Pointer_Nat)] */
  assign x1adj_destruct_d = {lizzieLet18_1Succ_d[17:2],
                             lizzieLet18_1Succ_d[0]};
  assign lizzieLet18_1Succ_r = x1adj_destruct_r;
  
  /* demux (Ty Nat,
       Ty Nat) : (lizzieLet18_2,Nat) (lizzieLet18_1,Nat) > [(_22,Nat),
                                                            (lizzieLet18_1Succ,Nat)] */
  logic [1:0] lizzieLet18_1_onehotd;
  always_comb
    if ((lizzieLet18_2_d[0] && lizzieLet18_1_d[0]))
      unique case (lizzieLet18_2_d[1:1])
        1'd0: lizzieLet18_1_onehotd = 2'd1;
        1'd1: lizzieLet18_1_onehotd = 2'd2;
        default: lizzieLet18_1_onehotd = 2'd0;
      endcase
    else lizzieLet18_1_onehotd = 2'd0;
  assign _22_d = {lizzieLet18_1_d[17:1], lizzieLet18_1_onehotd[0]};
  assign lizzieLet18_1Succ_d = {lizzieLet18_1_d[17:1],
                                lizzieLet18_1_onehotd[1]};
  assign lizzieLet18_1_r = (| (lizzieLet18_1_onehotd & {lizzieLet18_1Succ_r,
                                                        _22_r}));
  assign lizzieLet18_2_r = lizzieLet18_1_r;
  
  /* demux (Ty Nat,
       Ty Go) : (lizzieLet18_3,Nat) (go_9_goMux_data,Go) > [(lizzieLet18_3Zero,Go),
                                                            (lizzieLet18_3Succ,Go)] */
  logic [1:0] go_9_goMux_data_onehotd;
  always_comb
    if ((lizzieLet18_3_d[0] && go_9_goMux_data_d[0]))
      unique case (lizzieLet18_3_d[1:1])
        1'd0: go_9_goMux_data_onehotd = 2'd1;
        1'd1: go_9_goMux_data_onehotd = 2'd2;
        default: go_9_goMux_data_onehotd = 2'd0;
      endcase
    else go_9_goMux_data_onehotd = 2'd0;
  assign lizzieLet18_3Zero_d = go_9_goMux_data_onehotd[0];
  assign lizzieLet18_3Succ_d = go_9_goMux_data_onehotd[1];
  assign go_9_goMux_data_r = (| (go_9_goMux_data_onehotd & {lizzieLet18_3Succ_r,
                                                            lizzieLet18_3Zero_r}));
  assign lizzieLet18_3_r = go_9_goMux_data_r;
  
  /* demux (Ty Nat,
       Ty Nat) : (lizzieLet18_4,Nat) (readPointer_Natyadh_1_argbuf_rwb,Nat) > [(lizzieLet18_4Zero,Nat),
                                                                               (lizzieLet18_4Succ,Nat)] */
  logic [1:0] readPointer_Natyadh_1_argbuf_rwb_onehotd;
  always_comb
    if ((lizzieLet18_4_d[0] && readPointer_Natyadh_1_argbuf_rwb_d[0]))
      unique case (lizzieLet18_4_d[1:1])
        1'd0: readPointer_Natyadh_1_argbuf_rwb_onehotd = 2'd1;
        1'd1: readPointer_Natyadh_1_argbuf_rwb_onehotd = 2'd2;
        default: readPointer_Natyadh_1_argbuf_rwb_onehotd = 2'd0;
      endcase
    else readPointer_Natyadh_1_argbuf_rwb_onehotd = 2'd0;
  assign lizzieLet18_4Zero_d = {readPointer_Natyadh_1_argbuf_rwb_d[17:1],
                                readPointer_Natyadh_1_argbuf_rwb_onehotd[0]};
  assign lizzieLet18_4Succ_d = {readPointer_Natyadh_1_argbuf_rwb_d[17:1],
                                readPointer_Natyadh_1_argbuf_rwb_onehotd[1]};
  assign readPointer_Natyadh_1_argbuf_rwb_r = (| (readPointer_Natyadh_1_argbuf_rwb_onehotd & {lizzieLet18_4Succ_r,
                                                                                              lizzieLet18_4Zero_r}));
  assign lizzieLet18_4_r = readPointer_Natyadh_1_argbuf_rwb_r;
  
  /* fork (Ty Nat) : (lizzieLet18_4Succ,Nat) > [(lizzieLet18_4Succ_1,Nat),
                                           (lizzieLet18_4Succ_2,Nat),
                                           (lizzieLet18_4Succ_3,Nat),
                                           (lizzieLet18_4Succ_4,Nat)] */
  logic [3:0] lizzieLet18_4Succ_emitted;
  logic [3:0] lizzieLet18_4Succ_done;
  assign lizzieLet18_4Succ_1_d = {lizzieLet18_4Succ_d[17:1],
                                  (lizzieLet18_4Succ_d[0] && (! lizzieLet18_4Succ_emitted[0]))};
  assign lizzieLet18_4Succ_2_d = {lizzieLet18_4Succ_d[17:1],
                                  (lizzieLet18_4Succ_d[0] && (! lizzieLet18_4Succ_emitted[1]))};
  assign lizzieLet18_4Succ_3_d = {lizzieLet18_4Succ_d[17:1],
                                  (lizzieLet18_4Succ_d[0] && (! lizzieLet18_4Succ_emitted[2]))};
  assign lizzieLet18_4Succ_4_d = {lizzieLet18_4Succ_d[17:1],
                                  (lizzieLet18_4Succ_d[0] && (! lizzieLet18_4Succ_emitted[3]))};
  assign lizzieLet18_4Succ_done = (lizzieLet18_4Succ_emitted | ({lizzieLet18_4Succ_4_d[0],
                                                                 lizzieLet18_4Succ_3_d[0],
                                                                 lizzieLet18_4Succ_2_d[0],
                                                                 lizzieLet18_4Succ_1_d[0]} & {lizzieLet18_4Succ_4_r,
                                                                                              lizzieLet18_4Succ_3_r,
                                                                                              lizzieLet18_4Succ_2_r,
                                                                                              lizzieLet18_4Succ_1_r}));
  assign lizzieLet18_4Succ_r = (& lizzieLet18_4Succ_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_4Succ_emitted <= 4'd0;
    else
      lizzieLet18_4Succ_emitted <= (lizzieLet18_4Succ_r ? 4'd0 :
                                    lizzieLet18_4Succ_done);
  
  /* destruct (Ty Nat,
          Dcon Succ) : (lizzieLet18_4Succ_1Succ,Nat) > [(y1adk_destruct,Pointer_Nat)] */
  assign y1adk_destruct_d = {lizzieLet18_4Succ_1Succ_d[17:2],
                             lizzieLet18_4Succ_1Succ_d[0]};
  assign lizzieLet18_4Succ_1Succ_r = y1adk_destruct_r;
  
  /* demux (Ty Nat,
       Ty Nat) : (lizzieLet18_4Succ_2,Nat) (lizzieLet18_4Succ_1,Nat) > [(_21,Nat),
                                                                        (lizzieLet18_4Succ_1Succ,Nat)] */
  logic [1:0] lizzieLet18_4Succ_1_onehotd;
  always_comb
    if ((lizzieLet18_4Succ_2_d[0] && lizzieLet18_4Succ_1_d[0]))
      unique case (lizzieLet18_4Succ_2_d[1:1])
        1'd0: lizzieLet18_4Succ_1_onehotd = 2'd1;
        1'd1: lizzieLet18_4Succ_1_onehotd = 2'd2;
        default: lizzieLet18_4Succ_1_onehotd = 2'd0;
      endcase
    else lizzieLet18_4Succ_1_onehotd = 2'd0;
  assign _21_d = {lizzieLet18_4Succ_1_d[17:1],
                  lizzieLet18_4Succ_1_onehotd[0]};
  assign lizzieLet18_4Succ_1Succ_d = {lizzieLet18_4Succ_1_d[17:1],
                                      lizzieLet18_4Succ_1_onehotd[1]};
  assign lizzieLet18_4Succ_1_r = (| (lizzieLet18_4Succ_1_onehotd & {lizzieLet18_4Succ_1Succ_r,
                                                                    _21_r}));
  assign lizzieLet18_4Succ_2_r = lizzieLet18_4Succ_1_r;
  
  /* demux (Ty Nat,
       Ty Go) : (lizzieLet18_4Succ_3,Nat) (lizzieLet18_3Succ,Go) > [(lizzieLet18_4Succ_3Zero,Go),
                                                                    (lizzieLet18_4Succ_3Succ,Go)] */
  logic [1:0] lizzieLet18_3Succ_onehotd;
  always_comb
    if ((lizzieLet18_4Succ_3_d[0] && lizzieLet18_3Succ_d[0]))
      unique case (lizzieLet18_4Succ_3_d[1:1])
        1'd0: lizzieLet18_3Succ_onehotd = 2'd1;
        1'd1: lizzieLet18_3Succ_onehotd = 2'd2;
        default: lizzieLet18_3Succ_onehotd = 2'd0;
      endcase
    else lizzieLet18_3Succ_onehotd = 2'd0;
  assign lizzieLet18_4Succ_3Zero_d = lizzieLet18_3Succ_onehotd[0];
  assign lizzieLet18_4Succ_3Succ_d = lizzieLet18_3Succ_onehotd[1];
  assign lizzieLet18_3Succ_r = (| (lizzieLet18_3Succ_onehotd & {lizzieLet18_4Succ_3Succ_r,
                                                                lizzieLet18_4Succ_3Zero_r}));
  assign lizzieLet18_4Succ_3_r = lizzieLet18_3Succ_r;
  
  /* buf (Ty Go) : (lizzieLet18_4Succ_3Succ,Go) > (lizzieLet18_4Succ_3Succ_1_argbuf,Go) */
  Go_t lizzieLet18_4Succ_3Succ_bufchan_d;
  logic lizzieLet18_4Succ_3Succ_bufchan_r;
  assign lizzieLet18_4Succ_3Succ_r = ((! lizzieLet18_4Succ_3Succ_bufchan_d[0]) || lizzieLet18_4Succ_3Succ_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_4Succ_3Succ_bufchan_d <= 1'd0;
    else
      if (lizzieLet18_4Succ_3Succ_r)
        lizzieLet18_4Succ_3Succ_bufchan_d <= lizzieLet18_4Succ_3Succ_d;
  Go_t lizzieLet18_4Succ_3Succ_bufchan_buf;
  assign lizzieLet18_4Succ_3Succ_bufchan_r = (! lizzieLet18_4Succ_3Succ_bufchan_buf[0]);
  assign lizzieLet18_4Succ_3Succ_1_argbuf_d = (lizzieLet18_4Succ_3Succ_bufchan_buf[0] ? lizzieLet18_4Succ_3Succ_bufchan_buf :
                                               lizzieLet18_4Succ_3Succ_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet18_4Succ_3Succ_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet18_4Succ_3Succ_1_argbuf_r && lizzieLet18_4Succ_3Succ_bufchan_buf[0]))
        lizzieLet18_4Succ_3Succ_bufchan_buf <= 1'd0;
      else if (((! lizzieLet18_4Succ_3Succ_1_argbuf_r) && (! lizzieLet18_4Succ_3Succ_bufchan_buf[0])))
        lizzieLet18_4Succ_3Succ_bufchan_buf <= lizzieLet18_4Succ_3Succ_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet18_4Succ_3Zero,Go)] > (lizzieLet18_4Succ_3Zero_1MyFalse,MyBool) */
  assign lizzieLet18_4Succ_3Zero_1MyFalse_d = MyFalse_dc((& {lizzieLet18_4Succ_3Zero_d[0]}), lizzieLet18_4Succ_3Zero_d);
  assign {lizzieLet18_4Succ_3Zero_r} = {1 {(lizzieLet18_4Succ_3Zero_1MyFalse_r && lizzieLet18_4Succ_3Zero_1MyFalse_d[0])}};
  
  /* demux (Ty Nat,
       Ty Pointer_Nat) : (lizzieLet18_4Succ_4,Nat) (x1adj_destruct,Pointer_Nat) > [(_20,Pointer_Nat),
                                                                                   (lizzieLet18_4Succ_4Succ,Pointer_Nat)] */
  logic [1:0] x1adj_destruct_onehotd;
  always_comb
    if ((lizzieLet18_4Succ_4_d[0] && x1adj_destruct_d[0]))
      unique case (lizzieLet18_4Succ_4_d[1:1])
        1'd0: x1adj_destruct_onehotd = 2'd1;
        1'd1: x1adj_destruct_onehotd = 2'd2;
        default: x1adj_destruct_onehotd = 2'd0;
      endcase
    else x1adj_destruct_onehotd = 2'd0;
  assign _20_d = {x1adj_destruct_d[16:1], x1adj_destruct_onehotd[0]};
  assign lizzieLet18_4Succ_4Succ_d = {x1adj_destruct_d[16:1],
                                      x1adj_destruct_onehotd[1]};
  assign x1adj_destruct_r = (| (x1adj_destruct_onehotd & {lizzieLet18_4Succ_4Succ_r,
                                                          _20_r}));
  assign lizzieLet18_4Succ_4_r = x1adj_destruct_r;
  
  /* buf (Ty Pointer_Nat) : (lizzieLet18_4Succ_4Succ,Pointer_Nat) > (lizzieLet18_4Succ_4Succ_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t lizzieLet18_4Succ_4Succ_bufchan_d;
  logic lizzieLet18_4Succ_4Succ_bufchan_r;
  assign lizzieLet18_4Succ_4Succ_r = ((! lizzieLet18_4Succ_4Succ_bufchan_d[0]) || lizzieLet18_4Succ_4Succ_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet18_4Succ_4Succ_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet18_4Succ_4Succ_r)
        lizzieLet18_4Succ_4Succ_bufchan_d <= lizzieLet18_4Succ_4Succ_d;
  Pointer_Nat_t lizzieLet18_4Succ_4Succ_bufchan_buf;
  assign lizzieLet18_4Succ_4Succ_bufchan_r = (! lizzieLet18_4Succ_4Succ_bufchan_buf[0]);
  assign lizzieLet18_4Succ_4Succ_1_argbuf_d = (lizzieLet18_4Succ_4Succ_bufchan_buf[0] ? lizzieLet18_4Succ_4Succ_bufchan_buf :
                                               lizzieLet18_4Succ_4Succ_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet18_4Succ_4Succ_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet18_4Succ_4Succ_1_argbuf_r && lizzieLet18_4Succ_4Succ_bufchan_buf[0]))
        lizzieLet18_4Succ_4Succ_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet18_4Succ_4Succ_1_argbuf_r) && (! lizzieLet18_4Succ_4Succ_bufchan_buf[0])))
        lizzieLet18_4Succ_4Succ_bufchan_buf <= lizzieLet18_4Succ_4Succ_bufchan_d;
  
  /* demux (Ty Nat,
       Ty Go) : (lizzieLet18_4Zero,Nat) (lizzieLet18_3Zero,Go) > [(lizzieLet18_4Zero_1Zero,Go),
                                                                  (lizzieLet18_4Zero_1Succ,Go)] */
  logic [1:0] lizzieLet18_3Zero_onehotd;
  always_comb
    if ((lizzieLet18_4Zero_d[0] && lizzieLet18_3Zero_d[0]))
      unique case (lizzieLet18_4Zero_d[1:1])
        1'd0: lizzieLet18_3Zero_onehotd = 2'd1;
        1'd1: lizzieLet18_3Zero_onehotd = 2'd2;
        default: lizzieLet18_3Zero_onehotd = 2'd0;
      endcase
    else lizzieLet18_3Zero_onehotd = 2'd0;
  assign lizzieLet18_4Zero_1Zero_d = lizzieLet18_3Zero_onehotd[0];
  assign lizzieLet18_4Zero_1Succ_d = lizzieLet18_3Zero_onehotd[1];
  assign lizzieLet18_3Zero_r = (| (lizzieLet18_3Zero_onehotd & {lizzieLet18_4Zero_1Succ_r,
                                                                lizzieLet18_4Zero_1Zero_r}));
  assign lizzieLet18_4Zero_r = lizzieLet18_3Zero_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet18_4Zero_1Succ,Go)] > (lizzieLet18_4Zero_1Succ_1MyFalse,MyBool) */
  assign lizzieLet18_4Zero_1Succ_1MyFalse_d = MyFalse_dc((& {lizzieLet18_4Zero_1Succ_d[0]}), lizzieLet18_4Zero_1Succ_d);
  assign {lizzieLet18_4Zero_1Succ_r} = {1 {(lizzieLet18_4Zero_1Succ_1MyFalse_r && lizzieLet18_4Zero_1Succ_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet18_4Zero_1Zero,Go)] > (lizzieLet18_4Zero_1Zero_1MyTrue,MyBool) */
  assign lizzieLet18_4Zero_1Zero_1MyTrue_d = MyTrue_dc((& {lizzieLet18_4Zero_1Zero_d[0]}), lizzieLet18_4Zero_1Zero_d);
  assign {lizzieLet18_4Zero_1Zero_r} = {1 {(lizzieLet18_4Zero_1Zero_1MyTrue_r && lizzieLet18_4Zero_1Zero_1MyTrue_d[0])}};
  
  /* merge (Ty MyBool) : [(lizzieLet18_4Zero_1Zero_1MyTrue,MyBool),
                     (lizzieLet18_4Zero_1Succ_1MyFalse,MyBool)] > (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge,MyBool) */
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected;
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_select;
  always_comb
    begin
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected = 2'd0;
      if ((| lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_select))
        lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected = lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_select;
      else
        if (lizzieLet18_4Zero_1Zero_1MyTrue_d[0])
          lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected[0] = 1'd1;
        else if (lizzieLet18_4Zero_1Succ_1MyFalse_d[0])
          lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_select <= 2'd0;
    else
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_select <= (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_r ? 2'd0 :
                                                                                       lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected);
  always_comb
    if (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected[0])
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d = lizzieLet18_4Zero_1Zero_1MyTrue_d;
    else if (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected[1])
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d = lizzieLet18_4Zero_1Succ_1MyFalse_d;
    else
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d = {1'd0,
                                                                                 1'd0};
  assign {lizzieLet18_4Zero_1Succ_1MyFalse_r,
          lizzieLet18_4Zero_1Zero_1MyTrue_r} = (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_r ? lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_selected :
                                                2'd0);
  
  /* merge (Ty MyBool) : [(lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge,MyBool),
                     (lizzieLet18_4Succ_3Zero_1MyFalse,MyBool)] > (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge,MyBool) */
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected;
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_select;
  always_comb
    begin
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected = 2'd0;
      if ((| lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_select))
        lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected = lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_select;
      else
        if (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d[0])
          lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected[0] = 1'd1;
        else if (lizzieLet18_4Succ_3Zero_1MyFalse_d[0])
          lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_select <= 2'd0;
    else
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_select <= (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_r ? 2'd0 :
                                                                                                                                   lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected);
  always_comb
    if (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected[0])
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d = lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_d;
    else if (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected[1])
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d = lizzieLet18_4Succ_3Zero_1MyFalse_d;
    else
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d = {1'd0,
                                                                                                                             1'd0};
  assign {lizzieLet18_4Succ_3Zero_1MyFalse_r,
          lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_merge_r} = (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_r ? lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_selected :
                                                                                      2'd0);
  
  /* fork (Ty MyBool) : (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge,MyBool) > [(lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1,MyBool),
                                                                                                                                                 (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2,MyBool)] */
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted;
  logic [1:0] lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_done;
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_d = {lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d[1:1],
                                                                                                                                       (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d[0] && (! lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted[0]))};
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d = {lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d[1:1],
                                                                                                                                       (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_d[0] && (! lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted[1]))};
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_done = (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted | ({lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_d[0],
                                                                                                                                                                                                                                                                 lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_d[0]} & {lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_2_r,
                                                                                                                                                                                                                                                                                                                                                                                                   lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_r}));
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_r = (& lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted <= 2'd0;
    else
      lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_emitted <= (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_r ? 2'd0 :
                                                                                                                                    lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_done);
  
  /* togo (Ty MyBool) : (lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1,MyBool) > (eqNat_goConst,Go) */
  assign eqNat_goConst_d = lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_d[0];
  assign lizzieLet18_4Zero_1Zero_1MyTruelizzieLet18_4Zero_1Succ_1MyFalse_mergelizzieLet18_4Succ_3Zero_1MyFalse_merge_merge_fork_1_r = eqNat_goConst_r;
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool0) : (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) > [(es_1_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_2_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_3_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_6_destruct,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted;
  logic [3:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_done;
  assign es_1_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[19:4],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[0]))};
  assign es_2_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[35:20],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[1]))};
  assign es_3_3_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[51:36],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[67:52],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted[3]))};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_done = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted | ({sc_0_6_destruct_d[0],
                                                                                                                       es_3_3_destruct_d[0],
                                                                                                                       es_2_2_destruct_d[0],
                                                                                                                       es_1_2_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                                                                es_3_3_destruct_r,
                                                                                                                                                es_2_2_destruct_r,
                                                                                                                                                es_1_2_destruct_r}));
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_r = (& lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted <= 4'd0;
    else
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_emitted <= (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_r ? 4'd0 :
                                                               lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool1) : (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) > [(es_2_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (es_3_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_5_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZad7_4_destruct,MyDTBool_Bool),
                                                                                                                               (gad8_4_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1adc_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2ada_4_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted;
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_done;
  assign es_2_1_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[19:4],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[35:20],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[51:36],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[2]))};
  assign isZad7_4_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[3]));
  assign gad8_4_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[4]));
  assign q1adc_3_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[67:52],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[5]))};
  assign m2ada_4_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[83:68],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted[6]))};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_done = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted | ({m2ada_4_destruct_d[0],
                                                                                                                       q1adc_3_destruct_d[0],
                                                                                                                       gad8_4_destruct_d[0],
                                                                                                                       isZad7_4_destruct_d[0],
                                                                                                                       sc_0_5_destruct_d[0],
                                                                                                                       es_3_2_destruct_d[0],
                                                                                                                       es_2_1_destruct_d[0]} & {m2ada_4_destruct_r,
                                                                                                                                                q1adc_3_destruct_r,
                                                                                                                                                gad8_4_destruct_r,
                                                                                                                                                isZad7_4_destruct_r,
                                                                                                                                                sc_0_5_destruct_r,
                                                                                                                                                es_3_2_destruct_r,
                                                                                                                                                es_2_1_destruct_r}));
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_r = (& lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted <= 7'd0;
    else
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_emitted <= (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_r ? 7'd0 :
                                                               lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool2) : (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) > [(es_3_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (sc_0_4_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZad7_3_destruct,MyDTBool_Bool),
                                                                                                                               (gad8_3_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1adc_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2ada_3_destruct,Pointer_QTree_Bool),
                                                                                                                               (q2add_2_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted;
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_done;
  assign es_3_1_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[19:4],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[35:20],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[1]))};
  assign isZad7_3_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[2]));
  assign gad8_3_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[3]));
  assign q1adc_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[51:36],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[4]))};
  assign m2ada_3_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[67:52],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[5]))};
  assign q2add_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[83:68],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted[6]))};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_done = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted | ({q2add_2_destruct_d[0],
                                                                                                                       m2ada_3_destruct_d[0],
                                                                                                                       q1adc_2_destruct_d[0],
                                                                                                                       gad8_3_destruct_d[0],
                                                                                                                       isZad7_3_destruct_d[0],
                                                                                                                       sc_0_4_destruct_d[0],
                                                                                                                       es_3_1_destruct_d[0]} & {q2add_2_destruct_r,
                                                                                                                                                m2ada_3_destruct_r,
                                                                                                                                                q1adc_2_destruct_r,
                                                                                                                                                gad8_3_destruct_r,
                                                                                                                                                isZad7_3_destruct_r,
                                                                                                                                                sc_0_4_destruct_r,
                                                                                                                                                es_3_1_destruct_r}));
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_r = (& lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted <= 7'd0;
    else
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_emitted <= (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_r ? 7'd0 :
                                                               lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_done);
  
  /* destruct (Ty CTkron_kron_Bool_Bool_Bool,
          Dcon Lcall_kron_kron_Bool_Bool_Bool3) : (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) > [(sc_0_3_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                               (isZad7_2_destruct,MyDTBool_Bool),
                                                                                                                               (gad8_2_destruct,MyDTBool_Bool_Bool),
                                                                                                                               (q1adc_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (m2ada_2_destruct,Pointer_QTree_Bool),
                                                                                                                               (q2add_1_destruct,Pointer_QTree_Bool),
                                                                                                                               (q3ade_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted;
  logic [6:0] lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_done;
  assign sc_0_3_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[19:4],
                              (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[0]))};
  assign isZad7_2_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[1]));
  assign gad8_2_destruct_d = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[2]));
  assign q1adc_1_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[35:20],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[3]))};
  assign m2ada_2_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[51:36],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[4]))};
  assign q2add_1_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[67:52],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[5]))};
  assign q3ade_1_destruct_d = {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[83:68],
                               (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d[0] && (! lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted[6]))};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_done = (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted | ({q3ade_1_destruct_d[0],
                                                                                                                       q2add_1_destruct_d[0],
                                                                                                                       m2ada_2_destruct_d[0],
                                                                                                                       q1adc_1_destruct_d[0],
                                                                                                                       gad8_2_destruct_d[0],
                                                                                                                       isZad7_2_destruct_d[0],
                                                                                                                       sc_0_3_destruct_d[0]} & {q3ade_1_destruct_r,
                                                                                                                                                q2add_1_destruct_r,
                                                                                                                                                m2ada_2_destruct_r,
                                                                                                                                                q1adc_1_destruct_r,
                                                                                                                                                gad8_2_destruct_r,
                                                                                                                                                isZad7_2_destruct_r,
                                                                                                                                                sc_0_3_destruct_r}));
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_r = (& lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted <= 7'd0;
    else
      lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_emitted <= (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_r ? 7'd0 :
                                                               lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_done);
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet24_2,CTkron_kron_Bool_Bool_Bool) (lizzieLet24_1,CTkron_kron_Bool_Bool_Bool) > [(_19,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool)] */
  logic [4:0] lizzieLet24_1_onehotd;
  always_comb
    if ((lizzieLet24_2_d[0] && lizzieLet24_1_d[0]))
      unique case (lizzieLet24_2_d[3:1])
        3'd0: lizzieLet24_1_onehotd = 5'd1;
        3'd1: lizzieLet24_1_onehotd = 5'd2;
        3'd2: lizzieLet24_1_onehotd = 5'd4;
        3'd3: lizzieLet24_1_onehotd = 5'd8;
        3'd4: lizzieLet24_1_onehotd = 5'd16;
        default: lizzieLet24_1_onehotd = 5'd0;
      endcase
    else lizzieLet24_1_onehotd = 5'd0;
  assign _19_d = {lizzieLet24_1_d[83:1], lizzieLet24_1_onehotd[0]};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_d = {lizzieLet24_1_d[83:1],
                                                           lizzieLet24_1_onehotd[1]};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_d = {lizzieLet24_1_d[83:1],
                                                           lizzieLet24_1_onehotd[2]};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_d = {lizzieLet24_1_d[83:1],
                                                           lizzieLet24_1_onehotd[3]};
  assign lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_d = {lizzieLet24_1_d[83:1],
                                                           lizzieLet24_1_onehotd[4]};
  assign lizzieLet24_1_r = (| (lizzieLet24_1_onehotd & {lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                        lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                        lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                        lizzieLet24_1Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                        _19_r}));
  assign lizzieLet24_2_r = lizzieLet24_1_r;
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty Go) : (lizzieLet24_3,CTkron_kron_Bool_Bool_Bool) (go_13_goMux_data,Go) > [(_18,Go),
                                                                                    (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3,Go),
                                                                                    (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2,Go),
                                                                                    (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1,Go),
                                                                                    (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0,Go)] */
  logic [4:0] go_13_goMux_data_onehotd;
  always_comb
    if ((lizzieLet24_3_d[0] && go_13_goMux_data_d[0]))
      unique case (lizzieLet24_3_d[3:1])
        3'd0: go_13_goMux_data_onehotd = 5'd1;
        3'd1: go_13_goMux_data_onehotd = 5'd2;
        3'd2: go_13_goMux_data_onehotd = 5'd4;
        3'd3: go_13_goMux_data_onehotd = 5'd8;
        3'd4: go_13_goMux_data_onehotd = 5'd16;
        default: go_13_goMux_data_onehotd = 5'd0;
      endcase
    else go_13_goMux_data_onehotd = 5'd0;
  assign _18_d = go_13_goMux_data_onehotd[0];
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_d = go_13_goMux_data_onehotd[1];
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_d = go_13_goMux_data_onehotd[2];
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_d = go_13_goMux_data_onehotd[3];
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_d = go_13_goMux_data_onehotd[4];
  assign go_13_goMux_data_r = (| (go_13_goMux_data_onehotd & {lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                              lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                              lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                              lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                              _18_r}));
  assign lizzieLet24_3_r = go_13_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0,Go) > (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_r = ((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d[0]) || lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_r)
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_d;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r = (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d = (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0] ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf :
                                                                    lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r && lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r) && (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0])))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1,Go) > (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_r = ((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d[0]) || lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_r)
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_d;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r = (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_d = (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0] ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf :
                                                                    lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r && lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_1_argbuf_r) && (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0])))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2,Go) > (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_r = ((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d[0]) || lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_r)
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_d;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r = (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_d = (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0] ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf :
                                                                    lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r && lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_1_argbuf_r) && (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0])))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3,Go) > (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf,Go) */
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  logic lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_r = ((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d[0]) || lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= 1'd0;
    else
      if (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_r)
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_d;
  Go_t lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf;
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r = (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]);
  assign lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_d = (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0] ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf :
                                                                    lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r && lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_1_argbuf_r) && (! lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0])))
        lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  
  /* demux (Ty CTkron_kron_Bool_Bool_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet24_4,CTkron_kron_Bool_Bool_Bool) (srtarg_0_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                                                                                      (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet24_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet24_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d = {srtarg_0_goMux_mux_d[16:1],
                                                         srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_d = {srtarg_0_goMux_mux_d[16:1],
                                                           srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_r,
                                                                  lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_r,
                                                                  lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_r,
                                                                  lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_r,
                                                                  lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_r}));
  assign lizzieLet24_4_r = srtarg_0_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0,Pointer_QTree_Bool),
                          (es_1_2_destruct,Pointer_QTree_Bool),
                          (es_2_2_destruct,Pointer_QTree_Bool),
                          (es_3_3_destruct,Pointer_QTree_Bool)] > (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) */
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d = QNode_Bool_dc((& {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_d[0],
                                                                                                                es_1_2_destruct_d[0],
                                                                                                                es_2_2_destruct_d[0],
                                                                                                                es_3_3_destruct_d[0]}), lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_d, es_1_2_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_r,
          es_1_2_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool,QTree_Bool) > (lizzieLet28_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r = ((! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d[0]) || lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d <= {66'd0,
                                                                                                     1'd0};
    else
      if (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_r)
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_d;
  QTree_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_r = (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0]);
  assign lizzieLet28_1_argbuf_d = (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0] ? lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf :
                                   lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                                       1'd0};
    else
      if ((lizzieLet28_1_argbuf_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0]))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= {66'd0,
                                                                                                         1'd0};
      else if (((! lizzieLet28_1_argbuf_r) && (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf[0])))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_buf <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool0_1es_1_2_1es_2_2_1es_3_3_1QNode_Bool_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool0) : [(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                               (es_2_1_destruct,Pointer_QTree_Bool),
                                               (es_3_2_destruct,Pointer_QTree_Bool),
                                               (sc_0_5_destruct,Pointer_CTkron_kron_Bool_Bool_Bool)] > (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d = Lcall_kron_kron_Bool_Bool_Bool0_dc((& {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_d[0],
                                                                                                                                                          es_2_1_destruct_d[0],
                                                                                                                                                          es_3_2_destruct_d[0],
                                                                                                                                                          sc_0_5_destruct_d[0]}), lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_d, es_2_1_destruct_d, es_3_2_destruct_d, sc_0_5_destruct_d);
  assign {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_r,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_5_destruct_r} = {4 {(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0,CTkron_kron_Bool_Bool_Bool) > (lizzieLet27_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r = ((! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d[0]) || lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= {83'd0,
                                                                                                                          1'd0};
    else
      if (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_r)
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_r = (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]);
  assign lizzieLet27_1_argbuf_d = (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0] ? lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf :
                                   lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= {83'd0,
                                                                                                                            1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0]))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= {83'd0,
                                                                                                                              1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf[0])))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_buf <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool1_1es_2_1_1es_3_2_1sc_0_5_1Lcall_kron_kron_Bool_Bool_Bool0_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool1) : [(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                               (es_3_1_destruct,Pointer_QTree_Bool),
                                               (sc_0_4_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (isZad7_3_1,MyDTBool_Bool),
                                               (gad8_3_1,MyDTBool_Bool_Bool),
                                               (q1adc_2_destruct,Pointer_QTree_Bool),
                                               (m2ada_3_1,Pointer_QTree_Bool)] > (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_d = Lcall_kron_kron_Bool_Bool_Bool1_dc((& {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_d[0],
                                                                                                                                                                                      es_3_1_destruct_d[0],
                                                                                                                                                                                      sc_0_4_destruct_d[0],
                                                                                                                                                                                      isZad7_3_1_d[0],
                                                                                                                                                                                      gad8_3_1_d[0],
                                                                                                                                                                                      q1adc_2_destruct_d[0],
                                                                                                                                                                                      m2ada_3_1_d[0]}), lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_d, es_3_1_destruct_d, sc_0_4_destruct_d, isZad7_3_1_d, gad8_3_1_d, q1adc_2_destruct_d, m2ada_3_1_d);
  assign {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_r,
          es_3_1_destruct_r,
          sc_0_4_destruct_r,
          isZad7_3_1_r,
          gad8_3_1_r,
          q1adc_2_destruct_r,
          m2ada_3_1_r} = {7 {(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1,CTkron_kron_Bool_Bool_Bool) > (lizzieLet26_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_r = ((! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d[0]) || lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= {83'd0,
                                                                                                                                                      1'd0};
    else
      if (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_r)
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_r = (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]);
  assign lizzieLet26_1_argbuf_d = (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0] ? lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf :
                                   lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= {83'd0,
                                                                                                                                                        1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0]))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= {83'd0,
                                                                                                                                                          1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf[0])))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_buf <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool2_1es_3_1_1sc_0_4_1isZad7_3_1gad8_3_1q1adc_2_1m2ada_3_1Lcall_kron_kron_Bool_Bool_Bool1_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool2) : [(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                               (sc_0_3_destruct,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (isZad7_2_1,MyDTBool_Bool),
                                               (gad8_2_1,MyDTBool_Bool_Bool),
                                               (q1adc_1_destruct,Pointer_QTree_Bool),
                                               (m2ada_2_1,Pointer_QTree_Bool),
                                               (q2add_1_destruct,Pointer_QTree_Bool)] > (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_d = Lcall_kron_kron_Bool_Bool_Bool2_dc((& {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_d[0],
                                                                                                                                                                                       sc_0_3_destruct_d[0],
                                                                                                                                                                                       isZad7_2_1_d[0],
                                                                                                                                                                                       gad8_2_1_d[0],
                                                                                                                                                                                       q1adc_1_destruct_d[0],
                                                                                                                                                                                       m2ada_2_1_d[0],
                                                                                                                                                                                       q2add_1_destruct_d[0]}), lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_d, sc_0_3_destruct_d, isZad7_2_1_d, gad8_2_1_d, q1adc_1_destruct_d, m2ada_2_1_d, q2add_1_destruct_d);
  assign {lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_r,
          sc_0_3_destruct_r,
          isZad7_2_1_r,
          gad8_2_1_r,
          q1adc_1_destruct_r,
          m2ada_2_1_r,
          q2add_1_destruct_r} = {7 {(lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2,CTkron_kron_Bool_Bool_Bool) > (lizzieLet25_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  logic lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_r = ((! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d[0]) || lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= {83'd0,
                                                                                                                                                       1'd0};
    else
      if (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_r)
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf;
  assign lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_r = (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]);
  assign lizzieLet25_1_argbuf_d = (lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0] ? lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf :
                                   lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= {83'd0,
                                                                                                                                                         1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0]))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= {83'd0,
                                                                                                                                                           1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf[0])))
        lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_buf <= lizzieLet24_4Lcall_kron_kron_Bool_Bool_Bool3_1sc_0_3_1isZad7_2_1gad8_2_1q1adc_1_1m2ada_2_1q2add_1_1Lcall_kron_kron_Bool_Bool_Bool2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                                  (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted;
  logic [1:0] lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_done;
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d = {lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d[16:1],
                                                                              (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d[0] && (! lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted[0]))};
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d = {lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d[16:1],
                                                                              (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_d[0] && (! lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted[1]))};
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_done = (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted | ({lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d[0],
                                                                                                                   lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r,
                                                                                                                                                                                            lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_r = (& lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted <= 2'd0;
    else
      lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_emitted <= (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_r ? 2'd0 :
                                                             lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_done);
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_kron_kron_Bool_Bool_Bool_goConst,Go) */
  assign call_kron_kron_Bool_Bool_Bool_goConst_d = lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r = call_kron_kron_Bool_Bool_Bool_goConst_r;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (kron_kron_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r = ((! lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                                    1'd0};
    else
      if (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r)
        lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Bool_t lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign kron_kron_Bool_Bool_Bool_resbuf_d = (lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf :
                                              lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                      1'd0};
    else
      if ((kron_kron_Bool_Bool_Bool_resbuf_r && lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                        1'd0};
      else if (((! kron_kron_Bool_Bool_Bool_resbuf_r) && (! lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet24_4Lkron_kron_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* destruct (Ty CTmain_map'_Bool_Nat,
          Dcon Lcall_main_map'_Bool_Nat0) : (lizzieLet29_1Lcall_main_map'_Bool_Nat0,CTmain_map'_Bool_Nat) > [(es_2_3_destruct,Pointer_QTree_Nat),
                                                                                                             (es_3_5_destruct,Pointer_QTree_Nat),
                                                                                                             (es_4_3_destruct,Pointer_QTree_Nat),
                                                                                                             (sc_0_10_destruct,Pointer_CTmain_map'_Bool_Nat)] */
  logic [3:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted ;
  logic [3:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat0_done ;
  assign es_2_3_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [19:4],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted [0]))};
  assign es_3_5_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [35:20],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted [1]))};
  assign es_4_3_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [51:36],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [67:52],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted [3]))};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat0_done  = (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted  | ({sc_0_10_destruct_d[0],
                                                                                                               es_4_3_destruct_d[0],
                                                                                                               es_3_5_destruct_d[0],
                                                                                                               es_2_3_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                                        es_4_3_destruct_r,
                                                                                                                                        es_3_5_destruct_r,
                                                                                                                                        es_2_3_destruct_r}));
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat0_r  = (& \lizzieLet29_1Lcall_main_map'_Bool_Nat0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted  <= 4'd0;
    else
      \lizzieLet29_1Lcall_main_map'_Bool_Nat0_emitted  <= (\lizzieLet29_1Lcall_main_map'_Bool_Nat0_r  ? 4'd0 :
                                                           \lizzieLet29_1Lcall_main_map'_Bool_Nat0_done );
  
  /* destruct (Ty CTmain_map'_Bool_Nat,
          Dcon Lcall_main_map'_Bool_Nat1) : (lizzieLet29_1Lcall_main_map'_Bool_Nat1,CTmain_map'_Bool_Nat) > [(es_3_4_destruct,Pointer_QTree_Nat),
                                                                                                             (es_4_2_destruct,Pointer_QTree_Nat),
                                                                                                             (sc_0_9_destruct,Pointer_CTmain_map'_Bool_Nat),
                                                                                                             (isZacQ_4_destruct,MyDTNat_Bool),
                                                                                                             (gacR_4_destruct,MyDTBool_Nat),
                                                                                                             (q1acU_3_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted ;
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat1_done ;
  assign es_3_4_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [19:4],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [0]))};
  assign es_4_2_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [35:20],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [51:36],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [2]))};
  assign isZacQ_4_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [3]));
  assign gacR_4_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [4]));
  assign q1acU_3_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [67:52],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted [5]))};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat1_done  = (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted  | ({q1acU_3_destruct_d[0],
                                                                                                               gacR_4_destruct_d[0],
                                                                                                               isZacQ_4_destruct_d[0],
                                                                                                               sc_0_9_destruct_d[0],
                                                                                                               es_4_2_destruct_d[0],
                                                                                                               es_3_4_destruct_d[0]} & {q1acU_3_destruct_r,
                                                                                                                                        gacR_4_destruct_r,
                                                                                                                                        isZacQ_4_destruct_r,
                                                                                                                                        sc_0_9_destruct_r,
                                                                                                                                        es_4_2_destruct_r,
                                                                                                                                        es_3_4_destruct_r}));
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat1_r  = (& \lizzieLet29_1Lcall_main_map'_Bool_Nat1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted  <= 6'd0;
    else
      \lizzieLet29_1Lcall_main_map'_Bool_Nat1_emitted  <= (\lizzieLet29_1Lcall_main_map'_Bool_Nat1_r  ? 6'd0 :
                                                           \lizzieLet29_1Lcall_main_map'_Bool_Nat1_done );
  
  /* destruct (Ty CTmain_map'_Bool_Nat,
          Dcon Lcall_main_map'_Bool_Nat2) : (lizzieLet29_1Lcall_main_map'_Bool_Nat2,CTmain_map'_Bool_Nat) > [(es_4_1_destruct,Pointer_QTree_Nat),
                                                                                                             (sc_0_8_destruct,Pointer_CTmain_map'_Bool_Nat),
                                                                                                             (isZacQ_3_destruct,MyDTNat_Bool),
                                                                                                             (gacR_3_destruct,MyDTBool_Nat),
                                                                                                             (q1acU_2_destruct,Pointer_QTree_Bool),
                                                                                                             (q2acV_2_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted ;
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat2_done ;
  assign es_4_1_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [19:4],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [35:20],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [1]))};
  assign isZacQ_3_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [2]));
  assign gacR_3_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [3]));
  assign q1acU_2_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [51:36],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [4]))};
  assign q2acV_2_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [67:52],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted [5]))};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat2_done  = (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted  | ({q2acV_2_destruct_d[0],
                                                                                                               q1acU_2_destruct_d[0],
                                                                                                               gacR_3_destruct_d[0],
                                                                                                               isZacQ_3_destruct_d[0],
                                                                                                               sc_0_8_destruct_d[0],
                                                                                                               es_4_1_destruct_d[0]} & {q2acV_2_destruct_r,
                                                                                                                                        q1acU_2_destruct_r,
                                                                                                                                        gacR_3_destruct_r,
                                                                                                                                        isZacQ_3_destruct_r,
                                                                                                                                        sc_0_8_destruct_r,
                                                                                                                                        es_4_1_destruct_r}));
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat2_r  = (& \lizzieLet29_1Lcall_main_map'_Bool_Nat2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted  <= 6'd0;
    else
      \lizzieLet29_1Lcall_main_map'_Bool_Nat2_emitted  <= (\lizzieLet29_1Lcall_main_map'_Bool_Nat2_r  ? 6'd0 :
                                                           \lizzieLet29_1Lcall_main_map'_Bool_Nat2_done );
  
  /* destruct (Ty CTmain_map'_Bool_Nat,
          Dcon Lcall_main_map'_Bool_Nat3) : (lizzieLet29_1Lcall_main_map'_Bool_Nat3,CTmain_map'_Bool_Nat) > [(sc_0_7_destruct,Pointer_CTmain_map'_Bool_Nat),
                                                                                                             (isZacQ_2_destruct,MyDTNat_Bool),
                                                                                                             (gacR_2_destruct,MyDTBool_Nat),
                                                                                                             (q1acU_1_destruct,Pointer_QTree_Bool),
                                                                                                             (q2acV_1_destruct,Pointer_QTree_Bool),
                                                                                                             (q3acW_1_destruct,Pointer_QTree_Bool)] */
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted ;
  logic [5:0] \lizzieLet29_1Lcall_main_map'_Bool_Nat3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [19:4],
                              (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [0]))};
  assign isZacQ_2_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [1]));
  assign gacR_2_destruct_d = (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [2]));
  assign q1acU_1_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [35:20],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [3]))};
  assign q2acV_1_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [51:36],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [4]))};
  assign q3acW_1_destruct_d = {\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [67:52],
                               (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_d [0] && (! \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted [5]))};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat3_done  = (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted  | ({q3acW_1_destruct_d[0],
                                                                                                               q2acV_1_destruct_d[0],
                                                                                                               q1acU_1_destruct_d[0],
                                                                                                               gacR_2_destruct_d[0],
                                                                                                               isZacQ_2_destruct_d[0],
                                                                                                               sc_0_7_destruct_d[0]} & {q3acW_1_destruct_r,
                                                                                                                                        q2acV_1_destruct_r,
                                                                                                                                        q1acU_1_destruct_r,
                                                                                                                                        gacR_2_destruct_r,
                                                                                                                                        isZacQ_2_destruct_r,
                                                                                                                                        sc_0_7_destruct_r}));
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat3_r  = (& \lizzieLet29_1Lcall_main_map'_Bool_Nat3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted  <= 6'd0;
    else
      \lizzieLet29_1Lcall_main_map'_Bool_Nat3_emitted  <= (\lizzieLet29_1Lcall_main_map'_Bool_Nat3_r  ? 6'd0 :
                                                           \lizzieLet29_1Lcall_main_map'_Bool_Nat3_done );
  
  /* demux (Ty CTmain_map'_Bool_Nat,
       Ty CTmain_map'_Bool_Nat) : (lizzieLet29_2,CTmain_map'_Bool_Nat) (lizzieLet29_1,CTmain_map'_Bool_Nat) > [(_17,CTmain_map'_Bool_Nat),
                                                                                                               (lizzieLet29_1Lcall_main_map'_Bool_Nat3,CTmain_map'_Bool_Nat),
                                                                                                               (lizzieLet29_1Lcall_main_map'_Bool_Nat2,CTmain_map'_Bool_Nat),
                                                                                                               (lizzieLet29_1Lcall_main_map'_Bool_Nat1,CTmain_map'_Bool_Nat),
                                                                                                               (lizzieLet29_1Lcall_main_map'_Bool_Nat0,CTmain_map'_Bool_Nat)] */
  logic [4:0] lizzieLet29_1_onehotd;
  always_comb
    if ((lizzieLet29_2_d[0] && lizzieLet29_1_d[0]))
      unique case (lizzieLet29_2_d[3:1])
        3'd0: lizzieLet29_1_onehotd = 5'd1;
        3'd1: lizzieLet29_1_onehotd = 5'd2;
        3'd2: lizzieLet29_1_onehotd = 5'd4;
        3'd3: lizzieLet29_1_onehotd = 5'd8;
        3'd4: lizzieLet29_1_onehotd = 5'd16;
        default: lizzieLet29_1_onehotd = 5'd0;
      endcase
    else lizzieLet29_1_onehotd = 5'd0;
  assign _17_d = {lizzieLet29_1_d[67:1], lizzieLet29_1_onehotd[0]};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat3_d  = {lizzieLet29_1_d[67:1],
                                                       lizzieLet29_1_onehotd[1]};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat2_d  = {lizzieLet29_1_d[67:1],
                                                       lizzieLet29_1_onehotd[2]};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat1_d  = {lizzieLet29_1_d[67:1],
                                                       lizzieLet29_1_onehotd[3]};
  assign \lizzieLet29_1Lcall_main_map'_Bool_Nat0_d  = {lizzieLet29_1_d[67:1],
                                                       lizzieLet29_1_onehotd[4]};
  assign lizzieLet29_1_r = (| (lizzieLet29_1_onehotd & {\lizzieLet29_1Lcall_main_map'_Bool_Nat0_r ,
                                                        \lizzieLet29_1Lcall_main_map'_Bool_Nat1_r ,
                                                        \lizzieLet29_1Lcall_main_map'_Bool_Nat2_r ,
                                                        \lizzieLet29_1Lcall_main_map'_Bool_Nat3_r ,
                                                        _17_r}));
  assign lizzieLet29_2_r = lizzieLet29_1_r;
  
  /* demux (Ty CTmain_map'_Bool_Nat,
       Ty Go) : (lizzieLet29_3,CTmain_map'_Bool_Nat) (go_14_goMux_data,Go) > [(_16,Go),
                                                                              (lizzieLet29_3Lcall_main_map'_Bool_Nat3,Go),
                                                                              (lizzieLet29_3Lcall_main_map'_Bool_Nat2,Go),
                                                                              (lizzieLet29_3Lcall_main_map'_Bool_Nat1,Go),
                                                                              (lizzieLet29_3Lcall_main_map'_Bool_Nat0,Go)] */
  logic [4:0] go_14_goMux_data_onehotd;
  always_comb
    if ((lizzieLet29_3_d[0] && go_14_goMux_data_d[0]))
      unique case (lizzieLet29_3_d[3:1])
        3'd0: go_14_goMux_data_onehotd = 5'd1;
        3'd1: go_14_goMux_data_onehotd = 5'd2;
        3'd2: go_14_goMux_data_onehotd = 5'd4;
        3'd3: go_14_goMux_data_onehotd = 5'd8;
        3'd4: go_14_goMux_data_onehotd = 5'd16;
        default: go_14_goMux_data_onehotd = 5'd0;
      endcase
    else go_14_goMux_data_onehotd = 5'd0;
  assign _16_d = go_14_goMux_data_onehotd[0];
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat3_d  = go_14_goMux_data_onehotd[1];
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat2_d  = go_14_goMux_data_onehotd[2];
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat1_d  = go_14_goMux_data_onehotd[3];
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat0_d  = go_14_goMux_data_onehotd[4];
  assign go_14_goMux_data_r = (| (go_14_goMux_data_onehotd & {\lizzieLet29_3Lcall_main_map'_Bool_Nat0_r ,
                                                              \lizzieLet29_3Lcall_main_map'_Bool_Nat1_r ,
                                                              \lizzieLet29_3Lcall_main_map'_Bool_Nat2_r ,
                                                              \lizzieLet29_3Lcall_main_map'_Bool_Nat3_r ,
                                                              _16_r}));
  assign lizzieLet29_3_r = go_14_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_main_map'_Bool_Nat0,Go) > (lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf,Go) */
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_r ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat0_r  = ((! \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d [0]) || \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet29_3Lcall_main_map'_Bool_Nat0_r )
        \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat0_d ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_r  = (! \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf [0]);
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_d  = (\lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf [0] ? \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf  :
                                                                \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_r  && \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf [0]))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_r ) && (! \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf [0])))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_buf  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_main_map'_Bool_Nat1,Go) > (lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf,Go) */
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_r ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat1_r  = ((! \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d [0]) || \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet29_3Lcall_main_map'_Bool_Nat1_r )
        \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat1_d ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_r  = (! \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf [0]);
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_d  = (\lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf [0] ? \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf  :
                                                                \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_r  && \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf [0]))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet29_3Lcall_main_map'_Bool_Nat1_1_argbuf_r ) && (! \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf [0])))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_buf  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_main_map'_Bool_Nat2,Go) > (lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf,Go) */
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_r ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat2_r  = ((! \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d [0]) || \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet29_3Lcall_main_map'_Bool_Nat2_r )
        \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat2_d ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_r  = (! \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf [0]);
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_d  = (\lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf [0] ? \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf  :
                                                                \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_r  && \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf [0]))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet29_3Lcall_main_map'_Bool_Nat2_1_argbuf_r ) && (! \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf [0])))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_buf  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet29_3Lcall_main_map'_Bool_Nat3,Go) > (lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf,Go) */
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d ;
  logic \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_r ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat3_r  = ((! \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d [0]) || \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet29_3Lcall_main_map'_Bool_Nat3_r )
        \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat3_d ;
  Go_t \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf ;
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_r  = (! \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf [0]);
  assign \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_d  = (\lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf [0] ? \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf  :
                                                                \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_r  && \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf [0]))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet29_3Lcall_main_map'_Bool_Nat3_1_argbuf_r ) && (! \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf [0])))
        \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_buf  <= \lizzieLet29_3Lcall_main_map'_Bool_Nat3_bufchan_d ;
  
  /* demux (Ty CTmain_map'_Bool_Nat,
       Ty Pointer_QTree_Nat) : (lizzieLet29_4,CTmain_map'_Bool_Nat) (srtarg_0_1_goMux_mux,Pointer_QTree_Nat) > [(lizzieLet29_4Lmain_map'_Bool_Natsbos,Pointer_QTree_Nat),
                                                                                                                (lizzieLet29_4Lcall_main_map'_Bool_Nat3,Pointer_QTree_Nat),
                                                                                                                (lizzieLet29_4Lcall_main_map'_Bool_Nat2,Pointer_QTree_Nat),
                                                                                                                (lizzieLet29_4Lcall_main_map'_Bool_Nat1,Pointer_QTree_Nat),
                                                                                                                (lizzieLet29_4Lcall_main_map'_Bool_Nat0,Pointer_QTree_Nat)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet29_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet29_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                     srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                       srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                       srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                       srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                       srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet29_4Lcall_main_map'_Bool_Nat0_r ,
                                                                      \lizzieLet29_4Lcall_main_map'_Bool_Nat1_r ,
                                                                      \lizzieLet29_4Lcall_main_map'_Bool_Nat2_r ,
                                                                      \lizzieLet29_4Lcall_main_map'_Bool_Nat3_r ,
                                                                      \lizzieLet29_4Lmain_map'_Bool_Natsbos_r }));
  assign lizzieLet29_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Nat,
      Dcon QNode_Nat) : [(lizzieLet29_4Lcall_main_map'_Bool_Nat0,Pointer_QTree_Nat),
                         (es_2_3_destruct,Pointer_QTree_Nat),
                         (es_3_5_destruct,Pointer_QTree_Nat),
                         (es_4_3_destruct,Pointer_QTree_Nat)] > (lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat,QTree_Nat) */
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_d  = QNode_Nat_dc((& {\lizzieLet29_4Lcall_main_map'_Bool_Nat0_d [0],
                                                                                                          es_2_3_destruct_d[0],
                                                                                                          es_3_5_destruct_d[0],
                                                                                                          es_4_3_destruct_d[0]}), \lizzieLet29_4Lcall_main_map'_Bool_Nat0_d , es_2_3_destruct_d, es_3_5_destruct_d, es_4_3_destruct_d);
  assign {\lizzieLet29_4Lcall_main_map'_Bool_Nat0_r ,
          es_2_3_destruct_r,
          es_3_5_destruct_r,
          es_4_3_destruct_r} = {4 {(\lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_r  && \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_d [0])}};
  
  /* buf (Ty QTree_Nat) : (lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat,QTree_Nat) > (lizzieLet33_1_argbuf,QTree_Nat) */
  QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_r ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_r  = ((! \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d [0]) || \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d  <= {66'd0,
                                                                                                1'd0};
    else
      if (\lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_r )
        \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_d ;
  QTree_Nat_t \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_r  = (! \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf [0]);
  assign lizzieLet33_1_argbuf_d = (\lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf [0] ? \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf  :
                                   \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf  <= {66'd0,
                                                                                                  1'd0};
    else
      if ((lizzieLet33_1_argbuf_r && \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf [0]))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf  <= {66'd0,
                                                                                                    1'd0};
      else if (((! lizzieLet33_1_argbuf_r) && (! \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf [0])))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_buf  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat0_1es_2_3_1es_3_5_1es_4_3_1QNode_Nat_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Bool_Nat,
      Dcon Lcall_main_map'_Bool_Nat0) : [(lizzieLet29_4Lcall_main_map'_Bool_Nat1,Pointer_QTree_Nat),
                                         (es_3_4_destruct,Pointer_QTree_Nat),
                                         (es_4_2_destruct,Pointer_QTree_Nat),
                                         (sc_0_9_destruct,Pointer_CTmain_map'_Bool_Nat)] > (lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0,CTmain_map'_Bool_Nat) */
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_d  = \Lcall_main_map'_Bool_Nat0_dc ((& {\lizzieLet29_4Lcall_main_map'_Bool_Nat1_d [0],
                                                                                                                                            es_3_4_destruct_d[0],
                                                                                                                                            es_4_2_destruct_d[0],
                                                                                                                                            sc_0_9_destruct_d[0]}), \lizzieLet29_4Lcall_main_map'_Bool_Nat1_d , es_3_4_destruct_d, es_4_2_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet29_4Lcall_main_map'_Bool_Nat1_r ,
          es_3_4_destruct_r,
          es_4_2_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_r  && \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_d [0])}};
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0,CTmain_map'_Bool_Nat) > (lizzieLet32_1_argbuf,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_r ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_r  = ((! \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d [0]) || \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d  <= {67'd0,
                                                                                                                1'd0};
    else
      if (\lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_r )
        \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_d ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_r  = (! \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf [0]);
  assign lizzieLet32_1_argbuf_d = (\lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf [0] ? \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf  :
                                   \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf  <= {67'd0,
                                                                                                                  1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf [0]))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf  <= {67'd0,
                                                                                                                    1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf [0])))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_buf  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat1_1es_3_4_1es_4_2_1sc_0_9_1Lcall_main_map'_Bool_Nat0_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Bool_Nat,
      Dcon Lcall_main_map'_Bool_Nat1) : [(lizzieLet29_4Lcall_main_map'_Bool_Nat2,Pointer_QTree_Nat),
                                         (es_4_1_destruct,Pointer_QTree_Nat),
                                         (sc_0_8_destruct,Pointer_CTmain_map'_Bool_Nat),
                                         (isZacQ_3_1,MyDTNat_Bool),
                                         (gacR_3_1,MyDTBool_Nat),
                                         (q1acU_2_destruct,Pointer_QTree_Bool)] > (lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1,CTmain_map'_Bool_Nat) */
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_d  = \Lcall_main_map'_Bool_Nat1_dc ((& {\lizzieLet29_4Lcall_main_map'_Bool_Nat2_d [0],
                                                                                                                                                               es_4_1_destruct_d[0],
                                                                                                                                                               sc_0_8_destruct_d[0],
                                                                                                                                                               isZacQ_3_1_d[0],
                                                                                                                                                               gacR_3_1_d[0],
                                                                                                                                                               q1acU_2_destruct_d[0]}), \lizzieLet29_4Lcall_main_map'_Bool_Nat2_d , es_4_1_destruct_d, sc_0_8_destruct_d, isZacQ_3_1_d, gacR_3_1_d, q1acU_2_destruct_d);
  assign {\lizzieLet29_4Lcall_main_map'_Bool_Nat2_r ,
          es_4_1_destruct_r,
          sc_0_8_destruct_r,
          isZacQ_3_1_r,
          gacR_3_1_r,
          q1acU_2_destruct_r} = {6 {(\lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_r  && \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_d [0])}};
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1,CTmain_map'_Bool_Nat) > (lizzieLet31_1_argbuf,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_r ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_r  = ((! \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d [0]) || \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d  <= {67'd0,
                                                                                                                                   1'd0};
    else
      if (\lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_r )
        \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_d ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_r  = (! \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf [0]);
  assign lizzieLet31_1_argbuf_d = (\lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf [0] ? \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf  :
                                   \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf  <= {67'd0,
                                                                                                                                     1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf [0]))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf  <= {67'd0,
                                                                                                                                       1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf [0])))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_buf  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat2_1es_4_1_1sc_0_8_1isZacQ_3_1gacR_3_1q1acU_2_1Lcall_main_map'_Bool_Nat1_bufchan_d ;
  
  /* dcon (Ty CTmain_map'_Bool_Nat,
      Dcon Lcall_main_map'_Bool_Nat2) : [(lizzieLet29_4Lcall_main_map'_Bool_Nat3,Pointer_QTree_Nat),
                                         (sc_0_7_destruct,Pointer_CTmain_map'_Bool_Nat),
                                         (isZacQ_2_1,MyDTNat_Bool),
                                         (gacR_2_1,MyDTBool_Nat),
                                         (q1acU_1_destruct,Pointer_QTree_Bool),
                                         (q2acV_1_destruct,Pointer_QTree_Bool)] > (lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2,CTmain_map'_Bool_Nat) */
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_d  = \Lcall_main_map'_Bool_Nat2_dc ((& {\lizzieLet29_4Lcall_main_map'_Bool_Nat3_d [0],
                                                                                                                                                                sc_0_7_destruct_d[0],
                                                                                                                                                                isZacQ_2_1_d[0],
                                                                                                                                                                gacR_2_1_d[0],
                                                                                                                                                                q1acU_1_destruct_d[0],
                                                                                                                                                                q2acV_1_destruct_d[0]}), \lizzieLet29_4Lcall_main_map'_Bool_Nat3_d , sc_0_7_destruct_d, isZacQ_2_1_d, gacR_2_1_d, q1acU_1_destruct_d, q2acV_1_destruct_d);
  assign {\lizzieLet29_4Lcall_main_map'_Bool_Nat3_r ,
          sc_0_7_destruct_r,
          isZacQ_2_1_r,
          gacR_2_1_r,
          q1acU_1_destruct_r,
          q2acV_1_destruct_r} = {6 {(\lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_r  && \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_d [0])}};
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2,CTmain_map'_Bool_Nat) > (lizzieLet30_1_argbuf,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d ;
  logic \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_r ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_r  = ((! \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d [0]) || \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d  <= {67'd0,
                                                                                                                                    1'd0};
    else
      if (\lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_r )
        \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_d ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf ;
  assign \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_r  = (! \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf [0]);
  assign lizzieLet30_1_argbuf_d = (\lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf [0] ? \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf  :
                                   \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf  <= {67'd0,
                                                                                                                                      1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf [0]))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf  <= {67'd0,
                                                                                                                                        1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf [0])))
        \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_buf  <= \lizzieLet29_4Lcall_main_map'_Bool_Nat3_1sc_0_7_1isZacQ_2_1gacR_2_1q1acU_1_1q2acV_1_1Lcall_main_map'_Bool_Nat2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Nat) : (lizzieLet29_4Lmain_map'_Bool_Natsbos,Pointer_QTree_Nat) > [(lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1,Pointer_QTree_Nat),
                                                                                          (lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2,Pointer_QTree_Nat)] */
  logic [1:0] \lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted ;
  logic [1:0] \lizzieLet29_4Lmain_map'_Bool_Natsbos_done ;
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_d  = {\lizzieLet29_4Lmain_map'_Bool_Natsbos_d [16:1],
                                                                          (\lizzieLet29_4Lmain_map'_Bool_Natsbos_d [0] && (! \lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted [0]))};
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_d  = {\lizzieLet29_4Lmain_map'_Bool_Natsbos_d [16:1],
                                                                          (\lizzieLet29_4Lmain_map'_Bool_Natsbos_d [0] && (! \lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted [1]))};
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_done  = (\lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted  | ({\lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_d [0],
                                                                                                           \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_r  = (& \lizzieLet29_4Lmain_map'_Bool_Natsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted  <= 2'd0;
    else
      \lizzieLet29_4Lmain_map'_Bool_Natsbos_emitted  <= (\lizzieLet29_4Lmain_map'_Bool_Natsbos_r  ? 2'd0 :
                                                         \lizzieLet29_4Lmain_map'_Bool_Natsbos_done );
  
  /* togo (Ty Pointer_QTree_Nat) : (lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1,Pointer_QTree_Nat) > (call_main_map'_Bool_Nat_goConst,Go) */
  assign \call_main_map'_Bool_Nat_goConst_d  = \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_1_r  = \call_main_map'_Bool_Nat_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Nat) : (lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2,Pointer_QTree_Nat) > (main_map'_Bool_Nat_resbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_r )
        \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Nat_t \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \main_map'_Bool_Nat_resbuf_d  = (\lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf  :
                                          \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((\main_map'_Bool_Nat_resbuf_r  && \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! \main_map'_Bool_Nat_resbuf_r ) && (! \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet29_4Lmain_map'_Bool_Natsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet2_1QNode_Bool,QTree_Bool) > [(q1adc_destruct,Pointer_QTree_Bool),
                                                                    (q2add_destruct,Pointer_QTree_Bool),
                                                                    (q3ade_destruct,Pointer_QTree_Bool),
                                                                    (q4adf_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet2_1QNode_Bool_emitted;
  logic [3:0] lizzieLet2_1QNode_Bool_done;
  assign q1adc_destruct_d = {lizzieLet2_1QNode_Bool_d[18:3],
                             (lizzieLet2_1QNode_Bool_d[0] && (! lizzieLet2_1QNode_Bool_emitted[0]))};
  assign q2add_destruct_d = {lizzieLet2_1QNode_Bool_d[34:19],
                             (lizzieLet2_1QNode_Bool_d[0] && (! lizzieLet2_1QNode_Bool_emitted[1]))};
  assign q3ade_destruct_d = {lizzieLet2_1QNode_Bool_d[50:35],
                             (lizzieLet2_1QNode_Bool_d[0] && (! lizzieLet2_1QNode_Bool_emitted[2]))};
  assign q4adf_destruct_d = {lizzieLet2_1QNode_Bool_d[66:51],
                             (lizzieLet2_1QNode_Bool_d[0] && (! lizzieLet2_1QNode_Bool_emitted[3]))};
  assign lizzieLet2_1QNode_Bool_done = (lizzieLet2_1QNode_Bool_emitted | ({q4adf_destruct_d[0],
                                                                           q3ade_destruct_d[0],
                                                                           q2add_destruct_d[0],
                                                                           q1adc_destruct_d[0]} & {q4adf_destruct_r,
                                                                                                   q3ade_destruct_r,
                                                                                                   q2add_destruct_r,
                                                                                                   q1adc_destruct_r}));
  assign lizzieLet2_1QNode_Bool_r = (& lizzieLet2_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet2_1QNode_Bool_emitted <= (lizzieLet2_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet2_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet2_1QVal_Bool,QTree_Bool) > [(vadb_destruct,MyBool)] */
  assign vadb_destruct_d = {lizzieLet2_1QVal_Bool_d[3:3],
                            lizzieLet2_1QVal_Bool_d[0]};
  assign lizzieLet2_1QVal_Bool_r = vadb_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet2_2,QTree_Bool) (lizzieLet2_1,QTree_Bool) > [(_15,QTree_Bool),
                                                                               (lizzieLet2_1QVal_Bool,QTree_Bool),
                                                                               (lizzieLet2_1QNode_Bool,QTree_Bool),
                                                                               (_14,QTree_Bool)] */
  logic [3:0] lizzieLet2_1_onehotd;
  always_comb
    if ((lizzieLet2_2_d[0] && lizzieLet2_1_d[0]))
      unique case (lizzieLet2_2_d[2:1])
        2'd0: lizzieLet2_1_onehotd = 4'd1;
        2'd1: lizzieLet2_1_onehotd = 4'd2;
        2'd2: lizzieLet2_1_onehotd = 4'd4;
        2'd3: lizzieLet2_1_onehotd = 4'd8;
        default: lizzieLet2_1_onehotd = 4'd0;
      endcase
    else lizzieLet2_1_onehotd = 4'd0;
  assign _15_d = {lizzieLet2_1_d[66:1], lizzieLet2_1_onehotd[0]};
  assign lizzieLet2_1QVal_Bool_d = {lizzieLet2_1_d[66:1],
                                    lizzieLet2_1_onehotd[1]};
  assign lizzieLet2_1QNode_Bool_d = {lizzieLet2_1_d[66:1],
                                     lizzieLet2_1_onehotd[2]};
  assign _14_d = {lizzieLet2_1_d[66:1], lizzieLet2_1_onehotd[3]};
  assign lizzieLet2_1_r = (| (lizzieLet2_1_onehotd & {_14_r,
                                                      lizzieLet2_1QNode_Bool_r,
                                                      lizzieLet2_1QVal_Bool_r,
                                                      _15_r}));
  assign lizzieLet2_2_r = lizzieLet2_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool_Bool) : (lizzieLet2_3,QTree_Bool) (gad8_goMux_mux,MyDTBool_Bool_Bool) > [(_13,MyDTBool_Bool_Bool),
                                                                                                 (lizzieLet2_3QVal_Bool,MyDTBool_Bool_Bool),
                                                                                                 (lizzieLet2_3QNode_Bool,MyDTBool_Bool_Bool),
                                                                                                 (_12,MyDTBool_Bool_Bool)] */
  logic [3:0] gad8_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_3_d[0] && gad8_goMux_mux_d[0]))
      unique case (lizzieLet2_3_d[2:1])
        2'd0: gad8_goMux_mux_onehotd = 4'd1;
        2'd1: gad8_goMux_mux_onehotd = 4'd2;
        2'd2: gad8_goMux_mux_onehotd = 4'd4;
        2'd3: gad8_goMux_mux_onehotd = 4'd8;
        default: gad8_goMux_mux_onehotd = 4'd0;
      endcase
    else gad8_goMux_mux_onehotd = 4'd0;
  assign _13_d = gad8_goMux_mux_onehotd[0];
  assign lizzieLet2_3QVal_Bool_d = gad8_goMux_mux_onehotd[1];
  assign lizzieLet2_3QNode_Bool_d = gad8_goMux_mux_onehotd[2];
  assign _12_d = gad8_goMux_mux_onehotd[3];
  assign gad8_goMux_mux_r = (| (gad8_goMux_mux_onehotd & {_12_r,
                                                          lizzieLet2_3QNode_Bool_r,
                                                          lizzieLet2_3QVal_Bool_r,
                                                          _13_r}));
  assign lizzieLet2_3_r = gad8_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool_Bool) : (lizzieLet2_3QNode_Bool,MyDTBool_Bool_Bool) > [(lizzieLet2_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                                                              (lizzieLet2_3QNode_Bool_2,MyDTBool_Bool_Bool)] */
  logic [1:0] lizzieLet2_3QNode_Bool_emitted;
  logic [1:0] lizzieLet2_3QNode_Bool_done;
  assign lizzieLet2_3QNode_Bool_1_d = (lizzieLet2_3QNode_Bool_d[0] && (! lizzieLet2_3QNode_Bool_emitted[0]));
  assign lizzieLet2_3QNode_Bool_2_d = (lizzieLet2_3QNode_Bool_d[0] && (! lizzieLet2_3QNode_Bool_emitted[1]));
  assign lizzieLet2_3QNode_Bool_done = (lizzieLet2_3QNode_Bool_emitted | ({lizzieLet2_3QNode_Bool_2_d[0],
                                                                           lizzieLet2_3QNode_Bool_1_d[0]} & {lizzieLet2_3QNode_Bool_2_r,
                                                                                                             lizzieLet2_3QNode_Bool_1_r}));
  assign lizzieLet2_3QNode_Bool_r = (& lizzieLet2_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet2_3QNode_Bool_emitted <= (lizzieLet2_3QNode_Bool_r ? 2'd0 :
                                         lizzieLet2_3QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet2_3QNode_Bool_2,MyDTBool_Bool_Bool) > (lizzieLet2_3QNode_Bool_2_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_2_bufchan_d;
  logic lizzieLet2_3QNode_Bool_2_bufchan_r;
  assign lizzieLet2_3QNode_Bool_2_r = ((! lizzieLet2_3QNode_Bool_2_bufchan_d[0]) || lizzieLet2_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_3QNode_Bool_2_r)
        lizzieLet2_3QNode_Bool_2_bufchan_d <= lizzieLet2_3QNode_Bool_2_d;
  MyDTBool_Bool_Bool_t lizzieLet2_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet2_3QNode_Bool_2_bufchan_r = (! lizzieLet2_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_3QNode_Bool_2_argbuf_d = (lizzieLet2_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet2_3QNode_Bool_2_bufchan_buf :
                                              lizzieLet2_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_3QNode_Bool_2_argbuf_r && lizzieLet2_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet2_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_3QNode_Bool_2_argbuf_r) && (! lizzieLet2_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet2_3QNode_Bool_2_bufchan_buf <= lizzieLet2_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool_Bool) : (lizzieLet2_3QVal_Bool,MyDTBool_Bool_Bool) > (lizzieLet2_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t lizzieLet2_3QVal_Bool_bufchan_d;
  logic lizzieLet2_3QVal_Bool_bufchan_r;
  assign lizzieLet2_3QVal_Bool_r = ((! lizzieLet2_3QVal_Bool_bufchan_d[0]) || lizzieLet2_3QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_3QVal_Bool_r)
        lizzieLet2_3QVal_Bool_bufchan_d <= lizzieLet2_3QVal_Bool_d;
  MyDTBool_Bool_Bool_t lizzieLet2_3QVal_Bool_bufchan_buf;
  assign lizzieLet2_3QVal_Bool_bufchan_r = (! lizzieLet2_3QVal_Bool_bufchan_buf[0]);
  assign lizzieLet2_3QVal_Bool_1_argbuf_d = (lizzieLet2_3QVal_Bool_bufchan_buf[0] ? lizzieLet2_3QVal_Bool_bufchan_buf :
                                             lizzieLet2_3QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_3QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_3QVal_Bool_1_argbuf_r && lizzieLet2_3QVal_Bool_bufchan_buf[0]))
        lizzieLet2_3QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_3QVal_Bool_1_argbuf_r) && (! lizzieLet2_3QVal_Bool_bufchan_buf[0])))
        lizzieLet2_3QVal_Bool_bufchan_buf <= lizzieLet2_3QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet2_4,QTree_Bool) (go_6_goMux_data,Go) > [(lizzieLet2_4QNone_Bool,Go),
                                                                  (lizzieLet2_4QVal_Bool,Go),
                                                                  (lizzieLet2_4QNode_Bool,Go),
                                                                  (lizzieLet2_4QError_Bool,Go)] */
  logic [3:0] go_6_goMux_data_onehotd;
  always_comb
    if ((lizzieLet2_4_d[0] && go_6_goMux_data_d[0]))
      unique case (lizzieLet2_4_d[2:1])
        2'd0: go_6_goMux_data_onehotd = 4'd1;
        2'd1: go_6_goMux_data_onehotd = 4'd2;
        2'd2: go_6_goMux_data_onehotd = 4'd4;
        2'd3: go_6_goMux_data_onehotd = 4'd8;
        default: go_6_goMux_data_onehotd = 4'd0;
      endcase
    else go_6_goMux_data_onehotd = 4'd0;
  assign lizzieLet2_4QNone_Bool_d = go_6_goMux_data_onehotd[0];
  assign lizzieLet2_4QVal_Bool_d = go_6_goMux_data_onehotd[1];
  assign lizzieLet2_4QNode_Bool_d = go_6_goMux_data_onehotd[2];
  assign lizzieLet2_4QError_Bool_d = go_6_goMux_data_onehotd[3];
  assign go_6_goMux_data_r = (| (go_6_goMux_data_onehotd & {lizzieLet2_4QError_Bool_r,
                                                            lizzieLet2_4QNode_Bool_r,
                                                            lizzieLet2_4QVal_Bool_r,
                                                            lizzieLet2_4QNone_Bool_r}));
  assign lizzieLet2_4_r = go_6_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet2_4QError_Bool,Go) > [(lizzieLet2_4QError_Bool_1,Go),
                                               (lizzieLet2_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet2_4QError_Bool_emitted;
  logic [1:0] lizzieLet2_4QError_Bool_done;
  assign lizzieLet2_4QError_Bool_1_d = (lizzieLet2_4QError_Bool_d[0] && (! lizzieLet2_4QError_Bool_emitted[0]));
  assign lizzieLet2_4QError_Bool_2_d = (lizzieLet2_4QError_Bool_d[0] && (! lizzieLet2_4QError_Bool_emitted[1]));
  assign lizzieLet2_4QError_Bool_done = (lizzieLet2_4QError_Bool_emitted | ({lizzieLet2_4QError_Bool_2_d[0],
                                                                             lizzieLet2_4QError_Bool_1_d[0]} & {lizzieLet2_4QError_Bool_2_r,
                                                                                                                lizzieLet2_4QError_Bool_1_r}));
  assign lizzieLet2_4QError_Bool_r = (& lizzieLet2_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet2_4QError_Bool_emitted <= (lizzieLet2_4QError_Bool_r ? 2'd0 :
                                          lizzieLet2_4QError_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QError_Bool) : [(lizzieLet2_4QError_Bool_1,Go)] > (lizzieLet2_4QError_Bool_1QError_Bool,QTree_Bool) */
  assign lizzieLet2_4QError_Bool_1QError_Bool_d = QError_Bool_dc((& {lizzieLet2_4QError_Bool_1_d[0]}), lizzieLet2_4QError_Bool_1_d);
  assign {lizzieLet2_4QError_Bool_1_r} = {1 {(lizzieLet2_4QError_Bool_1QError_Bool_r && lizzieLet2_4QError_Bool_1QError_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet2_4QError_Bool_1QError_Bool,QTree_Bool) > (lizzieLet5_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d;
  logic lizzieLet2_4QError_Bool_1QError_Bool_bufchan_r;
  assign lizzieLet2_4QError_Bool_1QError_Bool_r = ((! lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d[0]) || lizzieLet2_4QError_Bool_1QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet2_4QError_Bool_1QError_Bool_r)
        lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d <= lizzieLet2_4QError_Bool_1QError_Bool_d;
  QTree_Bool_t lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf;
  assign lizzieLet2_4QError_Bool_1QError_Bool_bufchan_r = (! lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf[0] ? lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf :
                                  lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf[0]))
        lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf[0])))
        lizzieLet2_4QError_Bool_1QError_Bool_bufchan_buf <= lizzieLet2_4QError_Bool_1QError_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QError_Bool_2,Go) > (lizzieLet2_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet2_4QError_Bool_2_bufchan_d;
  logic lizzieLet2_4QError_Bool_2_bufchan_r;
  assign lizzieLet2_4QError_Bool_2_r = ((! lizzieLet2_4QError_Bool_2_bufchan_d[0]) || lizzieLet2_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QError_Bool_2_r)
        lizzieLet2_4QError_Bool_2_bufchan_d <= lizzieLet2_4QError_Bool_2_d;
  Go_t lizzieLet2_4QError_Bool_2_bufchan_buf;
  assign lizzieLet2_4QError_Bool_2_bufchan_r = (! lizzieLet2_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_4QError_Bool_2_argbuf_d = (lizzieLet2_4QError_Bool_2_bufchan_buf[0] ? lizzieLet2_4QError_Bool_2_bufchan_buf :
                                               lizzieLet2_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QError_Bool_2_argbuf_r && lizzieLet2_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet2_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QError_Bool_2_argbuf_r) && (! lizzieLet2_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet2_4QError_Bool_2_bufchan_buf <= lizzieLet2_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNode_Bool,Go) > (lizzieLet2_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet2_4QNode_Bool_bufchan_d;
  logic lizzieLet2_4QNode_Bool_bufchan_r;
  assign lizzieLet2_4QNode_Bool_r = ((! lizzieLet2_4QNode_Bool_bufchan_d[0]) || lizzieLet2_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNode_Bool_r)
        lizzieLet2_4QNode_Bool_bufchan_d <= lizzieLet2_4QNode_Bool_d;
  Go_t lizzieLet2_4QNode_Bool_bufchan_buf;
  assign lizzieLet2_4QNode_Bool_bufchan_r = (! lizzieLet2_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet2_4QNode_Bool_1_argbuf_d = (lizzieLet2_4QNode_Bool_bufchan_buf[0] ? lizzieLet2_4QNode_Bool_bufchan_buf :
                                              lizzieLet2_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNode_Bool_1_argbuf_r && lizzieLet2_4QNode_Bool_bufchan_buf[0]))
        lizzieLet2_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNode_Bool_1_argbuf_r) && (! lizzieLet2_4QNode_Bool_bufchan_buf[0])))
        lizzieLet2_4QNode_Bool_bufchan_buf <= lizzieLet2_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet2_4QNone_Bool,Go) > [(lizzieLet2_4QNone_Bool_1,Go),
                                              (lizzieLet2_4QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet2_4QNone_Bool_emitted;
  logic [1:0] lizzieLet2_4QNone_Bool_done;
  assign lizzieLet2_4QNone_Bool_1_d = (lizzieLet2_4QNone_Bool_d[0] && (! lizzieLet2_4QNone_Bool_emitted[0]));
  assign lizzieLet2_4QNone_Bool_2_d = (lizzieLet2_4QNone_Bool_d[0] && (! lizzieLet2_4QNone_Bool_emitted[1]));
  assign lizzieLet2_4QNone_Bool_done = (lizzieLet2_4QNone_Bool_emitted | ({lizzieLet2_4QNone_Bool_2_d[0],
                                                                           lizzieLet2_4QNone_Bool_1_d[0]} & {lizzieLet2_4QNone_Bool_2_r,
                                                                                                             lizzieLet2_4QNone_Bool_1_r}));
  assign lizzieLet2_4QNone_Bool_r = (& lizzieLet2_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet2_4QNone_Bool_emitted <= (lizzieLet2_4QNone_Bool_r ? 2'd0 :
                                         lizzieLet2_4QNone_Bool_done);
  
  /* dcon (Ty QTree_Bool,
      Dcon QNone_Bool) : [(lizzieLet2_4QNone_Bool_1,Go)] > (lizzieLet2_4QNone_Bool_1QNone_Bool,QTree_Bool) */
  assign lizzieLet2_4QNone_Bool_1QNone_Bool_d = QNone_Bool_dc((& {lizzieLet2_4QNone_Bool_1_d[0]}), lizzieLet2_4QNone_Bool_1_d);
  assign {lizzieLet2_4QNone_Bool_1_r} = {1 {(lizzieLet2_4QNone_Bool_1QNone_Bool_r && lizzieLet2_4QNone_Bool_1QNone_Bool_d[0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet2_4QNone_Bool_1QNone_Bool,QTree_Bool) > (lizzieLet3_1_argbuf,QTree_Bool) */
  QTree_Bool_t lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d;
  logic lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_r;
  assign lizzieLet2_4QNone_Bool_1QNone_Bool_r = ((! lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d[0]) || lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet2_4QNone_Bool_1QNone_Bool_r)
        lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d <= lizzieLet2_4QNone_Bool_1QNone_Bool_d;
  QTree_Bool_t lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf;
  assign lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_r = (! lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf[0]);
  assign lizzieLet3_1_argbuf_d = (lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf[0] ? lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf :
                                  lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet3_1_argbuf_r && lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf[0]))
        lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet3_1_argbuf_r) && (! lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf[0])))
        lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_buf <= lizzieLet2_4QNone_Bool_1QNone_Bool_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet2_4QNone_Bool_2,Go) > (lizzieLet2_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet2_4QNone_Bool_2_bufchan_d;
  logic lizzieLet2_4QNone_Bool_2_bufchan_r;
  assign lizzieLet2_4QNone_Bool_2_r = ((! lizzieLet2_4QNone_Bool_2_bufchan_d[0]) || lizzieLet2_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QNone_Bool_2_r)
        lizzieLet2_4QNone_Bool_2_bufchan_d <= lizzieLet2_4QNone_Bool_2_d;
  Go_t lizzieLet2_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet2_4QNone_Bool_2_bufchan_r = (! lizzieLet2_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_4QNone_Bool_2_argbuf_d = (lizzieLet2_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet2_4QNone_Bool_2_bufchan_buf :
                                              lizzieLet2_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QNone_Bool_2_argbuf_r && lizzieLet2_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet2_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QNone_Bool_2_argbuf_r) && (! lizzieLet2_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet2_4QNone_Bool_2_bufchan_buf <= lizzieLet2_4QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet2_4QNone_Bool_2_argbuf,Go),
                           (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf,Go),
                           (lizzieLet2_4QVal_Bool_2_argbuf,Go),
                           (lizzieLet2_4QError_Bool_2_argbuf,Go)] > (go_13_goMux_choice,C4) (go_13_goMux_data,Go) */
  logic [3:0] lizzieLet2_4QNone_Bool_2_argbuf_select_d;
  assign lizzieLet2_4QNone_Bool_2_argbuf_select_d = ((| lizzieLet2_4QNone_Bool_2_argbuf_select_q) ? lizzieLet2_4QNone_Bool_2_argbuf_select_q :
                                                     (lizzieLet2_4QNone_Bool_2_argbuf_d[0] ? 4'd1 :
                                                      (lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d[0] ? 4'd2 :
                                                       (lizzieLet2_4QVal_Bool_2_argbuf_d[0] ? 4'd4 :
                                                        (lizzieLet2_4QError_Bool_2_argbuf_d[0] ? 4'd8 :
                                                         4'd0)))));
  logic [3:0] lizzieLet2_4QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNone_Bool_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet2_4QNone_Bool_2_argbuf_select_q <= (lizzieLet2_4QNone_Bool_2_argbuf_done ? 4'd0 :
                                                   lizzieLet2_4QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet2_4QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_4QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet2_4QNone_Bool_2_argbuf_emit_q <= (lizzieLet2_4QNone_Bool_2_argbuf_done ? 2'd0 :
                                                 lizzieLet2_4QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet2_4QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet2_4QNone_Bool_2_argbuf_emit_d = (lizzieLet2_4QNone_Bool_2_argbuf_emit_q | ({go_13_goMux_choice_d[0],
                                                                                              go_13_goMux_data_d[0]} & {go_13_goMux_choice_r,
                                                                                                                        go_13_goMux_data_r}));
  logic lizzieLet2_4QNone_Bool_2_argbuf_done;
  assign lizzieLet2_4QNone_Bool_2_argbuf_done = (& lizzieLet2_4QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet2_4QError_Bool_2_argbuf_r,
          lizzieLet2_4QVal_Bool_2_argbuf_r,
          lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_r,
          lizzieLet2_4QNone_Bool_2_argbuf_r} = (lizzieLet2_4QNone_Bool_2_argbuf_done ? lizzieLet2_4QNone_Bool_2_argbuf_select_d :
                                                4'd0);
  assign go_13_goMux_data_d = ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet2_4QNone_Bool_2_argbuf_d :
                               ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet24_3Lcall_kron_kron_Bool_Bool_Bool0_1_argbuf_d :
                                ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet2_4QVal_Bool_2_argbuf_d :
                                 ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet2_4QError_Bool_2_argbuf_d :
                                  1'd0))));
  assign go_13_goMux_choice_d = ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet2_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet2_4QNone_Bool_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet2_4QVal_Bool,Go) > [(lizzieLet2_4QVal_Bool_1,Go),
                                             (lizzieLet2_4QVal_Bool_2,Go)] */
  logic [1:0] lizzieLet2_4QVal_Bool_emitted;
  logic [1:0] lizzieLet2_4QVal_Bool_done;
  assign lizzieLet2_4QVal_Bool_1_d = (lizzieLet2_4QVal_Bool_d[0] && (! lizzieLet2_4QVal_Bool_emitted[0]));
  assign lizzieLet2_4QVal_Bool_2_d = (lizzieLet2_4QVal_Bool_d[0] && (! lizzieLet2_4QVal_Bool_emitted[1]));
  assign lizzieLet2_4QVal_Bool_done = (lizzieLet2_4QVal_Bool_emitted | ({lizzieLet2_4QVal_Bool_2_d[0],
                                                                         lizzieLet2_4QVal_Bool_1_d[0]} & {lizzieLet2_4QVal_Bool_2_r,
                                                                                                          lizzieLet2_4QVal_Bool_1_r}));
  assign lizzieLet2_4QVal_Bool_r = (& lizzieLet2_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Bool_emitted <= 2'd0;
    else
      lizzieLet2_4QVal_Bool_emitted <= (lizzieLet2_4QVal_Bool_r ? 2'd0 :
                                        lizzieLet2_4QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Bool_1,Go) > (lizzieLet2_4QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Bool_1_bufchan_d;
  logic lizzieLet2_4QVal_Bool_1_bufchan_r;
  assign lizzieLet2_4QVal_Bool_1_r = ((! lizzieLet2_4QVal_Bool_1_bufchan_d[0]) || lizzieLet2_4QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Bool_1_r)
        lizzieLet2_4QVal_Bool_1_bufchan_d <= lizzieLet2_4QVal_Bool_1_d;
  Go_t lizzieLet2_4QVal_Bool_1_bufchan_buf;
  assign lizzieLet2_4QVal_Bool_1_bufchan_r = (! lizzieLet2_4QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Bool_1_argbuf_d = (lizzieLet2_4QVal_Bool_1_bufchan_buf[0] ? lizzieLet2_4QVal_Bool_1_bufchan_buf :
                                             lizzieLet2_4QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Bool_1_argbuf_r && lizzieLet2_4QVal_Bool_1_bufchan_buf[0]))
        lizzieLet2_4QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Bool_1_argbuf_r) && (! lizzieLet2_4QVal_Bool_1_bufchan_buf[0])))
        lizzieLet2_4QVal_Bool_1_bufchan_buf <= lizzieLet2_4QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool,
      Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) : [(lizzieLet2_4QVal_Bool_1_argbuf,Go),
                                                                                        (lizzieLet2_5QVal_Bool_1_argbuf,MyDTBool_Bool),
                                                                                        (lizzieLet2_3QVal_Bool_1_argbuf,MyDTBool_Bool_Bool),
                                                                                        (vadb_1_argbuf,MyBool),
                                                                                        (lizzieLet2_6QVal_Bool_1_argbuf,Pointer_QTree_Bool)] > (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) */
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d  = TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_dc((& {lizzieLet2_4QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet2_5QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet2_3QVal_Bool_1_argbuf_d[0],
                                                                                                                                                                                                    vadb_1_argbuf_d[0],
                                                                                                                                                                                                    lizzieLet2_6QVal_Bool_1_argbuf_d[0]}), lizzieLet2_4QVal_Bool_1_argbuf_d, lizzieLet2_5QVal_Bool_1_argbuf_d, lizzieLet2_3QVal_Bool_1_argbuf_d, vadb_1_argbuf_d, lizzieLet2_6QVal_Bool_1_argbuf_d);
  assign {lizzieLet2_4QVal_Bool_1_argbuf_r,
          lizzieLet2_5QVal_Bool_1_argbuf_r,
          lizzieLet2_3QVal_Bool_1_argbuf_r,
          vadb_1_argbuf_r,
          lizzieLet2_6QVal_Bool_1_argbuf_r} = {5 {(\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet2_4QVal_Bool_2,Go) > (lizzieLet2_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet2_4QVal_Bool_2_bufchan_d;
  logic lizzieLet2_4QVal_Bool_2_bufchan_r;
  assign lizzieLet2_4QVal_Bool_2_r = ((! lizzieLet2_4QVal_Bool_2_bufchan_d[0]) || lizzieLet2_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_4QVal_Bool_2_r)
        lizzieLet2_4QVal_Bool_2_bufchan_d <= lizzieLet2_4QVal_Bool_2_d;
  Go_t lizzieLet2_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet2_4QVal_Bool_2_bufchan_r = (! lizzieLet2_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_4QVal_Bool_2_argbuf_d = (lizzieLet2_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet2_4QVal_Bool_2_bufchan_buf :
                                             lizzieLet2_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_4QVal_Bool_2_argbuf_r && lizzieLet2_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet2_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_4QVal_Bool_2_argbuf_r) && (! lizzieLet2_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet2_4QVal_Bool_2_bufchan_buf <= lizzieLet2_4QVal_Bool_2_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Bool) : (lizzieLet2_5,QTree_Bool) (isZad7_goMux_mux,MyDTBool_Bool) > [(_11,MyDTBool_Bool),
                                                                                         (lizzieLet2_5QVal_Bool,MyDTBool_Bool),
                                                                                         (lizzieLet2_5QNode_Bool,MyDTBool_Bool),
                                                                                         (_10,MyDTBool_Bool)] */
  logic [3:0] isZad7_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_5_d[0] && isZad7_goMux_mux_d[0]))
      unique case (lizzieLet2_5_d[2:1])
        2'd0: isZad7_goMux_mux_onehotd = 4'd1;
        2'd1: isZad7_goMux_mux_onehotd = 4'd2;
        2'd2: isZad7_goMux_mux_onehotd = 4'd4;
        2'd3: isZad7_goMux_mux_onehotd = 4'd8;
        default: isZad7_goMux_mux_onehotd = 4'd0;
      endcase
    else isZad7_goMux_mux_onehotd = 4'd0;
  assign _11_d = isZad7_goMux_mux_onehotd[0];
  assign lizzieLet2_5QVal_Bool_d = isZad7_goMux_mux_onehotd[1];
  assign lizzieLet2_5QNode_Bool_d = isZad7_goMux_mux_onehotd[2];
  assign _10_d = isZad7_goMux_mux_onehotd[3];
  assign isZad7_goMux_mux_r = (| (isZad7_goMux_mux_onehotd & {_10_r,
                                                              lizzieLet2_5QNode_Bool_r,
                                                              lizzieLet2_5QVal_Bool_r,
                                                              _11_r}));
  assign lizzieLet2_5_r = isZad7_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Bool) : (lizzieLet2_5QNode_Bool,MyDTBool_Bool) > [(lizzieLet2_5QNode_Bool_1,MyDTBool_Bool),
                                                                    (lizzieLet2_5QNode_Bool_2,MyDTBool_Bool)] */
  logic [1:0] lizzieLet2_5QNode_Bool_emitted;
  logic [1:0] lizzieLet2_5QNode_Bool_done;
  assign lizzieLet2_5QNode_Bool_1_d = (lizzieLet2_5QNode_Bool_d[0] && (! lizzieLet2_5QNode_Bool_emitted[0]));
  assign lizzieLet2_5QNode_Bool_2_d = (lizzieLet2_5QNode_Bool_d[0] && (! lizzieLet2_5QNode_Bool_emitted[1]));
  assign lizzieLet2_5QNode_Bool_done = (lizzieLet2_5QNode_Bool_emitted | ({lizzieLet2_5QNode_Bool_2_d[0],
                                                                           lizzieLet2_5QNode_Bool_1_d[0]} & {lizzieLet2_5QNode_Bool_2_r,
                                                                                                             lizzieLet2_5QNode_Bool_1_r}));
  assign lizzieLet2_5QNode_Bool_r = (& lizzieLet2_5QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_5QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet2_5QNode_Bool_emitted <= (lizzieLet2_5QNode_Bool_r ? 2'd0 :
                                         lizzieLet2_5QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet2_5QNode_Bool_2,MyDTBool_Bool) > (lizzieLet2_5QNode_Bool_2_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_2_bufchan_d;
  logic lizzieLet2_5QNode_Bool_2_bufchan_r;
  assign lizzieLet2_5QNode_Bool_2_r = ((! lizzieLet2_5QNode_Bool_2_bufchan_d[0]) || lizzieLet2_5QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_5QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_5QNode_Bool_2_r)
        lizzieLet2_5QNode_Bool_2_bufchan_d <= lizzieLet2_5QNode_Bool_2_d;
  MyDTBool_Bool_t lizzieLet2_5QNode_Bool_2_bufchan_buf;
  assign lizzieLet2_5QNode_Bool_2_bufchan_r = (! lizzieLet2_5QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_5QNode_Bool_2_argbuf_d = (lizzieLet2_5QNode_Bool_2_bufchan_buf[0] ? lizzieLet2_5QNode_Bool_2_bufchan_buf :
                                              lizzieLet2_5QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_5QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_5QNode_Bool_2_argbuf_r && lizzieLet2_5QNode_Bool_2_bufchan_buf[0]))
        lizzieLet2_5QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_5QNode_Bool_2_argbuf_r) && (! lizzieLet2_5QNode_Bool_2_bufchan_buf[0])))
        lizzieLet2_5QNode_Bool_2_bufchan_buf <= lizzieLet2_5QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Bool) : (lizzieLet2_5QVal_Bool,MyDTBool_Bool) > (lizzieLet2_5QVal_Bool_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t lizzieLet2_5QVal_Bool_bufchan_d;
  logic lizzieLet2_5QVal_Bool_bufchan_r;
  assign lizzieLet2_5QVal_Bool_r = ((! lizzieLet2_5QVal_Bool_bufchan_d[0]) || lizzieLet2_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_5QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet2_5QVal_Bool_r)
        lizzieLet2_5QVal_Bool_bufchan_d <= lizzieLet2_5QVal_Bool_d;
  MyDTBool_Bool_t lizzieLet2_5QVal_Bool_bufchan_buf;
  assign lizzieLet2_5QVal_Bool_bufchan_r = (! lizzieLet2_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet2_5QVal_Bool_1_argbuf_d = (lizzieLet2_5QVal_Bool_bufchan_buf[0] ? lizzieLet2_5QVal_Bool_bufchan_buf :
                                             lizzieLet2_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_5QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet2_5QVal_Bool_1_argbuf_r && lizzieLet2_5QVal_Bool_bufchan_buf[0]))
        lizzieLet2_5QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet2_5QVal_Bool_1_argbuf_r) && (! lizzieLet2_5QVal_Bool_bufchan_buf[0])))
        lizzieLet2_5QVal_Bool_bufchan_buf <= lizzieLet2_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet2_6,QTree_Bool) (m2ada_goMux_mux,Pointer_QTree_Bool) > [(_9,Pointer_QTree_Bool),
                                                                                                  (lizzieLet2_6QVal_Bool,Pointer_QTree_Bool),
                                                                                                  (lizzieLet2_6QNode_Bool,Pointer_QTree_Bool),
                                                                                                  (_8,Pointer_QTree_Bool)] */
  logic [3:0] m2ada_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_6_d[0] && m2ada_goMux_mux_d[0]))
      unique case (lizzieLet2_6_d[2:1])
        2'd0: m2ada_goMux_mux_onehotd = 4'd1;
        2'd1: m2ada_goMux_mux_onehotd = 4'd2;
        2'd2: m2ada_goMux_mux_onehotd = 4'd4;
        2'd3: m2ada_goMux_mux_onehotd = 4'd8;
        default: m2ada_goMux_mux_onehotd = 4'd0;
      endcase
    else m2ada_goMux_mux_onehotd = 4'd0;
  assign _9_d = {m2ada_goMux_mux_d[16:1],
                 m2ada_goMux_mux_onehotd[0]};
  assign lizzieLet2_6QVal_Bool_d = {m2ada_goMux_mux_d[16:1],
                                    m2ada_goMux_mux_onehotd[1]};
  assign lizzieLet2_6QNode_Bool_d = {m2ada_goMux_mux_d[16:1],
                                     m2ada_goMux_mux_onehotd[2]};
  assign _8_d = {m2ada_goMux_mux_d[16:1],
                 m2ada_goMux_mux_onehotd[3]};
  assign m2ada_goMux_mux_r = (| (m2ada_goMux_mux_onehotd & {_8_r,
                                                            lizzieLet2_6QNode_Bool_r,
                                                            lizzieLet2_6QVal_Bool_r,
                                                            _9_r}));
  assign lizzieLet2_6_r = m2ada_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet2_6QNode_Bool,Pointer_QTree_Bool) > [(lizzieLet2_6QNode_Bool_1,Pointer_QTree_Bool),
                                                                              (lizzieLet2_6QNode_Bool_2,Pointer_QTree_Bool)] */
  logic [1:0] lizzieLet2_6QNode_Bool_emitted;
  logic [1:0] lizzieLet2_6QNode_Bool_done;
  assign lizzieLet2_6QNode_Bool_1_d = {lizzieLet2_6QNode_Bool_d[16:1],
                                       (lizzieLet2_6QNode_Bool_d[0] && (! lizzieLet2_6QNode_Bool_emitted[0]))};
  assign lizzieLet2_6QNode_Bool_2_d = {lizzieLet2_6QNode_Bool_d[16:1],
                                       (lizzieLet2_6QNode_Bool_d[0] && (! lizzieLet2_6QNode_Bool_emitted[1]))};
  assign lizzieLet2_6QNode_Bool_done = (lizzieLet2_6QNode_Bool_emitted | ({lizzieLet2_6QNode_Bool_2_d[0],
                                                                           lizzieLet2_6QNode_Bool_1_d[0]} & {lizzieLet2_6QNode_Bool_2_r,
                                                                                                             lizzieLet2_6QNode_Bool_1_r}));
  assign lizzieLet2_6QNode_Bool_r = (& lizzieLet2_6QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet2_6QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet2_6QNode_Bool_emitted <= (lizzieLet2_6QNode_Bool_r ? 2'd0 :
                                         lizzieLet2_6QNode_Bool_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet2_6QNode_Bool_2,Pointer_QTree_Bool) > (lizzieLet2_6QNode_Bool_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_2_bufchan_d;
  logic lizzieLet2_6QNode_Bool_2_bufchan_r;
  assign lizzieLet2_6QNode_Bool_2_r = ((! lizzieLet2_6QNode_Bool_2_bufchan_d[0]) || lizzieLet2_6QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_6QNode_Bool_2_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_6QNode_Bool_2_r)
        lizzieLet2_6QNode_Bool_2_bufchan_d <= lizzieLet2_6QNode_Bool_2_d;
  Pointer_QTree_Bool_t lizzieLet2_6QNode_Bool_2_bufchan_buf;
  assign lizzieLet2_6QNode_Bool_2_bufchan_r = (! lizzieLet2_6QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet2_6QNode_Bool_2_argbuf_d = (lizzieLet2_6QNode_Bool_2_bufchan_buf[0] ? lizzieLet2_6QNode_Bool_2_bufchan_buf :
                                              lizzieLet2_6QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_6QNode_Bool_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_6QNode_Bool_2_argbuf_r && lizzieLet2_6QNode_Bool_2_bufchan_buf[0]))
        lizzieLet2_6QNode_Bool_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_6QNode_Bool_2_argbuf_r) && (! lizzieLet2_6QNode_Bool_2_bufchan_buf[0])))
        lizzieLet2_6QNode_Bool_2_bufchan_buf <= lizzieLet2_6QNode_Bool_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet2_6QVal_Bool,Pointer_QTree_Bool) > (lizzieLet2_6QVal_Bool_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t lizzieLet2_6QVal_Bool_bufchan_d;
  logic lizzieLet2_6QVal_Bool_bufchan_r;
  assign lizzieLet2_6QVal_Bool_r = ((! lizzieLet2_6QVal_Bool_bufchan_d[0]) || lizzieLet2_6QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_6QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_6QVal_Bool_r)
        lizzieLet2_6QVal_Bool_bufchan_d <= lizzieLet2_6QVal_Bool_d;
  Pointer_QTree_Bool_t lizzieLet2_6QVal_Bool_bufchan_buf;
  assign lizzieLet2_6QVal_Bool_bufchan_r = (! lizzieLet2_6QVal_Bool_bufchan_buf[0]);
  assign lizzieLet2_6QVal_Bool_1_argbuf_d = (lizzieLet2_6QVal_Bool_bufchan_buf[0] ? lizzieLet2_6QVal_Bool_bufchan_buf :
                                             lizzieLet2_6QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_6QVal_Bool_1_argbuf_r && lizzieLet2_6QVal_Bool_bufchan_buf[0]))
        lizzieLet2_6QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_6QVal_Bool_1_argbuf_r) && (! lizzieLet2_6QVal_Bool_bufchan_buf[0])))
        lizzieLet2_6QVal_Bool_bufchan_buf <= lizzieLet2_6QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet2_7,QTree_Bool) (sc_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) > [(lizzieLet2_7QNone_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet2_7QVal_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet2_7QNode_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                                                                                                                 (lizzieLet2_7QError_Bool,Pointer_CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet2_7_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet2_7_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet2_7QNone_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet2_7QVal_Bool_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet2_7QNode_Bool_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet2_7QError_Bool_d = {sc_0_goMux_mux_d[16:1],
                                      sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet2_7QError_Bool_r,
                                                          lizzieLet2_7QNode_Bool_r,
                                                          lizzieLet2_7QVal_Bool_r,
                                                          lizzieLet2_7QNone_Bool_r}));
  assign lizzieLet2_7_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet2_7QError_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet2_7QError_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QError_Bool_bufchan_d;
  logic lizzieLet2_7QError_Bool_bufchan_r;
  assign lizzieLet2_7QError_Bool_r = ((! lizzieLet2_7QError_Bool_bufchan_d[0]) || lizzieLet2_7QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_7QError_Bool_r)
        lizzieLet2_7QError_Bool_bufchan_d <= lizzieLet2_7QError_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QError_Bool_bufchan_buf;
  assign lizzieLet2_7QError_Bool_bufchan_r = (! lizzieLet2_7QError_Bool_bufchan_buf[0]);
  assign lizzieLet2_7QError_Bool_1_argbuf_d = (lizzieLet2_7QError_Bool_bufchan_buf[0] ? lizzieLet2_7QError_Bool_bufchan_buf :
                                               lizzieLet2_7QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_7QError_Bool_1_argbuf_r && lizzieLet2_7QError_Bool_bufchan_buf[0]))
        lizzieLet2_7QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_7QError_Bool_1_argbuf_r) && (! lizzieLet2_7QError_Bool_bufchan_buf[0])))
        lizzieLet2_7QError_Bool_bufchan_buf <= lizzieLet2_7QError_Bool_bufchan_d;
  
  /* dcon (Ty CTkron_kron_Bool_Bool_Bool,
      Dcon Lcall_kron_kron_Bool_Bool_Bool3) : [(lizzieLet2_7QNode_Bool,Pointer_CTkron_kron_Bool_Bool_Bool),
                                               (lizzieLet2_5QNode_Bool_1,MyDTBool_Bool),
                                               (lizzieLet2_3QNode_Bool_1,MyDTBool_Bool_Bool),
                                               (q1adc_destruct,Pointer_QTree_Bool),
                                               (lizzieLet2_6QNode_Bool_1,Pointer_QTree_Bool),
                                               (q2add_destruct,Pointer_QTree_Bool),
                                               (q3ade_destruct,Pointer_QTree_Bool)] > (lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) */
  assign lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_d = Lcall_kron_kron_Bool_Bool_Bool3_dc((& {lizzieLet2_7QNode_Bool_d[0],
                                                                                                                                                                                                         lizzieLet2_5QNode_Bool_1_d[0],
                                                                                                                                                                                                         lizzieLet2_3QNode_Bool_1_d[0],
                                                                                                                                                                                                         q1adc_destruct_d[0],
                                                                                                                                                                                                         lizzieLet2_6QNode_Bool_1_d[0],
                                                                                                                                                                                                         q2add_destruct_d[0],
                                                                                                                                                                                                         q3ade_destruct_d[0]}), lizzieLet2_7QNode_Bool_d, lizzieLet2_5QNode_Bool_1_d, lizzieLet2_3QNode_Bool_1_d, q1adc_destruct_d, lizzieLet2_6QNode_Bool_1_d, q2add_destruct_d, q3ade_destruct_d);
  assign {lizzieLet2_7QNode_Bool_r,
          lizzieLet2_5QNode_Bool_1_r,
          lizzieLet2_3QNode_Bool_1_r,
          q1adc_destruct_r,
          lizzieLet2_6QNode_Bool_1_r,
          q2add_destruct_r,
          q3ade_destruct_r} = {7 {(lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_r && lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_d[0])}};
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3,CTkron_kron_Bool_Bool_Bool) > (lizzieLet4_1_argbuf,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  logic lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r;
  assign lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_r = ((! lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d[0]) || lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= {83'd0,
                                                                                                                                                                         1'd0};
    else
      if (lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_r)
        lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d <= lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_d;
  CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf;
  assign lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_r = (! lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]);
  assign lizzieLet4_1_argbuf_d = (lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0] ? lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf :
                                  lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= {83'd0,
                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet4_1_argbuf_r && lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0]))
        lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= {83'd0,
                                                                                                                                                                             1'd0};
      else if (((! lizzieLet4_1_argbuf_r) && (! lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf[0])))
        lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_buf <= lizzieLet2_7QNode_Bool_1lizzieLet2_5QNode_Bool_1lizzieLet2_3QNode_Bool_1q1adc_1lizzieLet2_6QNode_Bool_1q2add_1q3ade_1Lcall_kron_kron_Bool_Bool_Bool3_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet2_7QNone_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet2_7QNone_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNone_Bool_bufchan_d;
  logic lizzieLet2_7QNone_Bool_bufchan_r;
  assign lizzieLet2_7QNone_Bool_r = ((! lizzieLet2_7QNone_Bool_bufchan_d[0]) || lizzieLet2_7QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_7QNone_Bool_r)
        lizzieLet2_7QNone_Bool_bufchan_d <= lizzieLet2_7QNone_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QNone_Bool_bufchan_buf;
  assign lizzieLet2_7QNone_Bool_bufchan_r = (! lizzieLet2_7QNone_Bool_bufchan_buf[0]);
  assign lizzieLet2_7QNone_Bool_1_argbuf_d = (lizzieLet2_7QNone_Bool_bufchan_buf[0] ? lizzieLet2_7QNone_Bool_bufchan_buf :
                                              lizzieLet2_7QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_7QNone_Bool_1_argbuf_r && lizzieLet2_7QNone_Bool_bufchan_buf[0]))
        lizzieLet2_7QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_7QNone_Bool_1_argbuf_r) && (! lizzieLet2_7QNone_Bool_bufchan_buf[0])))
        lizzieLet2_7QNone_Bool_bufchan_buf <= lizzieLet2_7QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (lizzieLet2_7QVal_Bool,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet2_7QVal_Bool_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QVal_Bool_bufchan_d;
  logic lizzieLet2_7QVal_Bool_bufchan_r;
  assign lizzieLet2_7QVal_Bool_r = ((! lizzieLet2_7QVal_Bool_bufchan_d[0]) || lizzieLet2_7QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QVal_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet2_7QVal_Bool_r)
        lizzieLet2_7QVal_Bool_bufchan_d <= lizzieLet2_7QVal_Bool_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t lizzieLet2_7QVal_Bool_bufchan_buf;
  assign lizzieLet2_7QVal_Bool_bufchan_r = (! lizzieLet2_7QVal_Bool_bufchan_buf[0]);
  assign lizzieLet2_7QVal_Bool_1_argbuf_d = (lizzieLet2_7QVal_Bool_bufchan_buf[0] ? lizzieLet2_7QVal_Bool_bufchan_buf :
                                             lizzieLet2_7QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet2_7QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_7QVal_Bool_1_argbuf_r && lizzieLet2_7QVal_Bool_bufchan_buf[0]))
        lizzieLet2_7QVal_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_7QVal_Bool_1_argbuf_r) && (! lizzieLet2_7QVal_Bool_bufchan_buf[0])))
        lizzieLet2_7QVal_Bool_bufchan_buf <= lizzieLet2_7QVal_Bool_bufchan_d;
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool0) : (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) > [(es_2_4_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_3_7_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_4_6_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_14_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted ;
  logic [3:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_done ;
  assign es_2_4_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [19:4],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [0]))};
  assign es_3_7_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [35:20],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [1]))};
  assign es_4_6_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [51:36],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [2]))};
  assign sc_0_14_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [67:52],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted [3]))};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_done  = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  | ({sc_0_14_destruct_d[0],
                                                                                                                               es_4_6_destruct_d[0],
                                                                                                                               es_3_7_destruct_d[0],
                                                                                                                               es_2_4_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                                                        es_4_6_destruct_r,
                                                                                                                                                        es_3_7_destruct_r,
                                                                                                                                                        es_2_4_destruct_r}));
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_r  = (& \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  <= 4'd0;
    else
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_emitted  <= (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_r  ? 4'd0 :
                                                                   \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool1) : (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) > [(es_3_6_destruct,Pointer_QTree_Bool),
                                                                                                                                     (es_4_5_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_13_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacY_4_destruct,MyDTBool_Bool),
                                                                                                                                     (gacZ_4_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'ad0_4_destruct,MyBool),
                                                                                                                                     (q1ad3_3_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted ;
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_done ;
  assign es_3_6_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [19:4],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [0]))};
  assign es_4_5_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [35:20],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [1]))};
  assign sc_0_13_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [51:36],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [2]))};
  assign isZacY_4_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [3]));
  assign gacZ_4_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [4]));
  assign \v'ad0_4_destruct_d  = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [52:52],
                                 (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [5]))};
  assign q1ad3_3_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [68:53],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted [6]))};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_done  = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  | ({q1ad3_3_destruct_d[0],
                                                                                                                               \v'ad0_4_destruct_d [0],
                                                                                                                               gacZ_4_destruct_d[0],
                                                                                                                               isZacY_4_destruct_d[0],
                                                                                                                               sc_0_13_destruct_d[0],
                                                                                                                               es_4_5_destruct_d[0],
                                                                                                                               es_3_6_destruct_d[0]} & {q1ad3_3_destruct_r,
                                                                                                                                                        \v'ad0_4_destruct_r ,
                                                                                                                                                        gacZ_4_destruct_r,
                                                                                                                                                        isZacY_4_destruct_r,
                                                                                                                                                        sc_0_13_destruct_r,
                                                                                                                                                        es_4_5_destruct_r,
                                                                                                                                                        es_3_6_destruct_r}));
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_r  = (& \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  <= 7'd0;
    else
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_emitted  <= (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_r  ? 7'd0 :
                                                                   \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool2) : (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) > [(es_4_4_destruct,Pointer_QTree_Bool),
                                                                                                                                     (sc_0_12_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacY_3_destruct,MyDTBool_Bool),
                                                                                                                                     (gacZ_3_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'ad0_3_destruct,MyBool),
                                                                                                                                     (q1ad3_2_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2ad4_2_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted ;
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_done ;
  assign es_4_4_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [19:4],
                              (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [0]))};
  assign sc_0_12_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [35:20],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [1]))};
  assign isZacY_3_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [2]));
  assign gacZ_3_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [3]));
  assign \v'ad0_3_destruct_d  = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [36:36],
                                 (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [4]))};
  assign q1ad3_2_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [52:37],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [5]))};
  assign q2ad4_2_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [68:53],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted [6]))};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_done  = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  | ({q2ad4_2_destruct_d[0],
                                                                                                                               q1ad3_2_destruct_d[0],
                                                                                                                               \v'ad0_3_destruct_d [0],
                                                                                                                               gacZ_3_destruct_d[0],
                                                                                                                               isZacY_3_destruct_d[0],
                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                               es_4_4_destruct_d[0]} & {q2ad4_2_destruct_r,
                                                                                                                                                        q1ad3_2_destruct_r,
                                                                                                                                                        \v'ad0_3_destruct_r ,
                                                                                                                                                        gacZ_3_destruct_r,
                                                                                                                                                        isZacY_3_destruct_r,
                                                                                                                                                        sc_0_12_destruct_r,
                                                                                                                                                        es_4_4_destruct_r}));
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_r  = (& \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  <= 7'd0;
    else
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_emitted  <= (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_r  ? 7'd0 :
                                                                   \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_done );
  
  /* destruct (Ty CTmap''_map''_Bool_Bool_Bool,
          Dcon Lcall_map''_map''_Bool_Bool_Bool3) : (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool) > [(sc_0_11_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                     (isZacY_2_destruct,MyDTBool_Bool),
                                                                                                                                     (gacZ_2_destruct,MyDTBool_Bool_Bool),
                                                                                                                                     (v'ad0_2_destruct,MyBool),
                                                                                                                                     (q1ad3_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q2ad4_1_destruct,Pointer_QTree_Bool),
                                                                                                                                     (q3ad5_1_destruct,Pointer_QTree_Bool)] */
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted ;
  logic [6:0] \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_done ;
  assign sc_0_11_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [19:4],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [0]))};
  assign isZacY_2_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [1]));
  assign gacZ_2_destruct_d = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [2]));
  assign \v'ad0_2_destruct_d  = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [20:20],
                                 (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [3]))};
  assign q1ad3_1_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [36:21],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [4]))};
  assign q2ad4_1_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [52:37],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [5]))};
  assign q3ad5_1_destruct_d = {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [68:53],
                               (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d [0] && (! \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted [6]))};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_done  = (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  | ({q3ad5_1_destruct_d[0],
                                                                                                                               q2ad4_1_destruct_d[0],
                                                                                                                               q1ad3_1_destruct_d[0],
                                                                                                                               \v'ad0_2_destruct_d [0],
                                                                                                                               gacZ_2_destruct_d[0],
                                                                                                                               isZacY_2_destruct_d[0],
                                                                                                                               sc_0_11_destruct_d[0]} & {q3ad5_1_destruct_r,
                                                                                                                                                         q2ad4_1_destruct_r,
                                                                                                                                                         q1ad3_1_destruct_r,
                                                                                                                                                         \v'ad0_2_destruct_r ,
                                                                                                                                                         gacZ_2_destruct_r,
                                                                                                                                                         isZacY_2_destruct_r,
                                                                                                                                                         sc_0_11_destruct_r}));
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_r  = (& \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  <= 7'd0;
    else
      \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_emitted  <= (\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_r  ? 7'd0 :
                                                                   \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_done );
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet34_2,CTmap''_map''_Bool_Bool_Bool) (lizzieLet34_1,CTmap''_map''_Bool_Bool_Bool) > [(_7,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                       (lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool)] */
  logic [4:0] lizzieLet34_1_onehotd;
  always_comb
    if ((lizzieLet34_2_d[0] && lizzieLet34_1_d[0]))
      unique case (lizzieLet34_2_d[3:1])
        3'd0: lizzieLet34_1_onehotd = 5'd1;
        3'd1: lizzieLet34_1_onehotd = 5'd2;
        3'd2: lizzieLet34_1_onehotd = 5'd4;
        3'd3: lizzieLet34_1_onehotd = 5'd8;
        3'd4: lizzieLet34_1_onehotd = 5'd16;
        default: lizzieLet34_1_onehotd = 5'd0;
      endcase
    else lizzieLet34_1_onehotd = 5'd0;
  assign _7_d = {lizzieLet34_1_d[68:1], lizzieLet34_1_onehotd[0]};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_d  = {lizzieLet34_1_d[68:1],
                                                               lizzieLet34_1_onehotd[1]};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_d  = {lizzieLet34_1_d[68:1],
                                                               lizzieLet34_1_onehotd[2]};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_d  = {lizzieLet34_1_d[68:1],
                                                               lizzieLet34_1_onehotd[3]};
  assign \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_d  = {lizzieLet34_1_d[68:1],
                                                               lizzieLet34_1_onehotd[4]};
  assign lizzieLet34_1_r = (| (lizzieLet34_1_onehotd & {\lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                        \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                        \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                        \lizzieLet34_1Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                        _7_r}));
  assign lizzieLet34_2_r = lizzieLet34_1_r;
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty Go) : (lizzieLet34_3,CTmap''_map''_Bool_Bool_Bool) (go_15_goMux_data,Go) > [(_6,Go),
                                                                                      (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3,Go),
                                                                                      (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2,Go),
                                                                                      (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1,Go),
                                                                                      (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet34_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet34_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _6_d = go_15_goMux_data_onehotd[0];
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_d  = go_15_goMux_data_onehotd[1];
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_d  = go_15_goMux_data_onehotd[2];
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_d  = go_15_goMux_data_onehotd[3];
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_d  = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                              \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                              \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                              \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                              _6_r}));
  assign lizzieLet34_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0,Go) > (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_r  = ((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d [0]) || \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_r )
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_d ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r  = (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_d  = (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0] ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  :
                                                                        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r  && \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_1_argbuf_r ) && (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0])))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1,Go) > (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_r  = ((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d [0]) || \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_r )
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_d ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r  = (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_d  = (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0] ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  :
                                                                        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r  && \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_1_argbuf_r ) && (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0])))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2,Go) > (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_r  = ((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d [0]) || \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_r )
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_d ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r  = (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_d  = (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0] ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  :
                                                                        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r  && \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_1_argbuf_r ) && (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0])))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3,Go) > (lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf,Go) */
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  logic \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_r  = ((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d [0]) || \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_r )
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_d ;
  Go_t \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf ;
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_r  = (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]);
  assign \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_d  = (\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0] ? \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  :
                                                                        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r  && \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0]))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_1_argbuf_r ) && (! \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf [0])))
        \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_buf  <= \lizzieLet34_3Lcall_map''_map''_Bool_Bool_Bool3_bufchan_d ;
  
  /* demux (Ty CTmap''_map''_Bool_Bool_Bool,
       Ty Pointer_QTree_Bool) : (lizzieLet34_4,CTmap''_map''_Bool_Bool_Bool) (srtarg_0_2_goMux_mux,Pointer_QTree_Bool) > [(lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                                                                                          (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0,Pointer_QTree_Bool)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet34_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet34_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                             srtarg_0_2_goMux_mux_onehotd[0]};
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[1]};
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[2]};
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[3]};
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_d  = {srtarg_0_2_goMux_mux_d[16:1],
                                                               srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_r ,
                                                                      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_r ,
                                                                      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_r ,
                                                                      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_r ,
                                                                      \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_r }));
  assign lizzieLet34_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Bool,
      Dcon QNode_Bool) : [(lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0,Pointer_QTree_Bool),
                          (es_2_4_destruct,Pointer_QTree_Bool),
                          (es_3_7_destruct,Pointer_QTree_Bool),
                          (es_4_6_destruct,Pointer_QTree_Bool)] > (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool,QTree_Bool) */
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_d  = QNode_Bool_dc((& {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_d [0],
                                                                                                                    es_2_4_destruct_d[0],
                                                                                                                    es_3_7_destruct_d[0],
                                                                                                                    es_4_6_destruct_d[0]}), \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_d , es_2_4_destruct_d, es_3_7_destruct_d, es_4_6_destruct_d);
  assign {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_r ,
          es_2_4_destruct_r,
          es_3_7_destruct_r,
          es_4_6_destruct_r} = {4 {(\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_r  && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_d [0])}};
  
  /* buf (Ty QTree_Bool) : (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool,QTree_Bool) > (lizzieLet38_1_argbuf,QTree_Bool) */
  QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_r ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_r  = ((! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d [0]) || \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d  <= {66'd0,
                                                                                                         1'd0};
    else
      if (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_r )
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_d ;
  QTree_Bool_t \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_r  = (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf [0]);
  assign lizzieLet38_1_argbuf_d = (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf [0] ? \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf  :
                                   \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                           1'd0};
    else
      if ((lizzieLet38_1_argbuf_r && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf [0]))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf  <= {66'd0,
                                                                                                             1'd0};
      else if (((! lizzieLet38_1_argbuf_r) && (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf [0])))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_buf  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool0_1es_2_4_1es_3_7_1es_4_6_1QNode_Bool_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool0) : [(lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1,Pointer_QTree_Bool),
                                                 (es_3_6_destruct,Pointer_QTree_Bool),
                                                 (es_4_5_destruct,Pointer_QTree_Bool),
                                                 (sc_0_13_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool)] > (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d  = \Lcall_map''_map''_Bool_Bool_Bool0_dc ((& {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_d [0],
                                                                                                                                                                     es_3_6_destruct_d[0],
                                                                                                                                                                     es_4_5_destruct_d[0],
                                                                                                                                                                     sc_0_13_destruct_d[0]}), \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_d , es_3_6_destruct_d, es_4_5_destruct_d, sc_0_13_destruct_d);
  assign {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_r ,
          es_3_6_destruct_r,
          es_4_5_destruct_r,
          sc_0_13_destruct_r} = {4 {(\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r  && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet37_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r  = ((! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d [0]) || \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= {68'd0,
                                                                                                                                 1'd0};
    else
      if (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_r )
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_r  = (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]);
  assign lizzieLet37_1_argbuf_d = (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0] ? \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  :
                                   \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= {68'd0,
                                                                                                                                   1'd0};
    else
      if ((lizzieLet37_1_argbuf_r && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0]))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= {68'd0,
                                                                                                                                     1'd0};
      else if (((! lizzieLet37_1_argbuf_r) && (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf [0])))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_buf  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool1_1es_3_6_1es_4_5_1sc_0_13_1Lcall_map''_map''_Bool_Bool_Bool0_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool1) : [(lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2,Pointer_QTree_Bool),
                                                 (es_4_4_destruct,Pointer_QTree_Bool),
                                                 (sc_0_12_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (isZacY_3_1,MyDTBool_Bool),
                                                 (gacZ_3_1,MyDTBool_Bool_Bool),
                                                 (v'ad0_3_1,MyBool),
                                                 (q1ad3_2_destruct,Pointer_QTree_Bool)] > (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_d  = \Lcall_map''_map''_Bool_Bool_Bool1_dc ((& {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_d [0],
                                                                                                                                                                                                 es_4_4_destruct_d[0],
                                                                                                                                                                                                 sc_0_12_destruct_d[0],
                                                                                                                                                                                                 isZacY_3_1_d[0],
                                                                                                                                                                                                 gacZ_3_1_d[0],
                                                                                                                                                                                                 \v'ad0_3_1_d [0],
                                                                                                                                                                                                 q1ad3_2_destruct_d[0]}), \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_d , es_4_4_destruct_d, sc_0_12_destruct_d, isZacY_3_1_d, gacZ_3_1_d, \v'ad0_3_1_d , q1ad3_2_destruct_d);
  assign {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_r ,
          es_4_4_destruct_r,
          sc_0_12_destruct_r,
          isZacY_3_1_r,
          gacZ_3_1_r,
          \v'ad0_3_1_r ,
          q1ad3_2_destruct_r} = {7 {(\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_r  && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet36_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_r  = ((! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d [0]) || \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= {68'd0,
                                                                                                                                                             1'd0};
    else
      if (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_r )
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_r  = (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]);
  assign lizzieLet36_1_argbuf_d = (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0] ? \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  :
                                   \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= {68'd0,
                                                                                                                                                               1'd0};
    else
      if ((lizzieLet36_1_argbuf_r && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0]))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= {68'd0,
                                                                                                                                                                 1'd0};
      else if (((! lizzieLet36_1_argbuf_r) && (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf [0])))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_buf  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool2_1es_4_4_1sc_0_12_1isZacY_3_1gacZ_3_1v'ad0_3_1q1ad3_2_1Lcall_map''_map''_Bool_Bool_Bool1_bufchan_d ;
  
  /* dcon (Ty CTmap''_map''_Bool_Bool_Bool,
      Dcon Lcall_map''_map''_Bool_Bool_Bool2) : [(lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3,Pointer_QTree_Bool),
                                                 (sc_0_11_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool),
                                                 (isZacY_2_1,MyDTBool_Bool),
                                                 (gacZ_2_1,MyDTBool_Bool_Bool),
                                                 (v'ad0_2_1,MyBool),
                                                 (q1ad3_1_destruct,Pointer_QTree_Bool),
                                                 (q2ad4_1_destruct,Pointer_QTree_Bool)] > (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) */
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_d  = \Lcall_map''_map''_Bool_Bool_Bool2_dc ((& {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_d [0],
                                                                                                                                                                                                  sc_0_11_destruct_d[0],
                                                                                                                                                                                                  isZacY_2_1_d[0],
                                                                                                                                                                                                  gacZ_2_1_d[0],
                                                                                                                                                                                                  \v'ad0_2_1_d [0],
                                                                                                                                                                                                  q1ad3_1_destruct_d[0],
                                                                                                                                                                                                  q2ad4_1_destruct_d[0]}), \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_d , sc_0_11_destruct_d, isZacY_2_1_d, gacZ_2_1_d, \v'ad0_2_1_d , q1ad3_1_destruct_d, q2ad4_1_destruct_d);
  assign {\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_r ,
          sc_0_11_destruct_r,
          isZacY_2_1_r,
          gacZ_2_1_r,
          \v'ad0_2_1_r ,
          q1ad3_1_destruct_r,
          q2ad4_1_destruct_r} = {7 {(\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_r  && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_d [0])}};
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2,CTmap''_map''_Bool_Bool_Bool) > (lizzieLet35_1_argbuf,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  logic \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_r  = ((! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d [0]) || \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= {68'd0,
                                                                                                                                                              1'd0};
    else
      if (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_r )
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf ;
  assign \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_r  = (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]);
  assign lizzieLet35_1_argbuf_d = (\lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0] ? \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  :
                                   \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= {68'd0,
                                                                                                                                                                1'd0};
    else
      if ((lizzieLet35_1_argbuf_r && \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0]))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= {68'd0,
                                                                                                                                                                  1'd0};
      else if (((! lizzieLet35_1_argbuf_r) && (! \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf [0])))
        \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_buf  <= \lizzieLet34_4Lcall_map''_map''_Bool_Bool_Bool3_1sc_0_11_1isZacY_2_1gacZ_2_1v'ad0_2_1q1ad3_1_1q2ad4_1_1Lcall_map''_map''_Bool_Bool_Bool2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Bool) : (lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos,Pointer_QTree_Bool) > [(lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool),
                                                                                                    (lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool)] */
  logic [1:0] \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted ;
  logic [1:0] \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_done ;
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d  = {\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d [16:1],
                                                                                  (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d [0] && (! \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted [0]))};
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d  = {\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d [16:1],
                                                                                  (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_d [0] && (! \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted [1]))};
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_done  = (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  | ({\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d [0],
                                                                                                                           \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                                        \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_r  = (& \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  <= 2'd0;
    else
      \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_emitted  <= (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_r  ? 2'd0 :
                                                                 \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_done );
  
  /* togo (Ty Pointer_QTree_Bool) : (lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1,Pointer_QTree_Bool) > (call_map''_map''_Bool_Bool_Bool_goConst,Go) */
  assign \call_map''_map''_Bool_Bool_Bool_goConst_d  = \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_1_r  = \call_map''_map''_Bool_Bool_Bool_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Bool) : (lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2,Pointer_QTree_Bool) > (map''_map''_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                        1'd0};
    else
      if (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_r )
        \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Bool_t \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \map''_map''_Bool_Bool_Bool_resbuf_d  = (\lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  :
                                                  \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                          1'd0};
    else
      if ((\map''_map''_Bool_Bool_Bool_resbuf_r  && \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                            1'd0};
      else if (((! \map''_map''_Bool_Bool_Bool_resbuf_r ) && (! \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet34_4Lmap''_map''_Bool_Bool_Boolsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty QTree_Bool,
          Dcon QNode_Bool) : (lizzieLet6_1QNode_Bool,QTree_Bool) > [(q1acU_destruct,Pointer_QTree_Bool),
                                                                    (q2acV_destruct,Pointer_QTree_Bool),
                                                                    (q3acW_destruct,Pointer_QTree_Bool),
                                                                    (q4acX_destruct,Pointer_QTree_Bool)] */
  logic [3:0] lizzieLet6_1QNode_Bool_emitted;
  logic [3:0] lizzieLet6_1QNode_Bool_done;
  assign q1acU_destruct_d = {lizzieLet6_1QNode_Bool_d[18:3],
                             (lizzieLet6_1QNode_Bool_d[0] && (! lizzieLet6_1QNode_Bool_emitted[0]))};
  assign q2acV_destruct_d = {lizzieLet6_1QNode_Bool_d[34:19],
                             (lizzieLet6_1QNode_Bool_d[0] && (! lizzieLet6_1QNode_Bool_emitted[1]))};
  assign q3acW_destruct_d = {lizzieLet6_1QNode_Bool_d[50:35],
                             (lizzieLet6_1QNode_Bool_d[0] && (! lizzieLet6_1QNode_Bool_emitted[2]))};
  assign q4acX_destruct_d = {lizzieLet6_1QNode_Bool_d[66:51],
                             (lizzieLet6_1QNode_Bool_d[0] && (! lizzieLet6_1QNode_Bool_emitted[3]))};
  assign lizzieLet6_1QNode_Bool_done = (lizzieLet6_1QNode_Bool_emitted | ({q4acX_destruct_d[0],
                                                                           q3acW_destruct_d[0],
                                                                           q2acV_destruct_d[0],
                                                                           q1acU_destruct_d[0]} & {q4acX_destruct_r,
                                                                                                   q3acW_destruct_r,
                                                                                                   q2acV_destruct_r,
                                                                                                   q1acU_destruct_r}));
  assign lizzieLet6_1QNode_Bool_r = (& lizzieLet6_1QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Bool_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Bool_emitted <= (lizzieLet6_1QNode_Bool_r ? 4'd0 :
                                         lizzieLet6_1QNode_Bool_done);
  
  /* destruct (Ty QTree_Bool,
          Dcon QVal_Bool) : (lizzieLet6_1QVal_Bool,QTree_Bool) > [(vacT_destruct,MyBool)] */
  assign vacT_destruct_d = {lizzieLet6_1QVal_Bool_d[3:3],
                            lizzieLet6_1QVal_Bool_d[0]};
  assign lizzieLet6_1QVal_Bool_r = vacT_destruct_r;
  
  /* demux (Ty QTree_Bool,
       Ty QTree_Bool) : (lizzieLet6_2,QTree_Bool) (lizzieLet6_1,QTree_Bool) > [(_5,QTree_Bool),
                                                                               (lizzieLet6_1QVal_Bool,QTree_Bool),
                                                                               (lizzieLet6_1QNode_Bool,QTree_Bool),
                                                                               (_4,QTree_Bool)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _5_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Bool_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Bool_d = {lizzieLet6_1_d[66:1],
                                     lizzieLet6_1_onehotd[2]};
  assign _4_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_4_r,
                                                      lizzieLet6_1QNode_Bool_r,
                                                      lizzieLet6_1QVal_Bool_r,
                                                      _5_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Bool,
       Ty MyDTBool_Nat) : (lizzieLet6_3,QTree_Bool) (gacR_goMux_mux,MyDTBool_Nat) > [(_3,MyDTBool_Nat),
                                                                                     (lizzieLet6_3QVal_Bool,MyDTBool_Nat),
                                                                                     (lizzieLet6_3QNode_Bool,MyDTBool_Nat),
                                                                                     (_2,MyDTBool_Nat)] */
  logic [3:0] gacR_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && gacR_goMux_mux_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: gacR_goMux_mux_onehotd = 4'd1;
        2'd1: gacR_goMux_mux_onehotd = 4'd2;
        2'd2: gacR_goMux_mux_onehotd = 4'd4;
        2'd3: gacR_goMux_mux_onehotd = 4'd8;
        default: gacR_goMux_mux_onehotd = 4'd0;
      endcase
    else gacR_goMux_mux_onehotd = 4'd0;
  assign _3_d = gacR_goMux_mux_onehotd[0];
  assign lizzieLet6_3QVal_Bool_d = gacR_goMux_mux_onehotd[1];
  assign lizzieLet6_3QNode_Bool_d = gacR_goMux_mux_onehotd[2];
  assign _2_d = gacR_goMux_mux_onehotd[3];
  assign gacR_goMux_mux_r = (| (gacR_goMux_mux_onehotd & {_2_r,
                                                          lizzieLet6_3QNode_Bool_r,
                                                          lizzieLet6_3QVal_Bool_r,
                                                          _3_r}));
  assign lizzieLet6_3_r = gacR_goMux_mux_r;
  
  /* fork (Ty MyDTBool_Nat) : (lizzieLet6_3QNode_Bool,MyDTBool_Nat) > [(lizzieLet6_3QNode_Bool_1,MyDTBool_Nat),
                                                                  (lizzieLet6_3QNode_Bool_2,MyDTBool_Nat)] */
  logic [1:0] lizzieLet6_3QNode_Bool_emitted;
  logic [1:0] lizzieLet6_3QNode_Bool_done;
  assign lizzieLet6_3QNode_Bool_1_d = (lizzieLet6_3QNode_Bool_d[0] && (! lizzieLet6_3QNode_Bool_emitted[0]));
  assign lizzieLet6_3QNode_Bool_2_d = (lizzieLet6_3QNode_Bool_d[0] && (! lizzieLet6_3QNode_Bool_emitted[1]));
  assign lizzieLet6_3QNode_Bool_done = (lizzieLet6_3QNode_Bool_emitted | ({lizzieLet6_3QNode_Bool_2_d[0],
                                                                           lizzieLet6_3QNode_Bool_1_d[0]} & {lizzieLet6_3QNode_Bool_2_r,
                                                                                                             lizzieLet6_3QNode_Bool_1_r}));
  assign lizzieLet6_3QNode_Bool_r = (& lizzieLet6_3QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet6_3QNode_Bool_emitted <= (lizzieLet6_3QNode_Bool_r ? 2'd0 :
                                         lizzieLet6_3QNode_Bool_done);
  
  /* buf (Ty MyDTBool_Nat) : (lizzieLet6_3QNode_Bool_2,MyDTBool_Nat) > (lizzieLet6_3QNode_Bool_2_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_2_bufchan_d;
  logic lizzieLet6_3QNode_Bool_2_bufchan_r;
  assign lizzieLet6_3QNode_Bool_2_r = ((! lizzieLet6_3QNode_Bool_2_bufchan_d[0]) || lizzieLet6_3QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNode_Bool_2_r)
        lizzieLet6_3QNode_Bool_2_bufchan_d <= lizzieLet6_3QNode_Bool_2_d;
  MyDTBool_Nat_t lizzieLet6_3QNode_Bool_2_bufchan_buf;
  assign lizzieLet6_3QNode_Bool_2_bufchan_r = (! lizzieLet6_3QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet6_3QNode_Bool_2_argbuf_d = (lizzieLet6_3QNode_Bool_2_bufchan_buf[0] ? lizzieLet6_3QNode_Bool_2_bufchan_buf :
                                              lizzieLet6_3QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNode_Bool_2_argbuf_r && lizzieLet6_3QNode_Bool_2_bufchan_buf[0]))
        lizzieLet6_3QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNode_Bool_2_argbuf_r) && (! lizzieLet6_3QNode_Bool_2_bufchan_buf[0])))
        lizzieLet6_3QNode_Bool_2_bufchan_buf <= lizzieLet6_3QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTBool_Nat) : (lizzieLet6_3QVal_Bool,MyDTBool_Nat) > (lizzieLet6_3QVal_Bool_1_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t lizzieLet6_3QVal_Bool_bufchan_d;
  logic lizzieLet6_3QVal_Bool_bufchan_r;
  assign lizzieLet6_3QVal_Bool_r = ((! lizzieLet6_3QVal_Bool_bufchan_d[0]) || lizzieLet6_3QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QVal_Bool_r)
        lizzieLet6_3QVal_Bool_bufchan_d <= lizzieLet6_3QVal_Bool_d;
  MyDTBool_Nat_t lizzieLet6_3QVal_Bool_bufchan_buf;
  assign lizzieLet6_3QVal_Bool_bufchan_r = (! lizzieLet6_3QVal_Bool_bufchan_buf[0]);
  assign lizzieLet6_3QVal_Bool_1_argbuf_d = (lizzieLet6_3QVal_Bool_bufchan_buf[0] ? lizzieLet6_3QVal_Bool_bufchan_buf :
                                             lizzieLet6_3QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QVal_Bool_1_argbuf_r && lizzieLet6_3QVal_Bool_bufchan_buf[0]))
        lizzieLet6_3QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QVal_Bool_1_argbuf_r) && (! lizzieLet6_3QVal_Bool_bufchan_buf[0])))
        lizzieLet6_3QVal_Bool_bufchan_buf <= lizzieLet6_3QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Go) : (lizzieLet6_4,QTree_Bool) (go_7_goMux_data,Go) > [(lizzieLet6_4QNone_Bool,Go),
                                                                  (lizzieLet6_4QVal_Bool,Go),
                                                                  (lizzieLet6_4QNode_Bool,Go),
                                                                  (lizzieLet6_4QError_Bool,Go)] */
  logic [3:0] go_7_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && go_7_goMux_data_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: go_7_goMux_data_onehotd = 4'd1;
        2'd1: go_7_goMux_data_onehotd = 4'd2;
        2'd2: go_7_goMux_data_onehotd = 4'd4;
        2'd3: go_7_goMux_data_onehotd = 4'd8;
        default: go_7_goMux_data_onehotd = 4'd0;
      endcase
    else go_7_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_4QNone_Bool_d = go_7_goMux_data_onehotd[0];
  assign lizzieLet6_4QVal_Bool_d = go_7_goMux_data_onehotd[1];
  assign lizzieLet6_4QNode_Bool_d = go_7_goMux_data_onehotd[2];
  assign lizzieLet6_4QError_Bool_d = go_7_goMux_data_onehotd[3];
  assign go_7_goMux_data_r = (| (go_7_goMux_data_onehotd & {lizzieLet6_4QError_Bool_r,
                                                            lizzieLet6_4QNode_Bool_r,
                                                            lizzieLet6_4QVal_Bool_r,
                                                            lizzieLet6_4QNone_Bool_r}));
  assign lizzieLet6_4_r = go_7_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_4QError_Bool,Go) > [(lizzieLet6_4QError_Bool_1,Go),
                                               (lizzieLet6_4QError_Bool_2,Go)] */
  logic [1:0] lizzieLet6_4QError_Bool_emitted;
  logic [1:0] lizzieLet6_4QError_Bool_done;
  assign lizzieLet6_4QError_Bool_1_d = (lizzieLet6_4QError_Bool_d[0] && (! lizzieLet6_4QError_Bool_emitted[0]));
  assign lizzieLet6_4QError_Bool_2_d = (lizzieLet6_4QError_Bool_d[0] && (! lizzieLet6_4QError_Bool_emitted[1]));
  assign lizzieLet6_4QError_Bool_done = (lizzieLet6_4QError_Bool_emitted | ({lizzieLet6_4QError_Bool_2_d[0],
                                                                             lizzieLet6_4QError_Bool_1_d[0]} & {lizzieLet6_4QError_Bool_2_r,
                                                                                                                lizzieLet6_4QError_Bool_1_r}));
  assign lizzieLet6_4QError_Bool_r = (& lizzieLet6_4QError_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Bool_emitted <= 2'd0;
    else
      lizzieLet6_4QError_Bool_emitted <= (lizzieLet6_4QError_Bool_r ? 2'd0 :
                                          lizzieLet6_4QError_Bool_done);
  
  /* dcon (Ty QTree_Nat,
      Dcon QError_Nat) : [(lizzieLet6_4QError_Bool_1,Go)] > (lizzieLet6_4QError_Bool_1QError_Nat,QTree_Nat) */
  assign lizzieLet6_4QError_Bool_1QError_Nat_d = QError_Nat_dc((& {lizzieLet6_4QError_Bool_1_d[0]}), lizzieLet6_4QError_Bool_1_d);
  assign {lizzieLet6_4QError_Bool_1_r} = {1 {(lizzieLet6_4QError_Bool_1QError_Nat_r && lizzieLet6_4QError_Bool_1QError_Nat_d[0])}};
  
  /* buf (Ty QTree_Nat) : (lizzieLet6_4QError_Bool_1QError_Nat,QTree_Nat) > (lizzieLet11_1_1_argbuf,QTree_Nat) */
  QTree_Nat_t lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d;
  logic lizzieLet6_4QError_Bool_1QError_Nat_bufchan_r;
  assign lizzieLet6_4QError_Bool_1QError_Nat_r = ((! lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d[0]) || lizzieLet6_4QError_Bool_1QError_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QError_Bool_1QError_Nat_r)
        lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d <= lizzieLet6_4QError_Bool_1QError_Nat_d;
  QTree_Nat_t lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf;
  assign lizzieLet6_4QError_Bool_1QError_Nat_bufchan_r = (! lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf[0] ? lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf :
                                     lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf[0]))
        lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf[0])))
        lizzieLet6_4QError_Bool_1QError_Nat_bufchan_buf <= lizzieLet6_4QError_Bool_1QError_Nat_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QError_Bool_2,Go) > (lizzieLet6_4QError_Bool_2_argbuf,Go) */
  Go_t lizzieLet6_4QError_Bool_2_bufchan_d;
  logic lizzieLet6_4QError_Bool_2_bufchan_r;
  assign lizzieLet6_4QError_Bool_2_r = ((! lizzieLet6_4QError_Bool_2_bufchan_d[0]) || lizzieLet6_4QError_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QError_Bool_2_r)
        lizzieLet6_4QError_Bool_2_bufchan_d <= lizzieLet6_4QError_Bool_2_d;
  Go_t lizzieLet6_4QError_Bool_2_bufchan_buf;
  assign lizzieLet6_4QError_Bool_2_bufchan_r = (! lizzieLet6_4QError_Bool_2_bufchan_buf[0]);
  assign lizzieLet6_4QError_Bool_2_argbuf_d = (lizzieLet6_4QError_Bool_2_bufchan_buf[0] ? lizzieLet6_4QError_Bool_2_bufchan_buf :
                                               lizzieLet6_4QError_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QError_Bool_2_argbuf_r && lizzieLet6_4QError_Bool_2_bufchan_buf[0]))
        lizzieLet6_4QError_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QError_Bool_2_argbuf_r) && (! lizzieLet6_4QError_Bool_2_bufchan_buf[0])))
        lizzieLet6_4QError_Bool_2_bufchan_buf <= lizzieLet6_4QError_Bool_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNode_Bool,Go) > (lizzieLet6_4QNode_Bool_1_argbuf,Go) */
  Go_t lizzieLet6_4QNode_Bool_bufchan_d;
  logic lizzieLet6_4QNode_Bool_bufchan_r;
  assign lizzieLet6_4QNode_Bool_r = ((! lizzieLet6_4QNode_Bool_bufchan_d[0]) || lizzieLet6_4QNode_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNode_Bool_r)
        lizzieLet6_4QNode_Bool_bufchan_d <= lizzieLet6_4QNode_Bool_d;
  Go_t lizzieLet6_4QNode_Bool_bufchan_buf;
  assign lizzieLet6_4QNode_Bool_bufchan_r = (! lizzieLet6_4QNode_Bool_bufchan_buf[0]);
  assign lizzieLet6_4QNode_Bool_1_argbuf_d = (lizzieLet6_4QNode_Bool_bufchan_buf[0] ? lizzieLet6_4QNode_Bool_bufchan_buf :
                                              lizzieLet6_4QNode_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNode_Bool_1_argbuf_r && lizzieLet6_4QNode_Bool_bufchan_buf[0]))
        lizzieLet6_4QNode_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNode_Bool_1_argbuf_r) && (! lizzieLet6_4QNode_Bool_bufchan_buf[0])))
        lizzieLet6_4QNode_Bool_bufchan_buf <= lizzieLet6_4QNode_Bool_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4QNone_Bool,Go) > [(lizzieLet6_4QNone_Bool_1,Go),
                                              (lizzieLet6_4QNone_Bool_2,Go)] */
  logic [1:0] lizzieLet6_4QNone_Bool_emitted;
  logic [1:0] lizzieLet6_4QNone_Bool_done;
  assign lizzieLet6_4QNone_Bool_1_d = (lizzieLet6_4QNone_Bool_d[0] && (! lizzieLet6_4QNone_Bool_emitted[0]));
  assign lizzieLet6_4QNone_Bool_2_d = (lizzieLet6_4QNone_Bool_d[0] && (! lizzieLet6_4QNone_Bool_emitted[1]));
  assign lizzieLet6_4QNone_Bool_done = (lizzieLet6_4QNone_Bool_emitted | ({lizzieLet6_4QNone_Bool_2_d[0],
                                                                           lizzieLet6_4QNone_Bool_1_d[0]} & {lizzieLet6_4QNone_Bool_2_r,
                                                                                                             lizzieLet6_4QNone_Bool_1_r}));
  assign lizzieLet6_4QNone_Bool_r = (& lizzieLet6_4QNone_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Bool_emitted <= 2'd0;
    else
      lizzieLet6_4QNone_Bool_emitted <= (lizzieLet6_4QNone_Bool_r ? 2'd0 :
                                         lizzieLet6_4QNone_Bool_done);
  
  /* dcon (Ty QTree_Nat,
      Dcon QNone_Nat) : [(lizzieLet6_4QNone_Bool_1,Go)] > (lizzieLet6_4QNone_Bool_1QNone_Nat,QTree_Nat) */
  assign lizzieLet6_4QNone_Bool_1QNone_Nat_d = QNone_Nat_dc((& {lizzieLet6_4QNone_Bool_1_d[0]}), lizzieLet6_4QNone_Bool_1_d);
  assign {lizzieLet6_4QNone_Bool_1_r} = {1 {(lizzieLet6_4QNone_Bool_1QNone_Nat_r && lizzieLet6_4QNone_Bool_1QNone_Nat_d[0])}};
  
  /* buf (Ty QTree_Nat) : (lizzieLet6_4QNone_Bool_1QNone_Nat,QTree_Nat) > (lizzieLet7_1_argbuf,QTree_Nat) */
  QTree_Nat_t lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d;
  logic lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_r;
  assign lizzieLet6_4QNone_Bool_1QNone_Nat_r = ((! lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d[0]) || lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QNone_Bool_1QNone_Nat_r)
        lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d <= lizzieLet6_4QNone_Bool_1QNone_Nat_d;
  QTree_Nat_t lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf;
  assign lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_r = (! lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf[0] ? lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf :
                                  lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf[0]))
        lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf[0])))
        lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_buf <= lizzieLet6_4QNone_Bool_1QNone_Nat_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNone_Bool_2,Go) > (lizzieLet6_4QNone_Bool_2_argbuf,Go) */
  Go_t lizzieLet6_4QNone_Bool_2_bufchan_d;
  logic lizzieLet6_4QNone_Bool_2_bufchan_r;
  assign lizzieLet6_4QNone_Bool_2_r = ((! lizzieLet6_4QNone_Bool_2_bufchan_d[0]) || lizzieLet6_4QNone_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNone_Bool_2_r)
        lizzieLet6_4QNone_Bool_2_bufchan_d <= lizzieLet6_4QNone_Bool_2_d;
  Go_t lizzieLet6_4QNone_Bool_2_bufchan_buf;
  assign lizzieLet6_4QNone_Bool_2_bufchan_r = (! lizzieLet6_4QNone_Bool_2_bufchan_buf[0]);
  assign lizzieLet6_4QNone_Bool_2_argbuf_d = (lizzieLet6_4QNone_Bool_2_bufchan_buf[0] ? lizzieLet6_4QNone_Bool_2_bufchan_buf :
                                              lizzieLet6_4QNone_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNone_Bool_2_argbuf_r && lizzieLet6_4QNone_Bool_2_bufchan_buf[0]))
        lizzieLet6_4QNone_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNone_Bool_2_argbuf_r) && (! lizzieLet6_4QNone_Bool_2_bufchan_buf[0])))
        lizzieLet6_4QNone_Bool_2_bufchan_buf <= lizzieLet6_4QNone_Bool_2_bufchan_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(lizzieLet6_4QNone_Bool_2_argbuf,Go),
                           (lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf,Go),
                           (es_0_1_1MyFalse_1_argbuf,Go),
                           (es_0_1_1MyTrue_2_argbuf,Go),
                           (lizzieLet6_4QError_Bool_2_argbuf,Go)] > (go_14_goMux_choice,C5) (go_14_goMux_data,Go) */
  logic [4:0] lizzieLet6_4QNone_Bool_2_argbuf_select_d;
  assign lizzieLet6_4QNone_Bool_2_argbuf_select_d = ((| lizzieLet6_4QNone_Bool_2_argbuf_select_q) ? lizzieLet6_4QNone_Bool_2_argbuf_select_q :
                                                     (lizzieLet6_4QNone_Bool_2_argbuf_d[0] ? 5'd1 :
                                                      (\lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_d [0] ? 5'd2 :
                                                       (es_0_1_1MyFalse_1_argbuf_d[0] ? 5'd4 :
                                                        (es_0_1_1MyTrue_2_argbuf_d[0] ? 5'd8 :
                                                         (lizzieLet6_4QError_Bool_2_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] lizzieLet6_4QNone_Bool_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Bool_2_argbuf_select_q <= 5'd0;
    else
      lizzieLet6_4QNone_Bool_2_argbuf_select_q <= (lizzieLet6_4QNone_Bool_2_argbuf_done ? 5'd0 :
                                                   lizzieLet6_4QNone_Bool_2_argbuf_select_d);
  logic [1:0] lizzieLet6_4QNone_Bool_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Bool_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_4QNone_Bool_2_argbuf_emit_q <= (lizzieLet6_4QNone_Bool_2_argbuf_done ? 2'd0 :
                                                 lizzieLet6_4QNone_Bool_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_4QNone_Bool_2_argbuf_emit_d;
  assign lizzieLet6_4QNone_Bool_2_argbuf_emit_d = (lizzieLet6_4QNone_Bool_2_argbuf_emit_q | ({go_14_goMux_choice_d[0],
                                                                                              go_14_goMux_data_d[0]} & {go_14_goMux_choice_r,
                                                                                                                        go_14_goMux_data_r}));
  logic lizzieLet6_4QNone_Bool_2_argbuf_done;
  assign lizzieLet6_4QNone_Bool_2_argbuf_done = (& lizzieLet6_4QNone_Bool_2_argbuf_emit_d);
  assign {lizzieLet6_4QError_Bool_2_argbuf_r,
          es_0_1_1MyTrue_2_argbuf_r,
          es_0_1_1MyFalse_1_argbuf_r,
          \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_r ,
          lizzieLet6_4QNone_Bool_2_argbuf_r} = (lizzieLet6_4QNone_Bool_2_argbuf_done ? lizzieLet6_4QNone_Bool_2_argbuf_select_d :
                                                5'd0);
  assign go_14_goMux_data_d = ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet6_4QNone_Bool_2_argbuf_d :
                               ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[0])) ? \lizzieLet29_3Lcall_main_map'_Bool_Nat0_1_argbuf_d  :
                                ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_1_1MyFalse_1_argbuf_d :
                                 ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[0])) ? es_0_1_1MyTrue_2_argbuf_d :
                                  ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[0])) ? lizzieLet6_4QError_Bool_2_argbuf_d :
                                   1'd0)))));
  assign go_14_goMux_choice_d = ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((lizzieLet6_4QNone_Bool_2_argbuf_select_d[4] && (! lizzieLet6_4QNone_Bool_2_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (lizzieLet6_4QVal_Bool,Go) > [(lizzieLet6_4QVal_Bool_1,Go),
                                             (lizzieLet6_4QVal_Bool_2,Go),
                                             (lizzieLet6_4QVal_Bool_3,Go)] */
  logic [2:0] lizzieLet6_4QVal_Bool_emitted;
  logic [2:0] lizzieLet6_4QVal_Bool_done;
  assign lizzieLet6_4QVal_Bool_1_d = (lizzieLet6_4QVal_Bool_d[0] && (! lizzieLet6_4QVal_Bool_emitted[0]));
  assign lizzieLet6_4QVal_Bool_2_d = (lizzieLet6_4QVal_Bool_d[0] && (! lizzieLet6_4QVal_Bool_emitted[1]));
  assign lizzieLet6_4QVal_Bool_3_d = (lizzieLet6_4QVal_Bool_d[0] && (! lizzieLet6_4QVal_Bool_emitted[2]));
  assign lizzieLet6_4QVal_Bool_done = (lizzieLet6_4QVal_Bool_emitted | ({lizzieLet6_4QVal_Bool_3_d[0],
                                                                         lizzieLet6_4QVal_Bool_2_d[0],
                                                                         lizzieLet6_4QVal_Bool_1_d[0]} & {lizzieLet6_4QVal_Bool_3_r,
                                                                                                          lizzieLet6_4QVal_Bool_2_r,
                                                                                                          lizzieLet6_4QVal_Bool_1_r}));
  assign lizzieLet6_4QVal_Bool_r = (& lizzieLet6_4QVal_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Bool_emitted <= 3'd0;
    else
      lizzieLet6_4QVal_Bool_emitted <= (lizzieLet6_4QVal_Bool_r ? 3'd0 :
                                        lizzieLet6_4QVal_Bool_done);
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Bool_1,Go) > (lizzieLet6_4QVal_Bool_1_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Bool_1_bufchan_d;
  logic lizzieLet6_4QVal_Bool_1_bufchan_r;
  assign lizzieLet6_4QVal_Bool_1_r = ((! lizzieLet6_4QVal_Bool_1_bufchan_d[0]) || lizzieLet6_4QVal_Bool_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Bool_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Bool_1_r)
        lizzieLet6_4QVal_Bool_1_bufchan_d <= lizzieLet6_4QVal_Bool_1_d;
  Go_t lizzieLet6_4QVal_Bool_1_bufchan_buf;
  assign lizzieLet6_4QVal_Bool_1_bufchan_r = (! lizzieLet6_4QVal_Bool_1_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Bool_1_argbuf_d = (lizzieLet6_4QVal_Bool_1_bufchan_buf[0] ? lizzieLet6_4QVal_Bool_1_bufchan_buf :
                                             lizzieLet6_4QVal_Bool_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Bool_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Bool_1_argbuf_r && lizzieLet6_4QVal_Bool_1_bufchan_buf[0]))
        lizzieLet6_4QVal_Bool_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Bool_1_argbuf_r) && (! lizzieLet6_4QVal_Bool_1_bufchan_buf[0])))
        lizzieLet6_4QVal_Bool_1_bufchan_buf <= lizzieLet6_4QVal_Bool_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTBool_Nat___MyBool,
      Dcon TupGo___MyDTBool_Nat___MyBool) : [(lizzieLet6_4QVal_Bool_1_argbuf,Go),
                                             (lizzieLet6_3QVal_Bool_1_argbuf,MyDTBool_Nat),
                                             (vacT_1_argbuf,MyBool)] > (applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1,TupGo___MyDTBool_Nat___MyBool) */
  assign applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d = TupGo___MyDTBool_Nat___MyBool_dc((& {lizzieLet6_4QVal_Bool_1_argbuf_d[0],
                                                                                                   lizzieLet6_3QVal_Bool_1_argbuf_d[0],
                                                                                                   vacT_1_argbuf_d[0]}), lizzieLet6_4QVal_Bool_1_argbuf_d, lizzieLet6_3QVal_Bool_1_argbuf_d, vacT_1_argbuf_d);
  assign {lizzieLet6_4QVal_Bool_1_argbuf_r,
          lizzieLet6_3QVal_Bool_1_argbuf_r,
          vacT_1_argbuf_r} = {3 {(applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_r && applyfnBool_Nat_5TupGo___MyDTBool_Nat___MyBool_1_d[0])}};
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Bool_2,Go) > (lizzieLet6_4QVal_Bool_2_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Bool_2_bufchan_d;
  logic lizzieLet6_4QVal_Bool_2_bufchan_r;
  assign lizzieLet6_4QVal_Bool_2_r = ((! lizzieLet6_4QVal_Bool_2_bufchan_d[0]) || lizzieLet6_4QVal_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Bool_2_r)
        lizzieLet6_4QVal_Bool_2_bufchan_d <= lizzieLet6_4QVal_Bool_2_d;
  Go_t lizzieLet6_4QVal_Bool_2_bufchan_buf;
  assign lizzieLet6_4QVal_Bool_2_bufchan_r = (! lizzieLet6_4QVal_Bool_2_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Bool_2_argbuf_d = (lizzieLet6_4QVal_Bool_2_bufchan_buf[0] ? lizzieLet6_4QVal_Bool_2_bufchan_buf :
                                             lizzieLet6_4QVal_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Bool_2_argbuf_r && lizzieLet6_4QVal_Bool_2_bufchan_buf[0]))
        lizzieLet6_4QVal_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Bool_2_argbuf_r) && (! lizzieLet6_4QVal_Bool_2_bufchan_buf[0])))
        lizzieLet6_4QVal_Bool_2_bufchan_buf <= lizzieLet6_4QVal_Bool_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTNat_Bool___Pointer_Nat,
      Dcon TupGo___MyDTNat_Bool___Pointer_Nat) : [(lizzieLet6_4QVal_Bool_2_argbuf,Go),
                                                  (lizzieLet6_5QVal_Bool_1_argbuf,MyDTNat_Bool),
                                                  (xacw_1_argbuf,Pointer_Nat)] > (applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1,TupGo___MyDTNat_Bool___Pointer_Nat) */
  assign applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d = TupGo___MyDTNat_Bool___Pointer_Nat_dc((& {lizzieLet6_4QVal_Bool_2_argbuf_d[0],
                                                                                                             lizzieLet6_5QVal_Bool_1_argbuf_d[0],
                                                                                                             xacw_1_argbuf_d[0]}), lizzieLet6_4QVal_Bool_2_argbuf_d, lizzieLet6_5QVal_Bool_1_argbuf_d, xacw_1_argbuf_d);
  assign {lizzieLet6_4QVal_Bool_2_argbuf_r,
          lizzieLet6_5QVal_Bool_1_argbuf_r,
          xacw_1_argbuf_r} = {3 {(applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_r && applyfnNat_Bool_5TupGo___MyDTNat_Bool___Pointer_Nat_1_d[0])}};
  
  /* demux (Ty QTree_Bool,
       Ty MyDTNat_Bool) : (lizzieLet6_5,QTree_Bool) (isZacQ_goMux_mux,MyDTNat_Bool) > [(_1,MyDTNat_Bool),
                                                                                       (lizzieLet6_5QVal_Bool,MyDTNat_Bool),
                                                                                       (lizzieLet6_5QNode_Bool,MyDTNat_Bool),
                                                                                       (_0,MyDTNat_Bool)] */
  logic [3:0] isZacQ_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && isZacQ_goMux_mux_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: isZacQ_goMux_mux_onehotd = 4'd1;
        2'd1: isZacQ_goMux_mux_onehotd = 4'd2;
        2'd2: isZacQ_goMux_mux_onehotd = 4'd4;
        2'd3: isZacQ_goMux_mux_onehotd = 4'd8;
        default: isZacQ_goMux_mux_onehotd = 4'd0;
      endcase
    else isZacQ_goMux_mux_onehotd = 4'd0;
  assign _1_d = isZacQ_goMux_mux_onehotd[0];
  assign lizzieLet6_5QVal_Bool_d = isZacQ_goMux_mux_onehotd[1];
  assign lizzieLet6_5QNode_Bool_d = isZacQ_goMux_mux_onehotd[2];
  assign _0_d = isZacQ_goMux_mux_onehotd[3];
  assign isZacQ_goMux_mux_r = (| (isZacQ_goMux_mux_onehotd & {_0_r,
                                                              lizzieLet6_5QNode_Bool_r,
                                                              lizzieLet6_5QVal_Bool_r,
                                                              _1_r}));
  assign lizzieLet6_5_r = isZacQ_goMux_mux_r;
  
  /* fork (Ty MyDTNat_Bool) : (lizzieLet6_5QNode_Bool,MyDTNat_Bool) > [(lizzieLet6_5QNode_Bool_1,MyDTNat_Bool),
                                                                  (lizzieLet6_5QNode_Bool_2,MyDTNat_Bool)] */
  logic [1:0] lizzieLet6_5QNode_Bool_emitted;
  logic [1:0] lizzieLet6_5QNode_Bool_done;
  assign lizzieLet6_5QNode_Bool_1_d = (lizzieLet6_5QNode_Bool_d[0] && (! lizzieLet6_5QNode_Bool_emitted[0]));
  assign lizzieLet6_5QNode_Bool_2_d = (lizzieLet6_5QNode_Bool_d[0] && (! lizzieLet6_5QNode_Bool_emitted[1]));
  assign lizzieLet6_5QNode_Bool_done = (lizzieLet6_5QNode_Bool_emitted | ({lizzieLet6_5QNode_Bool_2_d[0],
                                                                           lizzieLet6_5QNode_Bool_1_d[0]} & {lizzieLet6_5QNode_Bool_2_r,
                                                                                                             lizzieLet6_5QNode_Bool_1_r}));
  assign lizzieLet6_5QNode_Bool_r = (& lizzieLet6_5QNode_Bool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Bool_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Bool_emitted <= (lizzieLet6_5QNode_Bool_r ? 2'd0 :
                                         lizzieLet6_5QNode_Bool_done);
  
  /* buf (Ty MyDTNat_Bool) : (lizzieLet6_5QNode_Bool_2,MyDTNat_Bool) > (lizzieLet6_5QNode_Bool_2_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_2_bufchan_d;
  logic lizzieLet6_5QNode_Bool_2_bufchan_r;
  assign lizzieLet6_5QNode_Bool_2_r = ((! lizzieLet6_5QNode_Bool_2_bufchan_d[0]) || lizzieLet6_5QNode_Bool_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Bool_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Bool_2_r)
        lizzieLet6_5QNode_Bool_2_bufchan_d <= lizzieLet6_5QNode_Bool_2_d;
  MyDTNat_Bool_t lizzieLet6_5QNode_Bool_2_bufchan_buf;
  assign lizzieLet6_5QNode_Bool_2_bufchan_r = (! lizzieLet6_5QNode_Bool_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Bool_2_argbuf_d = (lizzieLet6_5QNode_Bool_2_bufchan_buf[0] ? lizzieLet6_5QNode_Bool_2_bufchan_buf :
                                              lizzieLet6_5QNode_Bool_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Bool_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Bool_2_argbuf_r && lizzieLet6_5QNode_Bool_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Bool_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Bool_2_argbuf_r) && (! lizzieLet6_5QNode_Bool_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Bool_2_bufchan_buf <= lizzieLet6_5QNode_Bool_2_bufchan_d;
  
  /* buf (Ty MyDTNat_Bool) : (lizzieLet6_5QVal_Bool,MyDTNat_Bool) > (lizzieLet6_5QVal_Bool_1_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t lizzieLet6_5QVal_Bool_bufchan_d;
  logic lizzieLet6_5QVal_Bool_bufchan_r;
  assign lizzieLet6_5QVal_Bool_r = ((! lizzieLet6_5QVal_Bool_bufchan_d[0]) || lizzieLet6_5QVal_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Bool_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Bool_r)
        lizzieLet6_5QVal_Bool_bufchan_d <= lizzieLet6_5QVal_Bool_d;
  MyDTNat_Bool_t lizzieLet6_5QVal_Bool_bufchan_buf;
  assign lizzieLet6_5QVal_Bool_bufchan_r = (! lizzieLet6_5QVal_Bool_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Bool_1_argbuf_d = (lizzieLet6_5QVal_Bool_bufchan_buf[0] ? lizzieLet6_5QVal_Bool_bufchan_buf :
                                             lizzieLet6_5QVal_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Bool_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Bool_1_argbuf_r && lizzieLet6_5QVal_Bool_bufchan_buf[0]))
        lizzieLet6_5QVal_Bool_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Bool_1_argbuf_r) && (! lizzieLet6_5QVal_Bool_bufchan_buf[0])))
        lizzieLet6_5QVal_Bool_bufchan_buf <= lizzieLet6_5QVal_Bool_bufchan_d;
  
  /* demux (Ty QTree_Bool,
       Ty Pointer_CTmain_map'_Bool_Nat) : (lizzieLet6_6,QTree_Bool) (sc_0_1_goMux_mux,Pointer_CTmain_map'_Bool_Nat) > [(lizzieLet6_6QNone_Bool,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                       (lizzieLet6_6QVal_Bool,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                       (lizzieLet6_6QNode_Bool,Pointer_CTmain_map'_Bool_Nat),
                                                                                                                       (lizzieLet6_6QError_Bool,Pointer_CTmain_map'_Bool_Nat)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_6QNone_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_6QVal_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_6QNode_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_6QError_Bool_d = {sc_0_1_goMux_mux_d[16:1],
                                      sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_6QError_Bool_r,
                                                              lizzieLet6_6QNode_Bool_r,
                                                              lizzieLet6_6QVal_Bool_r,
                                                              lizzieLet6_6QNone_Bool_r}));
  assign lizzieLet6_6_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (lizzieLet6_6QError_Bool,Pointer_CTmain_map'_Bool_Nat) > (lizzieLet6_6QError_Bool_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QError_Bool_bufchan_d;
  logic lizzieLet6_6QError_Bool_bufchan_r;
  assign lizzieLet6_6QError_Bool_r = ((! lizzieLet6_6QError_Bool_bufchan_d[0]) || lizzieLet6_6QError_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QError_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QError_Bool_r)
        lizzieLet6_6QError_Bool_bufchan_d <= lizzieLet6_6QError_Bool_d;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QError_Bool_bufchan_buf;
  assign lizzieLet6_6QError_Bool_bufchan_r = (! lizzieLet6_6QError_Bool_bufchan_buf[0]);
  assign lizzieLet6_6QError_Bool_1_argbuf_d = (lizzieLet6_6QError_Bool_bufchan_buf[0] ? lizzieLet6_6QError_Bool_bufchan_buf :
                                               lizzieLet6_6QError_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QError_Bool_1_argbuf_r && lizzieLet6_6QError_Bool_bufchan_buf[0]))
        lizzieLet6_6QError_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QError_Bool_1_argbuf_r) && (! lizzieLet6_6QError_Bool_bufchan_buf[0])))
        lizzieLet6_6QError_Bool_bufchan_buf <= lizzieLet6_6QError_Bool_bufchan_d;
  
  /* dcon (Ty CTmain_map'_Bool_Nat,
      Dcon Lcall_main_map'_Bool_Nat3) : [(lizzieLet6_6QNode_Bool,Pointer_CTmain_map'_Bool_Nat),
                                         (lizzieLet6_5QNode_Bool_1,MyDTNat_Bool),
                                         (lizzieLet6_3QNode_Bool_1,MyDTBool_Nat),
                                         (q1acU_destruct,Pointer_QTree_Bool),
                                         (q2acV_destruct,Pointer_QTree_Bool),
                                         (q3acW_destruct,Pointer_QTree_Bool)] > (lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3,CTmain_map'_Bool_Nat) */
  assign \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_d  = \Lcall_main_map'_Bool_Nat3_dc ((& {lizzieLet6_6QNode_Bool_d[0],
                                                                                                                                                                         lizzieLet6_5QNode_Bool_1_d[0],
                                                                                                                                                                         lizzieLet6_3QNode_Bool_1_d[0],
                                                                                                                                                                         q1acU_destruct_d[0],
                                                                                                                                                                         q2acV_destruct_d[0],
                                                                                                                                                                         q3acW_destruct_d[0]}), lizzieLet6_6QNode_Bool_d, lizzieLet6_5QNode_Bool_1_d, lizzieLet6_3QNode_Bool_1_d, q1acU_destruct_d, q2acV_destruct_d, q3acW_destruct_d);
  assign {lizzieLet6_6QNode_Bool_r,
          lizzieLet6_5QNode_Bool_1_r,
          lizzieLet6_3QNode_Bool_1_r,
          q1acU_destruct_r,
          q2acV_destruct_r,
          q3acW_destruct_r} = {6 {(\lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_r  && \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_d [0])}};
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3,CTmain_map'_Bool_Nat) > (lizzieLet10_1_argbuf,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d ;
  logic \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_r ;
  assign \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_r  = ((! \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d [0]) || \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d  <= {67'd0,
                                                                                                                                             1'd0};
    else
      if (\lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_r )
        \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d  <= \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_d ;
  \CTmain_map'_Bool_Nat_t  \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf ;
  assign \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_r  = (! \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf [0]);
  assign lizzieLet10_1_argbuf_d = (\lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf [0] ? \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf  :
                                   \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf  <= {67'd0,
                                                                                                                                               1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf [0]))
        \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf  <= {67'd0,
                                                                                                                                                 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf [0])))
        \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_buf  <= \lizzieLet6_6QNode_Bool_1lizzieLet6_5QNode_Bool_1lizzieLet6_3QNode_Bool_1q1acU_1q2acV_1q3acW_1Lcall_main_map'_Bool_Nat3_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (lizzieLet6_6QNone_Bool,Pointer_CTmain_map'_Bool_Nat) > (lizzieLet6_6QNone_Bool_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QNone_Bool_bufchan_d;
  logic lizzieLet6_6QNone_Bool_bufchan_r;
  assign lizzieLet6_6QNone_Bool_r = ((! lizzieLet6_6QNone_Bool_bufchan_d[0]) || lizzieLet6_6QNone_Bool_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNone_Bool_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_6QNone_Bool_r)
        lizzieLet6_6QNone_Bool_bufchan_d <= lizzieLet6_6QNone_Bool_d;
  \Pointer_CTmain_map'_Bool_Nat_t  lizzieLet6_6QNone_Bool_bufchan_buf;
  assign lizzieLet6_6QNone_Bool_bufchan_r = (! lizzieLet6_6QNone_Bool_bufchan_buf[0]);
  assign lizzieLet6_6QNone_Bool_1_argbuf_d = (lizzieLet6_6QNone_Bool_bufchan_buf[0] ? lizzieLet6_6QNone_Bool_bufchan_buf :
                                              lizzieLet6_6QNone_Bool_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_6QNone_Bool_1_argbuf_r && lizzieLet6_6QNone_Bool_bufchan_buf[0]))
        lizzieLet6_6QNone_Bool_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_6QNone_Bool_1_argbuf_r) && (! lizzieLet6_6QNone_Bool_bufchan_buf[0])))
        lizzieLet6_6QNone_Bool_bufchan_buf <= lizzieLet6_6QNone_Bool_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (m1ad9_goMux_mux,Pointer_QTree_Bool) > (m1ad9_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m1ad9_goMux_mux_bufchan_d;
  logic m1ad9_goMux_mux_bufchan_r;
  assign m1ad9_goMux_mux_r = ((! m1ad9_goMux_mux_bufchan_d[0]) || m1ad9_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad9_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1ad9_goMux_mux_r)
        m1ad9_goMux_mux_bufchan_d <= m1ad9_goMux_mux_d;
  Pointer_QTree_Bool_t m1ad9_goMux_mux_bufchan_buf;
  assign m1ad9_goMux_mux_bufchan_r = (! m1ad9_goMux_mux_bufchan_buf[0]);
  assign m1ad9_1_argbuf_d = (m1ad9_goMux_mux_bufchan_buf[0] ? m1ad9_goMux_mux_bufchan_buf :
                             m1ad9_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ad9_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1ad9_1_argbuf_r && m1ad9_goMux_mux_bufchan_buf[0]))
        m1ad9_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1ad9_1_argbuf_r) && (! m1ad9_goMux_mux_bufchan_buf[0])))
        m1ad9_goMux_mux_bufchan_buf <= m1ad9_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (m2ada_2_2,Pointer_QTree_Bool) > (m2ada_2_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2ada_2_2_bufchan_d;
  logic m2ada_2_2_bufchan_r;
  assign m2ada_2_2_r = ((! m2ada_2_2_bufchan_d[0]) || m2ada_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_2_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ada_2_2_r) m2ada_2_2_bufchan_d <= m2ada_2_2_d;
  Pointer_QTree_Bool_t m2ada_2_2_bufchan_buf;
  assign m2ada_2_2_bufchan_r = (! m2ada_2_2_bufchan_buf[0]);
  assign m2ada_2_2_argbuf_d = (m2ada_2_2_bufchan_buf[0] ? m2ada_2_2_bufchan_buf :
                               m2ada_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_2_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ada_2_2_argbuf_r && m2ada_2_2_bufchan_buf[0]))
        m2ada_2_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ada_2_2_argbuf_r) && (! m2ada_2_2_bufchan_buf[0])))
        m2ada_2_2_bufchan_buf <= m2ada_2_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2ada_2_destruct,Pointer_QTree_Bool) > [(m2ada_2_1,Pointer_QTree_Bool),
                                                                        (m2ada_2_2,Pointer_QTree_Bool)] */
  logic [1:0] m2ada_2_destruct_emitted;
  logic [1:0] m2ada_2_destruct_done;
  assign m2ada_2_1_d = {m2ada_2_destruct_d[16:1],
                        (m2ada_2_destruct_d[0] && (! m2ada_2_destruct_emitted[0]))};
  assign m2ada_2_2_d = {m2ada_2_destruct_d[16:1],
                        (m2ada_2_destruct_d[0] && (! m2ada_2_destruct_emitted[1]))};
  assign m2ada_2_destruct_done = (m2ada_2_destruct_emitted | ({m2ada_2_2_d[0],
                                                               m2ada_2_1_d[0]} & {m2ada_2_2_r,
                                                                                  m2ada_2_1_r}));
  assign m2ada_2_destruct_r = (& m2ada_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_2_destruct_emitted <= 2'd0;
    else
      m2ada_2_destruct_emitted <= (m2ada_2_destruct_r ? 2'd0 :
                                   m2ada_2_destruct_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2ada_3_2,Pointer_QTree_Bool) > (m2ada_3_2_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2ada_3_2_bufchan_d;
  logic m2ada_3_2_bufchan_r;
  assign m2ada_3_2_r = ((! m2ada_3_2_bufchan_d[0]) || m2ada_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_3_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ada_3_2_r) m2ada_3_2_bufchan_d <= m2ada_3_2_d;
  Pointer_QTree_Bool_t m2ada_3_2_bufchan_buf;
  assign m2ada_3_2_bufchan_r = (! m2ada_3_2_bufchan_buf[0]);
  assign m2ada_3_2_argbuf_d = (m2ada_3_2_bufchan_buf[0] ? m2ada_3_2_bufchan_buf :
                               m2ada_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_3_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ada_3_2_argbuf_r && m2ada_3_2_bufchan_buf[0]))
        m2ada_3_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ada_3_2_argbuf_r) && (! m2ada_3_2_bufchan_buf[0])))
        m2ada_3_2_bufchan_buf <= m2ada_3_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Bool) : (m2ada_3_destruct,Pointer_QTree_Bool) > [(m2ada_3_1,Pointer_QTree_Bool),
                                                                        (m2ada_3_2,Pointer_QTree_Bool)] */
  logic [1:0] m2ada_3_destruct_emitted;
  logic [1:0] m2ada_3_destruct_done;
  assign m2ada_3_1_d = {m2ada_3_destruct_d[16:1],
                        (m2ada_3_destruct_d[0] && (! m2ada_3_destruct_emitted[0]))};
  assign m2ada_3_2_d = {m2ada_3_destruct_d[16:1],
                        (m2ada_3_destruct_d[0] && (! m2ada_3_destruct_emitted[1]))};
  assign m2ada_3_destruct_done = (m2ada_3_destruct_emitted | ({m2ada_3_2_d[0],
                                                               m2ada_3_1_d[0]} & {m2ada_3_2_r,
                                                                                  m2ada_3_1_r}));
  assign m2ada_3_destruct_r = (& m2ada_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_3_destruct_emitted <= 2'd0;
    else
      m2ada_3_destruct_emitted <= (m2ada_3_destruct_r ? 2'd0 :
                                   m2ada_3_destruct_done);
  
  /* buf (Ty Pointer_QTree_Bool) : (m2ada_4_destruct,Pointer_QTree_Bool) > (m2ada_4_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t m2ada_4_destruct_bufchan_d;
  logic m2ada_4_destruct_bufchan_r;
  assign m2ada_4_destruct_r = ((! m2ada_4_destruct_bufchan_d[0]) || m2ada_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2ada_4_destruct_r)
        m2ada_4_destruct_bufchan_d <= m2ada_4_destruct_d;
  Pointer_QTree_Bool_t m2ada_4_destruct_bufchan_buf;
  assign m2ada_4_destruct_bufchan_r = (! m2ada_4_destruct_bufchan_buf[0]);
  assign m2ada_4_1_argbuf_d = (m2ada_4_destruct_bufchan_buf[0] ? m2ada_4_destruct_bufchan_buf :
                               m2ada_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ada_4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ada_4_1_argbuf_r && m2ada_4_destruct_bufchan_buf[0]))
        m2ada_4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ada_4_1_argbuf_r) && (! m2ada_4_destruct_bufchan_buf[0])))
        m2ada_4_destruct_bufchan_buf <= m2ada_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (macS_goMux_mux,Pointer_QTree_Bool) > (macS_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t macS_goMux_mux_bufchan_d;
  logic macS_goMux_mux_bufchan_r;
  assign macS_goMux_mux_r = ((! macS_goMux_mux_bufchan_d[0]) || macS_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macS_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (macS_goMux_mux_r) macS_goMux_mux_bufchan_d <= macS_goMux_mux_d;
  Pointer_QTree_Bool_t macS_goMux_mux_bufchan_buf;
  assign macS_goMux_mux_bufchan_r = (! macS_goMux_mux_bufchan_buf[0]);
  assign macS_1_argbuf_d = (macS_goMux_mux_bufchan_buf[0] ? macS_goMux_mux_bufchan_buf :
                            macS_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) macS_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((macS_1_argbuf_r && macS_goMux_mux_bufchan_buf[0]))
        macS_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! macS_1_argbuf_r) && (! macS_goMux_mux_bufchan_buf[0])))
        macS_goMux_mux_bufchan_buf <= macS_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (mad1_goMux_mux,Pointer_QTree_Bool) > (mad1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t mad1_goMux_mux_bufchan_d;
  logic mad1_goMux_mux_bufchan_r;
  assign mad1_goMux_mux_r = ((! mad1_goMux_mux_bufchan_d[0]) || mad1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mad1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (mad1_goMux_mux_r) mad1_goMux_mux_bufchan_d <= mad1_goMux_mux_d;
  Pointer_QTree_Bool_t mad1_goMux_mux_bufchan_buf;
  assign mad1_goMux_mux_bufchan_r = (! mad1_goMux_mux_bufchan_buf[0]);
  assign mad1_1_argbuf_d = (mad1_goMux_mux_bufchan_buf[0] ? mad1_goMux_mux_bufchan_buf :
                            mad1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mad1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mad1_1_argbuf_r && mad1_goMux_mux_bufchan_buf[0]))
        mad1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mad1_1_argbuf_r) && (! mad1_goMux_mux_bufchan_buf[0])))
        mad1_goMux_mux_bufchan_buf <= mad1_goMux_mux_bufchan_d;
  
  /* destruct (Ty TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool,
          Dcon TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool) : (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1,TupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool) > [(main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11,Go),
                                                                                                                                                                                                                      (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1,MyDTNat_Bool),
                                                                                                                                                                                                                      (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1,MyDTBool_Nat),
                                                                                                                                                                                                                      (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1,Pointer_QTree_Bool)] */
  logic [3:0] \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted ;
  logic [3:0] \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_done ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_d  = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted [0]));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_d  = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted [1]));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_d  = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted [2]));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_d  = {\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [16:1],
                                                                                                 (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted [3]))};
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_done  = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted  | ({\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_d [0],
                                                                                                                                                                                           \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_d [0],
                                                                                                                                                                                           \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_d [0],
                                                                                                                                                                                           \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_d [0]} & {\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_r ,
                                                                                                                                                                                                                                                                                      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_r }));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_r  = (& \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted  <= 4'd0;
    else
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_emitted  <= (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_r  ? 4'd0 :
                                                                                                 \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Bool_1_done );
  
  /* buf (Ty MyDTBool_Nat) : (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1,MyDTBool_Nat) > (gacR_1_1_argbuf,MyDTBool_Nat) */
  MyDTBool_Nat_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_r ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_r  = ((! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d [0]) || \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_r )
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_d ;
  MyDTBool_Nat_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_r  = (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf [0]);
  assign gacR_1_1_argbuf_d = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf [0] ? \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf  :
                              \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf  <= 1'd0;
    else
      if ((gacR_1_1_argbuf_r && \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf [0]))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf  <= 1'd0;
      else if (((! gacR_1_1_argbuf_r) && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf [0])))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_buf  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolgacR_1_bufchan_d ;
  
  /* fork (Ty Go) : (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11,Go) > [(go_11_1,Go),
                                                                                                       (go_11_2,Go)] */
  logic [1:0] \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted ;
  logic [1:0] \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_done ;
  assign go_11_1_d = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted [0]));
  assign go_11_2_d = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_d [0] && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted [1]));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_done  = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted  | ({go_11_2_d[0],
                                                                                                                                                                                                 go_11_1_d[0]} & {go_11_2_r,
                                                                                                                                                                                                                  go_11_1_r}));
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_r  = (& \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted  <= 2'd0;
    else
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_emitted  <= (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_r  ? 2'd0 :
                                                                                                    \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_Boolgo_11_done );
  
  /* buf (Ty MyDTNat_Bool) : (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1,MyDTNat_Bool) > (isZacQ_1_1_argbuf,MyDTNat_Bool) */
  MyDTNat_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_r ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_r  = ((! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d [0]) || \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d  <= 1'd0;
    else
      if (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_r )
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_d ;
  MyDTNat_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_r  = (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf [0]);
  assign isZacQ_1_1_argbuf_d = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf [0] ? \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf  :
                                \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacQ_1_1_argbuf_r && \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf [0]))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf  <= 1'd0;
      else if (((! isZacQ_1_1_argbuf_r) && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf [0])))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_buf  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolisZacQ_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1,Pointer_QTree_Bool) > (macS_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d ;
  logic \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_r ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_r  = ((! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d [0]) || \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d  <= {16'd0,
                                                                                                       1'd0};
    else
      if (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_r )
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_d ;
  Pointer_QTree_Bool_t \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf ;
  assign \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_r  = (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf [0]);
  assign macS_1_1_argbuf_d = (\main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf [0] ? \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf  :
                              \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf  <= {16'd0,
                                                                                                         1'd0};
    else
      if ((macS_1_1_argbuf_r && \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf [0]))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf  <= {16'd0,
                                                                                                           1'd0};
      else if (((! macS_1_1_argbuf_r) && (! \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf [0])))
        \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_buf  <= \main_map'_Bool_NatTupGo___MyDTNat_Bool___MyDTBool_Nat___Pointer_QTree_BoolmacS_1_bufchan_d ;
  
  /* sink (Ty Pointer_QTree_Nat) : (main_map'_Bool_Nat_resbuf,Pointer_QTree_Nat) > */
  assign {\main_map'_Bool_Nat_resbuf_r ,
          \main_map'_Bool_Nat_resbuf_dout } = {\main_map'_Bool_Nat_resbuf_rout ,
                                               \main_map'_Bool_Nat_resbuf_d };
  
  /* destruct (Ty TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool,
          Dcon TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1,TupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool) > [(map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12,Go),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1,MyDTBool_Bool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1,MyDTBool_Bool_Bool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1,MyBool),
                                                                                                                                                                                                                                                                              (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1,Pointer_QTree_Bool)] */
  logic [4:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted ;
  logic [4:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [0]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [1]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [2]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_d  = {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [1:1],
                                                                                                                          (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [3]))};
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_d  = {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [17:2],
                                                                                                                         (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted [4]))};
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  | ({\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_d [0],
                                                                                                                                                                                                                                           \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_d [0]} & {\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_r ,
                                                                                                                                                                                                                                                                                                                                                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_r ,
                                                                                                                                                                                                                                                                                                                                                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_r ,
                                                                                                                                                                                                                                                                                                                                                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_r ,
                                                                                                                                                                                                                                                                                                                                                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_r }));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  = (& \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  <= 5'd0;
    else
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_emitted  <= (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_r  ? 5'd0 :
                                                                                                                         \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Bool_1_done );
  
  /* buf (Ty MyDTBool_Bool_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1,MyDTBool_Bool_Bool) > (gacZ_1_1_argbuf,MyDTBool_Bool_Bool) */
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_d ;
  MyDTBool_Bool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf [0]);
  assign gacZ_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf  :
                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf  <= 1'd0;
    else
      if ((gacZ_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf  <= 1'd0;
      else if (((! gacZ_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolgacZ_1_bufchan_d ;
  
  /* fork (Ty Go) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12,Go) > [(go_12_1,Go),
                                                                                                                               (go_12_2,Go)] */
  logic [1:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted ;
  logic [1:0] \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_done ;
  assign go_12_1_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted [0]));
  assign go_12_2_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_d [0] && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted [1]));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_done  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted  | ({go_12_2_d[0],
                                                                                                                                                                                                                                                 go_12_1_d[0]} & {go_12_2_r,
                                                                                                                                                                                                                                                                  go_12_1_r}));
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_r  = (& \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted  <= 2'd0;
    else
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_emitted  <= (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_r  ? 2'd0 :
                                                                                                                            \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolgo_12_done );
  
  /* buf (Ty MyDTBool_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1,MyDTBool_Bool) > (isZacY_1_1_argbuf,MyDTBool_Bool) */
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d  <= 1'd0;
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_d ;
  MyDTBool_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf [0]);
  assign isZacY_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf  :
                                \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf  <= 1'd0;
    else
      if ((isZacY_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf  <= 1'd0;
      else if (((! isZacY_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_BoolisZacY_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1,Pointer_QTree_Bool) > (mad1_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d  <= {16'd0,
                                                                                                                               1'd0};
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_d ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf [0]);
  assign mad1_1_1_argbuf_d = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf  :
                              \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf  <= {16'd0,
                                                                                                                                 1'd0};
    else
      if ((mad1_1_1_argbuf_r && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf  <= {16'd0,
                                                                                                                                   1'd0};
      else if (((! mad1_1_1_argbuf_r) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolmad1_1_bufchan_d ;
  
  /* buf (Ty MyBool) : (map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1,MyBool) > (v'ad0_1_1_argbuf,MyBool) */
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d ;
  logic \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_r ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_r  = ((! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d [0]) || \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d  <= {1'd0,
                                                                                                                                1'd0};
    else
      if (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_r )
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_d ;
  MyBool_t \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf ;
  assign \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_r  = (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf [0]);
  assign \v'ad0_1_1_argbuf_d  = (\map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf [0] ? \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf  :
                                 \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf  <= {1'd0,
                                                                                                                                  1'd0};
    else
      if ((\v'ad0_1_1_argbuf_r  && \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf [0]))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf  <= {1'd0,
                                                                                                                                    1'd0};
      else if (((! \v'ad0_1_1_argbuf_r ) && (! \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf [0])))
        \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_buf  <= \map''_map''_Bool_Bool_BoolTupGo___MyDTBool_Bool___MyDTBool_Bool_Bool___MyBool___Pointer_QTree_Boolv'ad0_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (map''_map''_Bool_Bool_Bool_resbuf,Pointer_QTree_Bool) > (lizzieLet12_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d ;
  logic \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r ;
  assign \map''_map''_Bool_Bool_Bool_resbuf_r  = ((! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d [0]) || \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\map''_map''_Bool_Bool_Bool_resbuf_r )
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d  <= \map''_map''_Bool_Bool_Bool_resbuf_d ;
  Pointer_QTree_Bool_t \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf ;
  assign \map''_map''_Bool_Bool_Bool_resbuf_bufchan_r  = (! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0]);
  assign lizzieLet12_1_argbuf_d = (\map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0] ? \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  :
                                   \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0]))
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf [0])))
        \map''_map''_Bool_Bool_Bool_resbuf_bufchan_buf  <= \map''_map''_Bool_Bool_Bool_resbuf_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1acU_3_destruct,Pointer_QTree_Bool) > (q1acU_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1acU_3_destruct_bufchan_d;
  logic q1acU_3_destruct_bufchan_r;
  assign q1acU_3_destruct_r = ((! q1acU_3_destruct_bufchan_d[0]) || q1acU_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acU_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1acU_3_destruct_r)
        q1acU_3_destruct_bufchan_d <= q1acU_3_destruct_d;
  Pointer_QTree_Bool_t q1acU_3_destruct_bufchan_buf;
  assign q1acU_3_destruct_bufchan_r = (! q1acU_3_destruct_bufchan_buf[0]);
  assign q1acU_3_1_argbuf_d = (q1acU_3_destruct_bufchan_buf[0] ? q1acU_3_destruct_bufchan_buf :
                               q1acU_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1acU_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1acU_3_1_argbuf_r && q1acU_3_destruct_bufchan_buf[0]))
        q1acU_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1acU_3_1_argbuf_r) && (! q1acU_3_destruct_bufchan_buf[0])))
        q1acU_3_destruct_bufchan_buf <= q1acU_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1ad3_3_destruct,Pointer_QTree_Bool) > (q1ad3_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1ad3_3_destruct_bufchan_d;
  logic q1ad3_3_destruct_bufchan_r;
  assign q1ad3_3_destruct_r = ((! q1ad3_3_destruct_bufchan_d[0]) || q1ad3_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ad3_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ad3_3_destruct_r)
        q1ad3_3_destruct_bufchan_d <= q1ad3_3_destruct_d;
  Pointer_QTree_Bool_t q1ad3_3_destruct_bufchan_buf;
  assign q1ad3_3_destruct_bufchan_r = (! q1ad3_3_destruct_bufchan_buf[0]);
  assign q1ad3_3_1_argbuf_d = (q1ad3_3_destruct_bufchan_buf[0] ? q1ad3_3_destruct_bufchan_buf :
                               q1ad3_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ad3_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ad3_3_1_argbuf_r && q1ad3_3_destruct_bufchan_buf[0]))
        q1ad3_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ad3_3_1_argbuf_r) && (! q1ad3_3_destruct_bufchan_buf[0])))
        q1ad3_3_destruct_bufchan_buf <= q1ad3_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q1adc_3_destruct,Pointer_QTree_Bool) > (q1adc_3_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q1adc_3_destruct_bufchan_d;
  logic q1adc_3_destruct_bufchan_r;
  assign q1adc_3_destruct_r = ((! q1adc_3_destruct_bufchan_d[0]) || q1adc_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1adc_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1adc_3_destruct_r)
        q1adc_3_destruct_bufchan_d <= q1adc_3_destruct_d;
  Pointer_QTree_Bool_t q1adc_3_destruct_bufchan_buf;
  assign q1adc_3_destruct_bufchan_r = (! q1adc_3_destruct_bufchan_buf[0]);
  assign q1adc_3_1_argbuf_d = (q1adc_3_destruct_bufchan_buf[0] ? q1adc_3_destruct_bufchan_buf :
                               q1adc_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1adc_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1adc_3_1_argbuf_r && q1adc_3_destruct_bufchan_buf[0]))
        q1adc_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1adc_3_1_argbuf_r) && (! q1adc_3_destruct_bufchan_buf[0])))
        q1adc_3_destruct_bufchan_buf <= q1adc_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2acV_2_destruct,Pointer_QTree_Bool) > (q2acV_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2acV_2_destruct_bufchan_d;
  logic q2acV_2_destruct_bufchan_r;
  assign q2acV_2_destruct_r = ((! q2acV_2_destruct_bufchan_d[0]) || q2acV_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acV_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2acV_2_destruct_r)
        q2acV_2_destruct_bufchan_d <= q2acV_2_destruct_d;
  Pointer_QTree_Bool_t q2acV_2_destruct_bufchan_buf;
  assign q2acV_2_destruct_bufchan_r = (! q2acV_2_destruct_bufchan_buf[0]);
  assign q2acV_2_1_argbuf_d = (q2acV_2_destruct_bufchan_buf[0] ? q2acV_2_destruct_bufchan_buf :
                               q2acV_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2acV_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2acV_2_1_argbuf_r && q2acV_2_destruct_bufchan_buf[0]))
        q2acV_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2acV_2_1_argbuf_r) && (! q2acV_2_destruct_bufchan_buf[0])))
        q2acV_2_destruct_bufchan_buf <= q2acV_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2ad4_2_destruct,Pointer_QTree_Bool) > (q2ad4_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2ad4_2_destruct_bufchan_d;
  logic q2ad4_2_destruct_bufchan_r;
  assign q2ad4_2_destruct_r = ((! q2ad4_2_destruct_bufchan_d[0]) || q2ad4_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ad4_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2ad4_2_destruct_r)
        q2ad4_2_destruct_bufchan_d <= q2ad4_2_destruct_d;
  Pointer_QTree_Bool_t q2ad4_2_destruct_bufchan_buf;
  assign q2ad4_2_destruct_bufchan_r = (! q2ad4_2_destruct_bufchan_buf[0]);
  assign q2ad4_2_1_argbuf_d = (q2ad4_2_destruct_bufchan_buf[0] ? q2ad4_2_destruct_bufchan_buf :
                               q2ad4_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ad4_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2ad4_2_1_argbuf_r && q2ad4_2_destruct_bufchan_buf[0]))
        q2ad4_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2ad4_2_1_argbuf_r) && (! q2ad4_2_destruct_bufchan_buf[0])))
        q2ad4_2_destruct_bufchan_buf <= q2ad4_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q2add_2_destruct,Pointer_QTree_Bool) > (q2add_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q2add_2_destruct_bufchan_d;
  logic q2add_2_destruct_bufchan_r;
  assign q2add_2_destruct_r = ((! q2add_2_destruct_bufchan_d[0]) || q2add_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2add_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2add_2_destruct_r)
        q2add_2_destruct_bufchan_d <= q2add_2_destruct_d;
  Pointer_QTree_Bool_t q2add_2_destruct_bufchan_buf;
  assign q2add_2_destruct_bufchan_r = (! q2add_2_destruct_bufchan_buf[0]);
  assign q2add_2_1_argbuf_d = (q2add_2_destruct_bufchan_buf[0] ? q2add_2_destruct_bufchan_buf :
                               q2add_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2add_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2add_2_1_argbuf_r && q2add_2_destruct_bufchan_buf[0]))
        q2add_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2add_2_1_argbuf_r) && (! q2add_2_destruct_bufchan_buf[0])))
        q2add_2_destruct_bufchan_buf <= q2add_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3acW_1_destruct,Pointer_QTree_Bool) > (q3acW_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3acW_1_destruct_bufchan_d;
  logic q3acW_1_destruct_bufchan_r;
  assign q3acW_1_destruct_r = ((! q3acW_1_destruct_bufchan_d[0]) || q3acW_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acW_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3acW_1_destruct_r)
        q3acW_1_destruct_bufchan_d <= q3acW_1_destruct_d;
  Pointer_QTree_Bool_t q3acW_1_destruct_bufchan_buf;
  assign q3acW_1_destruct_bufchan_r = (! q3acW_1_destruct_bufchan_buf[0]);
  assign q3acW_1_1_argbuf_d = (q3acW_1_destruct_bufchan_buf[0] ? q3acW_1_destruct_bufchan_buf :
                               q3acW_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3acW_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3acW_1_1_argbuf_r && q3acW_1_destruct_bufchan_buf[0]))
        q3acW_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3acW_1_1_argbuf_r) && (! q3acW_1_destruct_bufchan_buf[0])))
        q3acW_1_destruct_bufchan_buf <= q3acW_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3ad5_1_destruct,Pointer_QTree_Bool) > (q3ad5_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3ad5_1_destruct_bufchan_d;
  logic q3ad5_1_destruct_bufchan_r;
  assign q3ad5_1_destruct_r = ((! q3ad5_1_destruct_bufchan_d[0]) || q3ad5_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad5_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ad5_1_destruct_r)
        q3ad5_1_destruct_bufchan_d <= q3ad5_1_destruct_d;
  Pointer_QTree_Bool_t q3ad5_1_destruct_bufchan_buf;
  assign q3ad5_1_destruct_bufchan_r = (! q3ad5_1_destruct_bufchan_buf[0]);
  assign q3ad5_1_1_argbuf_d = (q3ad5_1_destruct_bufchan_buf[0] ? q3ad5_1_destruct_bufchan_buf :
                               q3ad5_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ad5_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ad5_1_1_argbuf_r && q3ad5_1_destruct_bufchan_buf[0]))
        q3ad5_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ad5_1_1_argbuf_r) && (! q3ad5_1_destruct_bufchan_buf[0])))
        q3ad5_1_destruct_bufchan_buf <= q3ad5_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q3ade_1_destruct,Pointer_QTree_Bool) > (q3ade_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q3ade_1_destruct_bufchan_d;
  logic q3ade_1_destruct_bufchan_r;
  assign q3ade_1_destruct_r = ((! q3ade_1_destruct_bufchan_d[0]) || q3ade_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ade_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ade_1_destruct_r)
        q3ade_1_destruct_bufchan_d <= q3ade_1_destruct_d;
  Pointer_QTree_Bool_t q3ade_1_destruct_bufchan_buf;
  assign q3ade_1_destruct_bufchan_r = (! q3ade_1_destruct_bufchan_buf[0]);
  assign q3ade_1_1_argbuf_d = (q3ade_1_destruct_bufchan_buf[0] ? q3ade_1_destruct_bufchan_buf :
                               q3ade_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ade_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ade_1_1_argbuf_r && q3ade_1_destruct_bufchan_buf[0]))
        q3ade_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ade_1_1_argbuf_r) && (! q3ade_1_destruct_bufchan_buf[0])))
        q3ade_1_destruct_bufchan_buf <= q3ade_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4acX_destruct,Pointer_QTree_Bool) > (q4acX_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4acX_destruct_bufchan_d;
  logic q4acX_destruct_bufchan_r;
  assign q4acX_destruct_r = ((! q4acX_destruct_bufchan_d[0]) || q4acX_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acX_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4acX_destruct_r) q4acX_destruct_bufchan_d <= q4acX_destruct_d;
  Pointer_QTree_Bool_t q4acX_destruct_bufchan_buf;
  assign q4acX_destruct_bufchan_r = (! q4acX_destruct_bufchan_buf[0]);
  assign q4acX_1_argbuf_d = (q4acX_destruct_bufchan_buf[0] ? q4acX_destruct_bufchan_buf :
                             q4acX_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4acX_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4acX_1_argbuf_r && q4acX_destruct_bufchan_buf[0]))
        q4acX_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4acX_1_argbuf_r) && (! q4acX_destruct_bufchan_buf[0])))
        q4acX_destruct_bufchan_buf <= q4acX_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4ad6_destruct,Pointer_QTree_Bool) > (q4ad6_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4ad6_destruct_bufchan_d;
  logic q4ad6_destruct_bufchan_r;
  assign q4ad6_destruct_r = ((! q4ad6_destruct_bufchan_d[0]) || q4ad6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ad6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4ad6_destruct_r) q4ad6_destruct_bufchan_d <= q4ad6_destruct_d;
  Pointer_QTree_Bool_t q4ad6_destruct_bufchan_buf;
  assign q4ad6_destruct_bufchan_r = (! q4ad6_destruct_bufchan_buf[0]);
  assign q4ad6_1_argbuf_d = (q4ad6_destruct_bufchan_buf[0] ? q4ad6_destruct_bufchan_buf :
                             q4ad6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ad6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4ad6_1_argbuf_r && q4ad6_destruct_bufchan_buf[0]))
        q4ad6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4ad6_1_argbuf_r) && (! q4ad6_destruct_bufchan_buf[0])))
        q4ad6_destruct_bufchan_buf <= q4ad6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (q4adf_destruct,Pointer_QTree_Bool) > (q4adf_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t q4adf_destruct_bufchan_d;
  logic q4adf_destruct_bufchan_r;
  assign q4adf_destruct_r = ((! q4adf_destruct_bufchan_d[0]) || q4adf_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4adf_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4adf_destruct_r) q4adf_destruct_bufchan_d <= q4adf_destruct_d;
  Pointer_QTree_Bool_t q4adf_destruct_bufchan_buf;
  assign q4adf_destruct_bufchan_r = (! q4adf_destruct_bufchan_buf[0]);
  assign q4adf_1_argbuf_d = (q4adf_destruct_bufchan_buf[0] ? q4adf_destruct_bufchan_buf :
                             q4adf_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4adf_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4adf_1_argbuf_r && q4adf_destruct_bufchan_buf[0]))
        q4adf_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4adf_1_argbuf_r) && (! q4adf_destruct_bufchan_buf[0])))
        q4adf_destruct_bufchan_buf <= q4adf_destruct_bufchan_d;
  
  /* buf (Ty CTkron_kron_Bool_Bool_Bool) : (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf,CTkron_kron_Bool_Bool_Bool) > (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb,CTkron_kron_Bool_Bool_Bool) */
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r = ((! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d <= {83'd0,
                                                                            1'd0};
    else
      if (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_r)
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d <= readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_d;
  CTkron_kron_Bool_Bool_Bool_t readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_r = (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d = (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf :
                                                                          readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= {83'd0,
                                                                              1'd0};
    else
      if ((readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r && readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= {83'd0,
                                                                                1'd0};
      else if (((! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r) && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_buf <= readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CTkron_kron_Bool_Bool_Bool) : (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb,CTkron_kron_Bool_Bool_Bool) > [(lizzieLet24_1,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet24_2,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet24_3,CTkron_kron_Bool_Bool_Bool),
                                                                                                                                   (lizzieLet24_4,CTkron_kron_Bool_Bool_Bool)] */
  logic [3:0] readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet24_1_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet24_2_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet24_3_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet24_4_d = {readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[83:1],
                            (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done = (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet24_4_d[0],
                                                                                                                                                     lizzieLet24_3_d[0],
                                                                                                                                                     lizzieLet24_2_d[0],
                                                                                                                                                     lizzieLet24_1_d[0]} & {lizzieLet24_4_r,
                                                                                                                                                                            lizzieLet24_3_r,
                                                                                                                                                                            lizzieLet24_2_r,
                                                                                                                                                                            lizzieLet24_1_r}));
  assign readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r = (& readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                                              readPointer_CTkron_kron_Bool_Bool_Boolscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTmain_map'_Bool_Nat) : (readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf,CTmain_map'_Bool_Nat) > (readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb,CTmain_map'_Bool_Nat) */
  \CTmain_map'_Bool_Nat_t  \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_r  = ((! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d  <= {67'd0,
                                                                          1'd0};
    else
      if (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_r )
        \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_d ;
  \CTmain_map'_Bool_Nat_t  \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf  :
                                                                        \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                            1'd0};
    else
      if ((\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf  <= {67'd0,
                                                                              1'd0};
      else if (((! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmain_map'_Bool_Nat) : (readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb,CTmain_map'_Bool_Nat) > [(lizzieLet29_1,CTmain_map'_Bool_Nat),
                                                                                                                   (lizzieLet29_2,CTmain_map'_Bool_Nat),
                                                                                                                   (lizzieLet29_3,CTmain_map'_Bool_Nat),
                                                                                                                   (lizzieLet29_4,CTmain_map'_Bool_Nat)] */
  logic [3:0] \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet29_1_d = {\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet29_2_d = {\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet29_3_d = {\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet29_4_d = {\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [67:1],
                            (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet29_4_d[0],
                                                                                                                                                 lizzieLet29_3_d[0],
                                                                                                                                                 lizzieLet29_2_d[0],
                                                                                                                                                 lizzieLet29_1_d[0]} & {lizzieLet29_4_r,
                                                                                                                                                                        lizzieLet29_3_r,
                                                                                                                                                                        lizzieLet29_2_r,
                                                                                                                                                                        lizzieLet29_1_r}));
  assign \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                            \readPointer_CTmain_map'_Bool_Natscfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTmap''_map''_Bool_Bool_Bool) : (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf,CTmap''_map''_Bool_Bool_Bool) > (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb,CTmap''_map''_Bool_Bool_Bool) */
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  logic \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r ;
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r  = ((! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d [0]) || \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d  <= {68'd0,
                                                                                  1'd0};
    else
      if (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_r )
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d  <= \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_d ;
  \CTmap''_map''_Bool_Bool_Bool_t  \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf ;
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_r  = (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d  = (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0] ? \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  :
                                                                                \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {68'd0,
                                                                                    1'd0};
    else
      if ((\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  && \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0]))
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= {68'd0,
                                                                                      1'd0};
      else if (((! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r ) && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf [0])))
        \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_buf  <= \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTmap''_map''_Bool_Bool_Bool) : (readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb,CTmap''_map''_Bool_Bool_Bool) > [(lizzieLet34_1,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet34_2,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet34_3,CTmap''_map''_Bool_Bool_Bool),
                                                                                                                                           (lizzieLet34_4,CTmap''_map''_Bool_Bool_Bool)] */
  logic [3:0] \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done ;
  assign lizzieLet34_1_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet34_2_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet34_3_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet34_4_d = {\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [68:1],
                            (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_d [0] && (! \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done  = (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  | ({lizzieLet34_4_d[0],
                                                                                                                                                                 lizzieLet34_3_d[0],
                                                                                                                                                                 lizzieLet34_2_d[0],
                                                                                                                                                                 lizzieLet34_1_d[0]} & {lizzieLet34_4_r,
                                                                                                                                                                                        lizzieLet34_3_r,
                                                                                                                                                                                        lizzieLet34_2_r,
                                                                                                                                                                                        lizzieLet34_1_r}));
  assign \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  = (& \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_emitted  <= (\readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_r  ? 4'd0 :
                                                                                    \readPointer_CTmap''_map''_Bool_Bool_Boolscfarg_0_2_1_argbuf_rwb_done );
  
  /* buf (Ty Nat) : (readPointer_Natxadg_1_argbuf,Nat) > (readPointer_Natxadg_1_argbuf_rwb,Nat) */
  Nat_t readPointer_Natxadg_1_argbuf_bufchan_d;
  logic readPointer_Natxadg_1_argbuf_bufchan_r;
  assign readPointer_Natxadg_1_argbuf_r = ((! readPointer_Natxadg_1_argbuf_bufchan_d[0]) || readPointer_Natxadg_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_Natxadg_1_argbuf_bufchan_d <= {17'd0, 1'd0};
    else
      if (readPointer_Natxadg_1_argbuf_r)
        readPointer_Natxadg_1_argbuf_bufchan_d <= readPointer_Natxadg_1_argbuf_d;
  Nat_t readPointer_Natxadg_1_argbuf_bufchan_buf;
  assign readPointer_Natxadg_1_argbuf_bufchan_r = (! readPointer_Natxadg_1_argbuf_bufchan_buf[0]);
  assign readPointer_Natxadg_1_argbuf_rwb_d = (readPointer_Natxadg_1_argbuf_bufchan_buf[0] ? readPointer_Natxadg_1_argbuf_bufchan_buf :
                                               readPointer_Natxadg_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_Natxadg_1_argbuf_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((readPointer_Natxadg_1_argbuf_rwb_r && readPointer_Natxadg_1_argbuf_bufchan_buf[0]))
        readPointer_Natxadg_1_argbuf_bufchan_buf <= {17'd0, 1'd0};
      else if (((! readPointer_Natxadg_1_argbuf_rwb_r) && (! readPointer_Natxadg_1_argbuf_bufchan_buf[0])))
        readPointer_Natxadg_1_argbuf_bufchan_buf <= readPointer_Natxadg_1_argbuf_bufchan_d;
  
  /* fork (Ty Nat) : (readPointer_Natxadg_1_argbuf_rwb,Nat) > [(lizzieLet18_1,Nat),
                                                          (lizzieLet18_2,Nat),
                                                          (lizzieLet18_3,Nat),
                                                          (lizzieLet18_4,Nat)] */
  logic [3:0] readPointer_Natxadg_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_Natxadg_1_argbuf_rwb_done;
  assign lizzieLet18_1_d = {readPointer_Natxadg_1_argbuf_rwb_d[17:1],
                            (readPointer_Natxadg_1_argbuf_rwb_d[0] && (! readPointer_Natxadg_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet18_2_d = {readPointer_Natxadg_1_argbuf_rwb_d[17:1],
                            (readPointer_Natxadg_1_argbuf_rwb_d[0] && (! readPointer_Natxadg_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet18_3_d = {readPointer_Natxadg_1_argbuf_rwb_d[17:1],
                            (readPointer_Natxadg_1_argbuf_rwb_d[0] && (! readPointer_Natxadg_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet18_4_d = {readPointer_Natxadg_1_argbuf_rwb_d[17:1],
                            (readPointer_Natxadg_1_argbuf_rwb_d[0] && (! readPointer_Natxadg_1_argbuf_rwb_emitted[3]))};
  assign readPointer_Natxadg_1_argbuf_rwb_done = (readPointer_Natxadg_1_argbuf_rwb_emitted | ({lizzieLet18_4_d[0],
                                                                                               lizzieLet18_3_d[0],
                                                                                               lizzieLet18_2_d[0],
                                                                                               lizzieLet18_1_d[0]} & {lizzieLet18_4_r,
                                                                                                                      lizzieLet18_3_r,
                                                                                                                      lizzieLet18_2_r,
                                                                                                                      lizzieLet18_1_r}));
  assign readPointer_Natxadg_1_argbuf_rwb_r = (& readPointer_Natxadg_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_Natxadg_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_Natxadg_1_argbuf_rwb_emitted <= (readPointer_Natxadg_1_argbuf_rwb_r ? 4'd0 :
                                                   readPointer_Natxadg_1_argbuf_rwb_done);
  
  /* buf (Ty Nat) : (readPointer_Natyadh_1_argbuf,Nat) > (readPointer_Natyadh_1_argbuf_rwb,Nat) */
  Nat_t readPointer_Natyadh_1_argbuf_bufchan_d;
  logic readPointer_Natyadh_1_argbuf_bufchan_r;
  assign readPointer_Natyadh_1_argbuf_r = ((! readPointer_Natyadh_1_argbuf_bufchan_d[0]) || readPointer_Natyadh_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_Natyadh_1_argbuf_bufchan_d <= {17'd0, 1'd0};
    else
      if (readPointer_Natyadh_1_argbuf_r)
        readPointer_Natyadh_1_argbuf_bufchan_d <= readPointer_Natyadh_1_argbuf_d;
  Nat_t readPointer_Natyadh_1_argbuf_bufchan_buf;
  assign readPointer_Natyadh_1_argbuf_bufchan_r = (! readPointer_Natyadh_1_argbuf_bufchan_buf[0]);
  assign readPointer_Natyadh_1_argbuf_rwb_d = (readPointer_Natyadh_1_argbuf_bufchan_buf[0] ? readPointer_Natyadh_1_argbuf_bufchan_buf :
                                               readPointer_Natyadh_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_Natyadh_1_argbuf_bufchan_buf <= {17'd0, 1'd0};
    else
      if ((readPointer_Natyadh_1_argbuf_rwb_r && readPointer_Natyadh_1_argbuf_bufchan_buf[0]))
        readPointer_Natyadh_1_argbuf_bufchan_buf <= {17'd0, 1'd0};
      else if (((! readPointer_Natyadh_1_argbuf_rwb_r) && (! readPointer_Natyadh_1_argbuf_bufchan_buf[0])))
        readPointer_Natyadh_1_argbuf_bufchan_buf <= readPointer_Natyadh_1_argbuf_bufchan_d;
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolm1ad9_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolm1ad9_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolm1ad9_1_argbuf_r = ((! readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolm1ad9_1_argbuf_r)
        readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d <= readPointer_QTree_Boolm1ad9_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_r = (! readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d = (readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolm1ad9_1_argbuf_rwb_r && readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_r) && (! readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_buf <= readPointer_QTree_Boolm1ad9_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolm1ad9_1_argbuf_rwb,QTree_Bool) > [(lizzieLet2_1,QTree_Bool),
                                                                                (lizzieLet2_2,QTree_Bool),
                                                                                (lizzieLet2_3,QTree_Bool),
                                                                                (lizzieLet2_4,QTree_Bool),
                                                                                (lizzieLet2_5,QTree_Bool),
                                                                                (lizzieLet2_6,QTree_Bool),
                                                                                (lizzieLet2_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Boolm1ad9_1_argbuf_rwb_done;
  assign lizzieLet2_1_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet2_2_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet2_3_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet2_4_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet2_5_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet2_6_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet2_7_d = {readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Boolm1ad9_1_argbuf_rwb_done = (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted | ({lizzieLet2_7_d[0],
                                                                                                               lizzieLet2_6_d[0],
                                                                                                               lizzieLet2_5_d[0],
                                                                                                               lizzieLet2_4_d[0],
                                                                                                               lizzieLet2_3_d[0],
                                                                                                               lizzieLet2_2_d[0],
                                                                                                               lizzieLet2_1_d[0]} & {lizzieLet2_7_r,
                                                                                                                                     lizzieLet2_6_r,
                                                                                                                                     lizzieLet2_5_r,
                                                                                                                                     lizzieLet2_4_r,
                                                                                                                                     lizzieLet2_3_r,
                                                                                                                                     lizzieLet2_2_r,
                                                                                                                                     lizzieLet2_1_r}));
  assign readPointer_QTree_Boolm1ad9_1_argbuf_rwb_r = (& readPointer_QTree_Boolm1ad9_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Boolm1ad9_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolm1ad9_1_argbuf_rwb_r ? 7'd0 :
                                                           readPointer_QTree_Boolm1ad9_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_BoolmacS_1_argbuf,QTree_Bool) > (readPointer_QTree_BoolmacS_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_BoolmacS_1_argbuf_bufchan_d;
  logic readPointer_QTree_BoolmacS_1_argbuf_bufchan_r;
  assign readPointer_QTree_BoolmacS_1_argbuf_r = ((! readPointer_QTree_BoolmacS_1_argbuf_bufchan_d[0]) || readPointer_QTree_BoolmacS_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacS_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_BoolmacS_1_argbuf_r)
        readPointer_QTree_BoolmacS_1_argbuf_bufchan_d <= readPointer_QTree_BoolmacS_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf;
  assign readPointer_QTree_BoolmacS_1_argbuf_bufchan_r = (! readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_BoolmacS_1_argbuf_rwb_d = (readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf[0] ? readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_BoolmacS_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_BoolmacS_1_argbuf_rwb_r && readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_BoolmacS_1_argbuf_rwb_r) && (! readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_BoolmacS_1_argbuf_bufchan_buf <= readPointer_QTree_BoolmacS_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_BoolmacS_1_argbuf_rwb,QTree_Bool) > [(lizzieLet6_1,QTree_Bool),
                                                                               (lizzieLet6_2,QTree_Bool),
                                                                               (lizzieLet6_3,QTree_Bool),
                                                                               (lizzieLet6_4,QTree_Bool),
                                                                               (lizzieLet6_5,QTree_Bool),
                                                                               (lizzieLet6_6,QTree_Bool)] */
  logic [5:0] readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted;
  logic [5:0] readPointer_QTree_BoolmacS_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_BoolmacS_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_BoolmacS_1_argbuf_rwb_d[0] && (! readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted[5]))};
  assign readPointer_QTree_BoolmacS_1_argbuf_rwb_done = (readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted | ({lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_BoolmacS_1_argbuf_rwb_r = (& readPointer_QTree_BoolmacS_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted <= 6'd0;
    else
      readPointer_QTree_BoolmacS_1_argbuf_rwb_emitted <= (readPointer_QTree_BoolmacS_1_argbuf_rwb_r ? 6'd0 :
                                                          readPointer_QTree_BoolmacS_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Bool) : (readPointer_QTree_Boolmad1_1_argbuf,QTree_Bool) > (readPointer_QTree_Boolmad1_1_argbuf_rwb,QTree_Bool) */
  QTree_Bool_t readPointer_QTree_Boolmad1_1_argbuf_bufchan_d;
  logic readPointer_QTree_Boolmad1_1_argbuf_bufchan_r;
  assign readPointer_QTree_Boolmad1_1_argbuf_r = ((! readPointer_QTree_Boolmad1_1_argbuf_bufchan_d[0]) || readPointer_QTree_Boolmad1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolmad1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Boolmad1_1_argbuf_r)
        readPointer_QTree_Boolmad1_1_argbuf_bufchan_d <= readPointer_QTree_Boolmad1_1_argbuf_d;
  QTree_Bool_t readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Boolmad1_1_argbuf_bufchan_r = (! readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Boolmad1_1_argbuf_rwb_d = (readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Boolmad1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Boolmad1_1_argbuf_rwb_r && readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Boolmad1_1_argbuf_rwb_r) && (! readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Boolmad1_1_argbuf_bufchan_buf <= readPointer_QTree_Boolmad1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Bool) : (readPointer_QTree_Boolmad1_1_argbuf_rwb,QTree_Bool) > [(lizzieLet12_1_1,QTree_Bool),
                                                                               (lizzieLet12_1_2,QTree_Bool),
                                                                               (lizzieLet12_1_3,QTree_Bool),
                                                                               (lizzieLet12_1_4,QTree_Bool),
                                                                               (lizzieLet12_1_5,QTree_Bool),
                                                                               (lizzieLet12_1_6,QTree_Bool),
                                                                               (lizzieLet12_1_7,QTree_Bool)] */
  logic [6:0] readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted;
  logic [6:0] readPointer_QTree_Boolmad1_1_argbuf_rwb_done;
  assign lizzieLet12_1_1_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet12_1_2_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet12_1_3_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet12_1_4_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet12_1_5_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet12_1_6_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet12_1_7_d = {readPointer_QTree_Boolmad1_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Boolmad1_1_argbuf_rwb_d[0] && (! readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted[6]))};
  assign readPointer_QTree_Boolmad1_1_argbuf_rwb_done = (readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted | ({lizzieLet12_1_7_d[0],
                                                                                                             lizzieLet12_1_6_d[0],
                                                                                                             lizzieLet12_1_5_d[0],
                                                                                                             lizzieLet12_1_4_d[0],
                                                                                                             lizzieLet12_1_3_d[0],
                                                                                                             lizzieLet12_1_2_d[0],
                                                                                                             lizzieLet12_1_1_d[0]} & {lizzieLet12_1_7_r,
                                                                                                                                      lizzieLet12_1_6_r,
                                                                                                                                      lizzieLet12_1_5_r,
                                                                                                                                      lizzieLet12_1_4_r,
                                                                                                                                      lizzieLet12_1_3_r,
                                                                                                                                      lizzieLet12_1_2_r,
                                                                                                                                      lizzieLet12_1_1_r}));
  assign readPointer_QTree_Boolmad1_1_argbuf_rwb_r = (& readPointer_QTree_Boolmad1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted <= 7'd0;
    else
      readPointer_QTree_Boolmad1_1_argbuf_rwb_emitted <= (readPointer_QTree_Boolmad1_1_argbuf_rwb_r ? 7'd0 :
                                                          readPointer_QTree_Boolmad1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (sc_0_10_destruct,Pointer_CTmain_map'_Bool_Nat) > (sc_0_10_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTmain_map'_Bool_Nat_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (sc_0_14_destruct,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sc_0_14_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (sc_0_6_destruct,Pointer_CTkron_kron_Bool_Bool_Bool) > (sc_0_6_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (scfarg_0_1_goMux_mux,Pointer_CTmain_map'_Bool_Nat) > (scfarg_0_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTmain_map'_Bool_Nat_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (scfarg_0_2_goMux_mux,Pointer_CTmap''_map''_Bool_Bool_Bool) > (scfarg_0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (scfarg_0_goMux_mux,Pointer_CTkron_kron_Bool_Bool_Bool) > (scfarg_0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* destruct (Ty TupGo,
          Dcon TupGo) : (to_nat1TupGo_1,TupGo) > [(to_nat1TupGogo_16,Go)] */
  assign to_nat1TupGogo_16_d = to_nat1TupGo_1_d[0];
  assign to_nat1TupGo_1_r = to_nat1TupGogo_16_r;
  
  /* dcon (Ty Nat,
      Dcon Zero) : [(to_nat1TupGogo_16,Go)] > (go_16_1Zero,Nat) */
  assign go_16_1Zero_d = Zero_dc((& {to_nat1TupGogo_16_d[0]}), to_nat1TupGogo_16_d);
  assign {to_nat1TupGogo_16_r} = {1 {(go_16_1Zero_r && go_16_1Zero_d[0])}};
  
  /* buf (Ty MyBool) : (v'ad0_2_2,MyBool) > (v'ad0_2_2_argbuf,MyBool) */
  MyBool_t \v'ad0_2_2_bufchan_d ;
  logic \v'ad0_2_2_bufchan_r ;
  assign \v'ad0_2_2_r  = ((! \v'ad0_2_2_bufchan_d [0]) || \v'ad0_2_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_2_2_bufchan_d  <= {1'd0, 1'd0};
    else if (\v'ad0_2_2_r ) \v'ad0_2_2_bufchan_d  <= \v'ad0_2_2_d ;
  MyBool_t \v'ad0_2_2_bufchan_buf ;
  assign \v'ad0_2_2_bufchan_r  = (! \v'ad0_2_2_bufchan_buf [0]);
  assign \v'ad0_2_2_argbuf_d  = (\v'ad0_2_2_bufchan_buf [0] ? \v'ad0_2_2_bufchan_buf  :
                                 \v'ad0_2_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_2_2_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'ad0_2_2_argbuf_r  && \v'ad0_2_2_bufchan_buf [0]))
        \v'ad0_2_2_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'ad0_2_2_argbuf_r ) && (! \v'ad0_2_2_bufchan_buf [0])))
        \v'ad0_2_2_bufchan_buf  <= \v'ad0_2_2_bufchan_d ;
  
  /* fork (Ty MyBool) : (v'ad0_2_destruct,MyBool) > [(v'ad0_2_1,MyBool),
                                                (v'ad0_2_2,MyBool)] */
  logic [1:0] \v'ad0_2_destruct_emitted ;
  logic [1:0] \v'ad0_2_destruct_done ;
  assign \v'ad0_2_1_d  = {\v'ad0_2_destruct_d [1:1],
                          (\v'ad0_2_destruct_d [0] && (! \v'ad0_2_destruct_emitted [0]))};
  assign \v'ad0_2_2_d  = {\v'ad0_2_destruct_d [1:1],
                          (\v'ad0_2_destruct_d [0] && (! \v'ad0_2_destruct_emitted [1]))};
  assign \v'ad0_2_destruct_done  = (\v'ad0_2_destruct_emitted  | ({\v'ad0_2_2_d [0],
                                                                   \v'ad0_2_1_d [0]} & {\v'ad0_2_2_r ,
                                                                                        \v'ad0_2_1_r }));
  assign \v'ad0_2_destruct_r  = (& \v'ad0_2_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_2_destruct_emitted  <= 2'd0;
    else
      \v'ad0_2_destruct_emitted  <= (\v'ad0_2_destruct_r  ? 2'd0 :
                                     \v'ad0_2_destruct_done );
  
  /* buf (Ty MyBool) : (v'ad0_3_2,MyBool) > (v'ad0_3_2_argbuf,MyBool) */
  MyBool_t \v'ad0_3_2_bufchan_d ;
  logic \v'ad0_3_2_bufchan_r ;
  assign \v'ad0_3_2_r  = ((! \v'ad0_3_2_bufchan_d [0]) || \v'ad0_3_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_3_2_bufchan_d  <= {1'd0, 1'd0};
    else if (\v'ad0_3_2_r ) \v'ad0_3_2_bufchan_d  <= \v'ad0_3_2_d ;
  MyBool_t \v'ad0_3_2_bufchan_buf ;
  assign \v'ad0_3_2_bufchan_r  = (! \v'ad0_3_2_bufchan_buf [0]);
  assign \v'ad0_3_2_argbuf_d  = (\v'ad0_3_2_bufchan_buf [0] ? \v'ad0_3_2_bufchan_buf  :
                                 \v'ad0_3_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_3_2_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'ad0_3_2_argbuf_r  && \v'ad0_3_2_bufchan_buf [0]))
        \v'ad0_3_2_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'ad0_3_2_argbuf_r ) && (! \v'ad0_3_2_bufchan_buf [0])))
        \v'ad0_3_2_bufchan_buf  <= \v'ad0_3_2_bufchan_d ;
  
  /* fork (Ty MyBool) : (v'ad0_3_destruct,MyBool) > [(v'ad0_3_1,MyBool),
                                                (v'ad0_3_2,MyBool)] */
  logic [1:0] \v'ad0_3_destruct_emitted ;
  logic [1:0] \v'ad0_3_destruct_done ;
  assign \v'ad0_3_1_d  = {\v'ad0_3_destruct_d [1:1],
                          (\v'ad0_3_destruct_d [0] && (! \v'ad0_3_destruct_emitted [0]))};
  assign \v'ad0_3_2_d  = {\v'ad0_3_destruct_d [1:1],
                          (\v'ad0_3_destruct_d [0] && (! \v'ad0_3_destruct_emitted [1]))};
  assign \v'ad0_3_destruct_done  = (\v'ad0_3_destruct_emitted  | ({\v'ad0_3_2_d [0],
                                                                   \v'ad0_3_1_d [0]} & {\v'ad0_3_2_r ,
                                                                                        \v'ad0_3_1_r }));
  assign \v'ad0_3_destruct_r  = (& \v'ad0_3_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_3_destruct_emitted  <= 2'd0;
    else
      \v'ad0_3_destruct_emitted  <= (\v'ad0_3_destruct_r  ? 2'd0 :
                                     \v'ad0_3_destruct_done );
  
  /* buf (Ty MyBool) : (v'ad0_4_destruct,MyBool) > (v'ad0_4_1_argbuf,MyBool) */
  MyBool_t \v'ad0_4_destruct_bufchan_d ;
  logic \v'ad0_4_destruct_bufchan_r ;
  assign \v'ad0_4_destruct_r  = ((! \v'ad0_4_destruct_bufchan_d [0]) || \v'ad0_4_destruct_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'ad0_4_destruct_bufchan_d  <= {1'd0, 1'd0};
    else
      if (\v'ad0_4_destruct_r )
        \v'ad0_4_destruct_bufchan_d  <= \v'ad0_4_destruct_d ;
  MyBool_t \v'ad0_4_destruct_bufchan_buf ;
  assign \v'ad0_4_destruct_bufchan_r  = (! \v'ad0_4_destruct_bufchan_buf [0]);
  assign \v'ad0_4_1_argbuf_d  = (\v'ad0_4_destruct_bufchan_buf [0] ? \v'ad0_4_destruct_bufchan_buf  :
                                 \v'ad0_4_destruct_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \v'ad0_4_destruct_bufchan_buf  <= {1'd0, 1'd0};
    else
      if ((\v'ad0_4_1_argbuf_r  && \v'ad0_4_destruct_bufchan_buf [0]))
        \v'ad0_4_destruct_bufchan_buf  <= {1'd0, 1'd0};
      else if (((! \v'ad0_4_1_argbuf_r ) && (! \v'ad0_4_destruct_bufchan_buf [0])))
        \v'ad0_4_destruct_bufchan_buf  <= \v'ad0_4_destruct_bufchan_d ;
  
  /* buf (Ty MyBool) : (vacT_destruct,MyBool) > (vacT_1_argbuf,MyBool) */
  MyBool_t vacT_destruct_bufchan_d;
  logic vacT_destruct_bufchan_r;
  assign vacT_destruct_r = ((! vacT_destruct_bufchan_d[0]) || vacT_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacT_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (vacT_destruct_r) vacT_destruct_bufchan_d <= vacT_destruct_d;
  MyBool_t vacT_destruct_bufchan_buf;
  assign vacT_destruct_bufchan_r = (! vacT_destruct_bufchan_buf[0]);
  assign vacT_1_argbuf_d = (vacT_destruct_bufchan_buf[0] ? vacT_destruct_bufchan_buf :
                            vacT_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vacT_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((vacT_1_argbuf_r && vacT_destruct_bufchan_buf[0]))
        vacT_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! vacT_1_argbuf_r) && (! vacT_destruct_bufchan_buf[0])))
        vacT_destruct_bufchan_buf <= vacT_destruct_bufchan_d;
  
  /* buf (Ty MyBool) : (vad2_destruct,MyBool) > (vad2_1_argbuf,MyBool) */
  MyBool_t vad2_destruct_bufchan_d;
  logic vad2_destruct_bufchan_r;
  assign vad2_destruct_r = ((! vad2_destruct_bufchan_d[0]) || vad2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vad2_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (vad2_destruct_r) vad2_destruct_bufchan_d <= vad2_destruct_d;
  MyBool_t vad2_destruct_bufchan_buf;
  assign vad2_destruct_bufchan_r = (! vad2_destruct_bufchan_buf[0]);
  assign vad2_1_argbuf_d = (vad2_destruct_bufchan_buf[0] ? vad2_destruct_bufchan_buf :
                            vad2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vad2_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((vad2_1_argbuf_r && vad2_destruct_bufchan_buf[0]))
        vad2_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! vad2_1_argbuf_r) && (! vad2_destruct_bufchan_buf[0])))
        vad2_destruct_bufchan_buf <= vad2_destruct_bufchan_d;
  
  /* buf (Ty MyBool) : (vadb_destruct,MyBool) > (vadb_1_argbuf,MyBool) */
  MyBool_t vadb_destruct_bufchan_d;
  logic vadb_destruct_bufchan_r;
  assign vadb_destruct_r = ((! vadb_destruct_bufchan_d[0]) || vadb_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vadb_destruct_bufchan_d <= {1'd0, 1'd0};
    else
      if (vadb_destruct_r) vadb_destruct_bufchan_d <= vadb_destruct_d;
  MyBool_t vadb_destruct_bufchan_buf;
  assign vadb_destruct_bufchan_r = (! vadb_destruct_bufchan_buf[0]);
  assign vadb_1_argbuf_d = (vadb_destruct_bufchan_buf[0] ? vadb_destruct_bufchan_buf :
                            vadb_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vadb_destruct_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((vadb_1_argbuf_r && vadb_destruct_bufchan_buf[0]))
        vadb_destruct_bufchan_buf <= {1'd0, 1'd0};
      else if (((! vadb_1_argbuf_r) && (! vadb_destruct_bufchan_buf[0])))
        vadb_destruct_bufchan_buf <= vadb_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (lizzieLet14_1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet14_1_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf :
                                     writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((lizzieLet14_1_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! lizzieLet14_1_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca2_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca2_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet25_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca1_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca1_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet26_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d <= {16'd0,
                                                                        1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf :
                                                                      writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                          1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf <= {16'd0,
                                                                            1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca0_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                            1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                              1'd0};
    else
      if ((sca0_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                                1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) > (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf[0]);
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf :
                                                                     writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_r && writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTkron_kron_Bool_Bool_Bool) : (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb,Pointer_CTkron_kron_Bool_Bool_Bool) > (sca3_1_argbuf,Pointer_CTkron_kron_Bool_Bool_Bool) */
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  logic writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_r;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_r = ((! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d[0]) || writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                           1'd0};
    else
      if (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_r)
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d <= writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_d;
  Pointer_CTkron_kron_Bool_Bool_Bool_t writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf;
  assign writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_r = (! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0] ? writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf :
                            writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                             1'd0};
    else
      if ((sca3_1_argbuf_r && writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0]))
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                               1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf[0])))
        writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_buf <= writeCTkron_kron_Bool_Bool_BoollizzieLet4_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > (writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_r )
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_d  = (\writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_r  && \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) > (sca3_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_r )
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet10_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > (writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_r )
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_d  = (\writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_r  && \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) > (lizzieLet5_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_r )
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet5_1_1_argbuf_d = (\writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet22_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > (writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_r )
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_d  = (\writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_r  && \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) > (sca2_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_r )
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet30_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > (writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_r )
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_d  = (\writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_r  && \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) > (sca1_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_r )
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet31_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf,Pointer_CTmain_map'_Bool_Nat) > (writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d  <= {16'd0,
                                                                    1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_r )
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf [0]);
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_d  = (\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf  :
                                                                  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf  <= {16'd0,
                                                                      1'd0};
    else
      if ((\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_r  && \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf  <= {16'd0,
                                                                        1'd0};
      else if (((! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_r ) && (! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmain_map'_Bool_Nat) : (writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb,Pointer_CTmain_map'_Bool_Nat) > (sca0_1_1_argbuf,Pointer_CTmain_map'_Bool_Nat) */
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_r  = ((! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d [0]) || \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                        1'd0};
    else
      if (\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_r )
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d  <= \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_d ;
  \Pointer_CTmain_map'_Bool_Nat_t  \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_r  = (! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                          1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                            1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_buf  <= \writeCTmain_map'_Bool_NatlizzieLet32_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca3_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca3_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet16_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (lizzieLet10_1_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet10_1_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  :
                                     \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet23_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca2_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca2_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet35_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca1_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca1_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet36_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) > (writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d  <= {16'd0,
                                                                            1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf [0]);
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_d  = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf  :
                                                                          \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                              1'd0};
    else
      if ((\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_r  && \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf  <= {16'd0,
                                                                                1'd0};
      else if (((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_r ) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTmap''_map''_Bool_Bool_Bool) : (writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb,Pointer_CTmap''_map''_Bool_Bool_Bool) > (sca0_2_1_argbuf,Pointer_CTmap''_map''_Bool_Bool_Bool) */
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d ;
  logic \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_r ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_r  = ((! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d [0]) || \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                                1'd0};
    else
      if (\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_r )
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_d ;
  \Pointer_CTmap''_map''_Bool_Bool_Bool_t  \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_r  = (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_2_1_argbuf_d = (\writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0] ? \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  :
                              \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                  1'd0};
    else
      if ((sca0_2_1_argbuf_r && \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                    1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_buf  <= \writeCTmap''_map''_Bool_Bool_BoollizzieLet37_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet0_1_argbuf,Pointer_Nat) > (writeNatlizzieLet0_1_argbuf_rwb,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_bufchan_d;
  logic writeNatlizzieLet0_1_argbuf_bufchan_r;
  assign writeNatlizzieLet0_1_argbuf_r = ((! writeNatlizzieLet0_1_argbuf_bufchan_d[0]) || writeNatlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet0_1_argbuf_r)
        writeNatlizzieLet0_1_argbuf_bufchan_d <= writeNatlizzieLet0_1_argbuf_d;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_bufchan_buf;
  assign writeNatlizzieLet0_1_argbuf_bufchan_r = (! writeNatlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeNatlizzieLet0_1_argbuf_rwb_d = (writeNatlizzieLet0_1_argbuf_bufchan_buf[0] ? writeNatlizzieLet0_1_argbuf_bufchan_buf :
                                              writeNatlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeNatlizzieLet0_1_argbuf_rwb_r && writeNatlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeNatlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeNatlizzieLet0_1_argbuf_rwb_r) && (! writeNatlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeNatlizzieLet0_1_argbuf_bufchan_buf <= writeNatlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux,Pointer_Nat) > (applyfnBool_Nat_5_resbuf,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d;
  logic writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_r;
  assign writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_r = ((! writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d[0]) || writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d <= {16'd0,
                                                                          1'd0};
    else
      if (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_r)
        writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d <= writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_d;
  Pointer_Nat_t writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf;
  assign writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_r = (! writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf[0]);
  assign applyfnBool_Nat_5_resbuf_d = (writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf[0] ? writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf :
                                       writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf <= {16'd0,
                                                                            1'd0};
    else
      if ((applyfnBool_Nat_5_resbuf_r && writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf[0]))
        writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf <= {16'd0,
                                                                              1'd0};
      else if (((! applyfnBool_Nat_5_resbuf_r) && (! writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf[0])))
        writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_buf <= writeNatlizzieLet0_1_argbuf_rwbto_nat1_resbuf_mux_mux_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet1_1_argbuf,Pointer_Nat) > (writeNatlizzieLet1_1_argbuf_rwb,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_bufchan_d;
  logic writeNatlizzieLet1_1_argbuf_bufchan_r;
  assign writeNatlizzieLet1_1_argbuf_r = ((! writeNatlizzieLet1_1_argbuf_bufchan_d[0]) || writeNatlizzieLet1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet1_1_argbuf_r)
        writeNatlizzieLet1_1_argbuf_bufchan_d <= writeNatlizzieLet1_1_argbuf_d;
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_bufchan_buf;
  assign writeNatlizzieLet1_1_argbuf_bufchan_r = (! writeNatlizzieLet1_1_argbuf_bufchan_buf[0]);
  assign writeNatlizzieLet1_1_argbuf_rwb_d = (writeNatlizzieLet1_1_argbuf_bufchan_buf[0] ? writeNatlizzieLet1_1_argbuf_bufchan_buf :
                                              writeNatlizzieLet1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeNatlizzieLet1_1_argbuf_rwb_r && writeNatlizzieLet1_1_argbuf_bufchan_buf[0]))
        writeNatlizzieLet1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeNatlizzieLet1_1_argbuf_rwb_r) && (! writeNatlizzieLet1_1_argbuf_bufchan_buf[0])))
        writeNatlizzieLet1_1_argbuf_bufchan_buf <= writeNatlizzieLet1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet1_1_argbuf_rwb,Pointer_Nat) > (es_1_1_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_rwb_bufchan_d;
  logic writeNatlizzieLet1_1_argbuf_rwb_bufchan_r;
  assign writeNatlizzieLet1_1_argbuf_rwb_r = ((! writeNatlizzieLet1_1_argbuf_rwb_bufchan_d[0]) || writeNatlizzieLet1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet1_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet1_1_argbuf_rwb_r)
        writeNatlizzieLet1_1_argbuf_rwb_bufchan_d <= writeNatlizzieLet1_1_argbuf_rwb_d;
  Pointer_Nat_t writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf;
  assign writeNatlizzieLet1_1_argbuf_rwb_bufchan_r = (! writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf[0]);
  assign es_1_1_1_argbuf_d = (writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf[0] ? writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf :
                              writeNatlizzieLet1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_1_1_1_argbuf_r && writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf[0]))
        writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_1_1_1_argbuf_r) && (! writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf[0])))
        writeNatlizzieLet1_1_argbuf_rwb_bufchan_buf <= writeNatlizzieLet1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet39_1_argbuf,Pointer_Nat) > (writeNatlizzieLet39_1_argbuf_rwb,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet39_1_argbuf_bufchan_d;
  logic writeNatlizzieLet39_1_argbuf_bufchan_r;
  assign writeNatlizzieLet39_1_argbuf_r = ((! writeNatlizzieLet39_1_argbuf_bufchan_d[0]) || writeNatlizzieLet39_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet39_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet39_1_argbuf_r)
        writeNatlizzieLet39_1_argbuf_bufchan_d <= writeNatlizzieLet39_1_argbuf_d;
  Pointer_Nat_t writeNatlizzieLet39_1_argbuf_bufchan_buf;
  assign writeNatlizzieLet39_1_argbuf_bufchan_r = (! writeNatlizzieLet39_1_argbuf_bufchan_buf[0]);
  assign writeNatlizzieLet39_1_argbuf_rwb_d = (writeNatlizzieLet39_1_argbuf_bufchan_buf[0] ? writeNatlizzieLet39_1_argbuf_bufchan_buf :
                                               writeNatlizzieLet39_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeNatlizzieLet39_1_argbuf_rwb_r && writeNatlizzieLet39_1_argbuf_bufchan_buf[0]))
        writeNatlizzieLet39_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeNatlizzieLet39_1_argbuf_rwb_r) && (! writeNatlizzieLet39_1_argbuf_bufchan_buf[0])))
        writeNatlizzieLet39_1_argbuf_bufchan_buf <= writeNatlizzieLet39_1_argbuf_bufchan_d;
  
  /* dcon (Ty Nat,
      Dcon Succ) : [(writeNatlizzieLet39_1_argbuf_rwb,Pointer_Nat)] > (lizzieLet0_1_1Succ,Nat) */
  assign lizzieLet0_1_1Succ_d = Succ_dc((& {writeNatlizzieLet39_1_argbuf_rwb_d[0]}), writeNatlizzieLet39_1_argbuf_rwb_d);
  assign {writeNatlizzieLet39_1_argbuf_rwb_r} = {1 {(lizzieLet0_1_1Succ_r && lizzieLet0_1_1Succ_d[0])}};
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet40_1_argbuf,Pointer_Nat) > (writeNatlizzieLet40_1_argbuf_rwb,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_bufchan_d;
  logic writeNatlizzieLet40_1_argbuf_bufchan_r;
  assign writeNatlizzieLet40_1_argbuf_r = ((! writeNatlizzieLet40_1_argbuf_bufchan_d[0]) || writeNatlizzieLet40_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet40_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet40_1_argbuf_r)
        writeNatlizzieLet40_1_argbuf_bufchan_d <= writeNatlizzieLet40_1_argbuf_d;
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_bufchan_buf;
  assign writeNatlizzieLet40_1_argbuf_bufchan_r = (! writeNatlizzieLet40_1_argbuf_bufchan_buf[0]);
  assign writeNatlizzieLet40_1_argbuf_rwb_d = (writeNatlizzieLet40_1_argbuf_bufchan_buf[0] ? writeNatlizzieLet40_1_argbuf_bufchan_buf :
                                               writeNatlizzieLet40_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeNatlizzieLet40_1_argbuf_rwb_r && writeNatlizzieLet40_1_argbuf_bufchan_buf[0]))
        writeNatlizzieLet40_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeNatlizzieLet40_1_argbuf_rwb_r) && (! writeNatlizzieLet40_1_argbuf_bufchan_buf[0])))
        writeNatlizzieLet40_1_argbuf_bufchan_buf <= writeNatlizzieLet40_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (writeNatlizzieLet40_1_argbuf_rwb,Pointer_Nat) > (to_nat1_resbuf,Pointer_Nat) */
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_rwb_bufchan_d;
  logic writeNatlizzieLet40_1_argbuf_rwb_bufchan_r;
  assign writeNatlizzieLet40_1_argbuf_rwb_r = ((! writeNatlizzieLet40_1_argbuf_rwb_bufchan_d[0]) || writeNatlizzieLet40_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet40_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeNatlizzieLet40_1_argbuf_rwb_r)
        writeNatlizzieLet40_1_argbuf_rwb_bufchan_d <= writeNatlizzieLet40_1_argbuf_rwb_d;
  Pointer_Nat_t writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf;
  assign writeNatlizzieLet40_1_argbuf_rwb_bufchan_r = (! writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf[0]);
  assign to_nat1_resbuf_d = (writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf[0] ? writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf :
                             writeNatlizzieLet40_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((to_nat1_resbuf_r && writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf[0]))
        writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! to_nat1_resbuf_r) && (! writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf[0])))
        writeNatlizzieLet40_1_argbuf_rwb_bufchan_buf <= writeNatlizzieLet40_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_r = ((! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_1_argbuf_r)
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet13_1_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d = (writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf :
                                                        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r && writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet13_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet13_1_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet6_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                              1'd0};
    else
      if (writeQTree_BoollizzieLet13_1_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet13_1_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet6_1_1_argbuf_d = (writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                  1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet13_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_r = ((! writeQTree_BoollizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_r)
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_d = (writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet14_1_argbuf_rwb_r && writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet14_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet14_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet14_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet15_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_argbuf_r = ((! writeQTree_BoollizzieLet15_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_argbuf_r)
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet15_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_d = (writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet15_1_argbuf_rwb_r && writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet15_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet15_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet15_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet15_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet8_1_1_argbuf_d = (writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet17_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet17_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet17_1_argbuf_r = ((! writeQTree_BoollizzieLet17_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet17_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet17_1_argbuf_r)
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet17_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet17_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_d = (writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet17_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet17_1_argbuf_rwb_r && writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet17_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet17_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet17_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet17_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet17_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet17_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet17_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_r = ((! writeQTree_BoollizzieLet28_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_r)
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_d = (writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet28_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet28_1_argbuf_rwb_r && writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet28_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet28_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet28_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet28_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf :
                                 writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_1_argbuf_r && writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet28_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet38_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet38_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet38_1_argbuf_r = ((! writeQTree_BoollizzieLet38_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet38_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet38_1_argbuf_r)
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet38_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet38_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_d = (writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf :
                                                      writeQTree_BoollizzieLet38_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet38_1_argbuf_rwb_r && writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet38_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet38_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet38_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet38_1_argbuf_rwb,Pointer_QTree_Bool) > (contRet_0_2_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet38_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet38_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet38_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_r = ((! writeQTree_BoollizzieLet3_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_r)
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_d = (writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet3_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet3_1_argbuf_rwb_r && writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet3_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet3_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet11_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet3_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet3_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet3_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf,Pointer_QTree_Bool) > (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_r = ((! writeQTree_BoollizzieLet5_1_argbuf_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_r)
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_d = (writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf :
                                                     writeQTree_BoollizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_BoollizzieLet5_1_argbuf_rwb_r && writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_BoollizzieLet5_1_argbuf_rwb_r) && (! writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Bool) : (writeQTree_BoollizzieLet5_1_argbuf_rwb,Pointer_QTree_Bool) > (lizzieLet13_1_argbuf,Pointer_QTree_Bool) */
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_r = ((! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_BoollizzieLet5_1_argbuf_rwb_r)
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d <= writeQTree_BoollizzieLet5_1_argbuf_rwb_d;
  Pointer_QTree_Bool_t writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_r = (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_buf <= writeQTree_BoollizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet11_1_1_argbuf,Pointer_QTree_Nat) > (writeQTree_NatlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d;
  logic writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_r;
  assign writeQTree_NatlizzieLet11_1_1_argbuf_r = ((! writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d[0]) || writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet11_1_1_argbuf_r)
        writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d <= writeQTree_NatlizzieLet11_1_1_argbuf_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf;
  assign writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_r = (! writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_NatlizzieLet11_1_1_argbuf_rwb_d = (writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf[0] ? writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf :
                                                       writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_NatlizzieLet11_1_1_argbuf_rwb_r && writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf[0]))
        writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_NatlizzieLet11_1_1_argbuf_rwb_r) && (! writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf[0])))
        writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_buf <= writeQTree_NatlizzieLet11_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet11_1_1_argbuf_rwb,Pointer_QTree_Nat) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_NatlizzieLet11_1_1_argbuf_rwb_r = ((! writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_NatlizzieLet11_1_1_argbuf_rwb_r)
        writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d <= writeQTree_NatlizzieLet11_1_1_argbuf_rwb_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_r = (! writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_buf <= writeQTree_NatlizzieLet11_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet33_1_argbuf,Pointer_QTree_Nat) > (writeQTree_NatlizzieLet33_1_argbuf_rwb,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_bufchan_d;
  logic writeQTree_NatlizzieLet33_1_argbuf_bufchan_r;
  assign writeQTree_NatlizzieLet33_1_argbuf_r = ((! writeQTree_NatlizzieLet33_1_argbuf_bufchan_d[0]) || writeQTree_NatlizzieLet33_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet33_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet33_1_argbuf_r)
        writeQTree_NatlizzieLet33_1_argbuf_bufchan_d <= writeQTree_NatlizzieLet33_1_argbuf_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf;
  assign writeQTree_NatlizzieLet33_1_argbuf_bufchan_r = (! writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf[0]);
  assign writeQTree_NatlizzieLet33_1_argbuf_rwb_d = (writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf[0] ? writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf :
                                                     writeQTree_NatlizzieLet33_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_NatlizzieLet33_1_argbuf_rwb_r && writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf[0]))
        writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_NatlizzieLet33_1_argbuf_rwb_r) && (! writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf[0])))
        writeQTree_NatlizzieLet33_1_argbuf_bufchan_buf <= writeQTree_NatlizzieLet33_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet33_1_argbuf_rwb,Pointer_QTree_Nat) > (contRet_0_1_1_argbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d;
  logic writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_r;
  assign writeQTree_NatlizzieLet33_1_argbuf_rwb_r = ((! writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d[0]) || writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet33_1_argbuf_rwb_r)
        writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d <= writeQTree_NatlizzieLet33_1_argbuf_rwb_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_r = (! writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_buf <= writeQTree_NatlizzieLet33_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet7_1_argbuf,Pointer_QTree_Nat) > (writeQTree_NatlizzieLet7_1_argbuf_rwb,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_NatlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_NatlizzieLet7_1_argbuf_r = ((! writeQTree_NatlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_NatlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet7_1_argbuf_r)
        writeQTree_NatlizzieLet7_1_argbuf_bufchan_d <= writeQTree_NatlizzieLet7_1_argbuf_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_NatlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_NatlizzieLet7_1_argbuf_rwb_d = (writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_NatlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_NatlizzieLet7_1_argbuf_rwb_r && writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_NatlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_NatlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_NatlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet7_1_argbuf_rwb,Pointer_QTree_Nat) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_NatlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet7_1_argbuf_rwb_r)
        writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_NatlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_NatlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet8_1_argbuf,Pointer_QTree_Nat) > (writeQTree_NatlizzieLet8_1_argbuf_rwb,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_bufchan_d;
  logic writeQTree_NatlizzieLet8_1_argbuf_bufchan_r;
  assign writeQTree_NatlizzieLet8_1_argbuf_r = ((! writeQTree_NatlizzieLet8_1_argbuf_bufchan_d[0]) || writeQTree_NatlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet8_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet8_1_argbuf_r)
        writeQTree_NatlizzieLet8_1_argbuf_bufchan_d <= writeQTree_NatlizzieLet8_1_argbuf_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf;
  assign writeQTree_NatlizzieLet8_1_argbuf_bufchan_r = (! writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeQTree_NatlizzieLet8_1_argbuf_rwb_d = (writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf[0] ? writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf :
                                                    writeQTree_NatlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_NatlizzieLet8_1_argbuf_rwb_r && writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_NatlizzieLet8_1_argbuf_rwb_r) && (! writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeQTree_NatlizzieLet8_1_argbuf_bufchan_buf <= writeQTree_NatlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet8_1_argbuf_rwb,Pointer_QTree_Nat) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeQTree_NatlizzieLet8_1_argbuf_rwb_r = ((! writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet8_1_argbuf_rwb_r)
        writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d <= writeQTree_NatlizzieLet8_1_argbuf_rwb_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeQTree_NatlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet9_1_argbuf,Pointer_QTree_Nat) > (writeQTree_NatlizzieLet9_1_argbuf_rwb,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_NatlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_NatlizzieLet9_1_argbuf_r = ((! writeQTree_NatlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_NatlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet9_1_argbuf_r)
        writeQTree_NatlizzieLet9_1_argbuf_bufchan_d <= writeQTree_NatlizzieLet9_1_argbuf_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_NatlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_NatlizzieLet9_1_argbuf_rwb_d = (writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_NatlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_NatlizzieLet9_1_argbuf_rwb_r && writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_NatlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_NatlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_NatlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Nat) : (writeQTree_NatlizzieLet9_1_argbuf_rwb,Pointer_QTree_Nat) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Nat) */
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_NatlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_NatlizzieLet9_1_argbuf_rwb_r)
        writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_NatlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Nat_t writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_NatlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (xacw_1,Pointer_Nat) > (xacw_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t xacw_1_bufchan_d;
  logic xacw_1_bufchan_r;
  assign xacw_1_r = ((! xacw_1_bufchan_d[0]) || xacw_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacw_1_bufchan_d <= {16'd0, 1'd0};
    else if (xacw_1_r) xacw_1_bufchan_d <= xacw_1_d;
  Pointer_Nat_t xacw_1_bufchan_buf;
  assign xacw_1_bufchan_r = (! xacw_1_bufchan_buf[0]);
  assign xacw_1_argbuf_d = (xacw_1_bufchan_buf[0] ? xacw_1_bufchan_buf :
                            xacw_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacw_1_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((xacw_1_argbuf_r && xacw_1_bufchan_buf[0]))
        xacw_1_bufchan_buf <= {16'd0, 1'd0};
      else if (((! xacw_1_argbuf_r) && (! xacw_1_bufchan_buf[0])))
        xacw_1_bufchan_buf <= xacw_1_bufchan_d;
  
  /* buf (Ty MyBool) : (xacw_1_1,MyBool) > (xacw_1_1_argbuf,MyBool) */
  MyBool_t xacw_1_1_bufchan_d;
  logic xacw_1_1_bufchan_r;
  assign xacw_1_1_r = ((! xacw_1_1_bufchan_d[0]) || xacw_1_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacw_1_1_bufchan_d <= {1'd0, 1'd0};
    else if (xacw_1_1_r) xacw_1_1_bufchan_d <= xacw_1_1_d;
  MyBool_t xacw_1_1_bufchan_buf;
  assign xacw_1_1_bufchan_r = (! xacw_1_1_bufchan_buf[0]);
  assign xacw_1_1_argbuf_d = (xacw_1_1_bufchan_buf[0] ? xacw_1_1_bufchan_buf :
                              xacw_1_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xacw_1_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((xacw_1_1_argbuf_r && xacw_1_1_bufchan_buf[0]))
        xacw_1_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! xacw_1_1_argbuf_r) && (! xacw_1_1_bufchan_buf[0])))
        xacw_1_1_bufchan_buf <= xacw_1_1_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (xadg_goMux_mux,Pointer_Nat) > (xadg_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t xadg_goMux_mux_bufchan_d;
  logic xadg_goMux_mux_bufchan_r;
  assign xadg_goMux_mux_r = ((! xadg_goMux_mux_bufchan_d[0]) || xadg_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xadg_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (xadg_goMux_mux_r) xadg_goMux_mux_bufchan_d <= xadg_goMux_mux_d;
  Pointer_Nat_t xadg_goMux_mux_bufchan_buf;
  assign xadg_goMux_mux_bufchan_r = (! xadg_goMux_mux_bufchan_buf[0]);
  assign xadg_1_argbuf_d = (xadg_goMux_mux_bufchan_buf[0] ? xadg_goMux_mux_bufchan_buf :
                            xadg_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) xadg_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((xadg_1_argbuf_r && xadg_goMux_mux_bufchan_buf[0]))
        xadg_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! xadg_1_argbuf_r) && (! xadg_goMux_mux_bufchan_buf[0])))
        xadg_goMux_mux_bufchan_buf <= xadg_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (y1adk_destruct,Pointer_Nat) > (y1adk_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t y1adk_destruct_bufchan_d;
  logic y1adk_destruct_bufchan_r;
  assign y1adk_destruct_r = ((! y1adk_destruct_bufchan_d[0]) || y1adk_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) y1adk_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (y1adk_destruct_r) y1adk_destruct_bufchan_d <= y1adk_destruct_d;
  Pointer_Nat_t y1adk_destruct_bufchan_buf;
  assign y1adk_destruct_bufchan_r = (! y1adk_destruct_bufchan_buf[0]);
  assign y1adk_1_argbuf_d = (y1adk_destruct_bufchan_buf[0] ? y1adk_destruct_bufchan_buf :
                             y1adk_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) y1adk_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((y1adk_1_argbuf_r && y1adk_destruct_bufchan_buf[0]))
        y1adk_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! y1adk_1_argbuf_r) && (! y1adk_destruct_bufchan_buf[0])))
        y1adk_destruct_bufchan_buf <= y1adk_destruct_bufchan_d;
  
  /* buf (Ty Pointer_Nat) : (yadh_goMux_mux,Pointer_Nat) > (yadh_1_argbuf,Pointer_Nat) */
  Pointer_Nat_t yadh_goMux_mux_bufchan_d;
  logic yadh_goMux_mux_bufchan_r;
  assign yadh_goMux_mux_r = ((! yadh_goMux_mux_bufchan_d[0]) || yadh_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) yadh_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (yadh_goMux_mux_r) yadh_goMux_mux_bufchan_d <= yadh_goMux_mux_d;
  Pointer_Nat_t yadh_goMux_mux_bufchan_buf;
  assign yadh_goMux_mux_bufchan_r = (! yadh_goMux_mux_bufchan_buf[0]);
  assign yadh_1_argbuf_d = (yadh_goMux_mux_bufchan_buf[0] ? yadh_goMux_mux_bufchan_buf :
                            yadh_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) yadh_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((yadh_1_argbuf_r && yadh_goMux_mux_bufchan_buf[0]))
        yadh_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! yadh_1_argbuf_r) && (! yadh_goMux_mux_bufchan_buf[0])))
        yadh_goMux_mux_bufchan_buf <= yadh_goMux_mux_bufchan_d;
endmodule