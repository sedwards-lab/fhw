`timescale 1ns/1ns
package mMaskAdd_package ;
    typedef logic [4:0] \Int4#_t ;
    typedef logic [8:0] \Int8#_t ;
    typedef logic [16:0] \Int16#_t ;
    typedef logic [32:0] \Int#_t ;
    typedef logic [4:0] \Word4#_t ;
    typedef logic [8:0] \Word8#_t ;
    typedef logic [16:0] \Word16#_t ;
    typedef logic [32:0] \Word#_t ;
    typedef logic [5:0] C30_t;
    function C30_t C1_30_dc (logic valid);
      begin
        C1_30_dc = 6'bx;
        C1_30_dc[0:0] = valid;
        C1_30_dc[5:1] = 5'd0;
      end
    endfunction
    function C30_t C2_30_dc (logic valid);
      begin
        C2_30_dc = 6'bx;
        C2_30_dc[0:0] = valid;
        C2_30_dc[5:1] = 5'd1;
      end
    endfunction
    function C30_t C3_30_dc (logic valid);
      begin
        C3_30_dc = 6'bx;
        C3_30_dc[0:0] = valid;
        C3_30_dc[5:1] = 5'd2;
      end
    endfunction
    function C30_t C4_30_dc (logic valid);
      begin
        C4_30_dc = 6'bx;
        C4_30_dc[0:0] = valid;
        C4_30_dc[5:1] = 5'd3;
      end
    endfunction
    function C30_t C5_30_dc (logic valid);
      begin
        C5_30_dc = 6'bx;
        C5_30_dc[0:0] = valid;
        C5_30_dc[5:1] = 5'd4;
      end
    endfunction
    function C30_t C6_30_dc (logic valid);
      begin
        C6_30_dc = 6'bx;
        C6_30_dc[0:0] = valid;
        C6_30_dc[5:1] = 5'd5;
      end
    endfunction
    function C30_t C7_30_dc (logic valid);
      begin
        C7_30_dc = 6'bx;
        C7_30_dc[0:0] = valid;
        C7_30_dc[5:1] = 5'd6;
      end
    endfunction
    function C30_t C8_30_dc (logic valid);
      begin
        C8_30_dc = 6'bx;
        C8_30_dc[0:0] = valid;
        C8_30_dc[5:1] = 5'd7;
      end
    endfunction
    function C30_t C9_30_dc (logic valid);
      begin
        C9_30_dc = 6'bx;
        C9_30_dc[0:0] = valid;
        C9_30_dc[5:1] = 5'd8;
      end
    endfunction
    function C30_t C10_30_dc (logic valid);
      begin
        C10_30_dc = 6'bx;
        C10_30_dc[0:0] = valid;
        C10_30_dc[5:1] = 5'd9;
      end
    endfunction
    function C30_t C11_30_dc (logic valid);
      begin
        C11_30_dc = 6'bx;
        C11_30_dc[0:0] = valid;
        C11_30_dc[5:1] = 5'd10;
      end
    endfunction
    function C30_t C12_30_dc (logic valid);
      begin
        C12_30_dc = 6'bx;
        C12_30_dc[0:0] = valid;
        C12_30_dc[5:1] = 5'd11;
      end
    endfunction
    function C30_t C13_30_dc (logic valid);
      begin
        C13_30_dc = 6'bx;
        C13_30_dc[0:0] = valid;
        C13_30_dc[5:1] = 5'd12;
      end
    endfunction
    function C30_t C14_30_dc (logic valid);
      begin
        C14_30_dc = 6'bx;
        C14_30_dc[0:0] = valid;
        C14_30_dc[5:1] = 5'd13;
      end
    endfunction
    function C30_t C15_30_dc (logic valid);
      begin
        C15_30_dc = 6'bx;
        C15_30_dc[0:0] = valid;
        C15_30_dc[5:1] = 5'd14;
      end
    endfunction
    function C30_t C16_30_dc (logic valid);
      begin
        C16_30_dc = 6'bx;
        C16_30_dc[0:0] = valid;
        C16_30_dc[5:1] = 5'd15;
      end
    endfunction
    function C30_t C17_30_dc (logic valid);
      begin
        C17_30_dc = 6'bx;
        C17_30_dc[0:0] = valid;
        C17_30_dc[5:1] = 5'd16;
      end
    endfunction
    function C30_t C18_30_dc (logic valid);
      begin
        C18_30_dc = 6'bx;
        C18_30_dc[0:0] = valid;
        C18_30_dc[5:1] = 5'd17;
      end
    endfunction
    function C30_t C19_30_dc (logic valid);
      begin
        C19_30_dc = 6'bx;
        C19_30_dc[0:0] = valid;
        C19_30_dc[5:1] = 5'd18;
      end
    endfunction
    function C30_t C20_30_dc (logic valid);
      begin
        C20_30_dc = 6'bx;
        C20_30_dc[0:0] = valid;
        C20_30_dc[5:1] = 5'd19;
      end
    endfunction
    function C30_t C21_30_dc (logic valid);
      begin
        C21_30_dc = 6'bx;
        C21_30_dc[0:0] = valid;
        C21_30_dc[5:1] = 5'd20;
      end
    endfunction
    function C30_t C22_30_dc (logic valid);
      begin
        C22_30_dc = 6'bx;
        C22_30_dc[0:0] = valid;
        C22_30_dc[5:1] = 5'd21;
      end
    endfunction
    function C30_t C23_30_dc (logic valid);
      begin
        C23_30_dc = 6'bx;
        C23_30_dc[0:0] = valid;
        C23_30_dc[5:1] = 5'd22;
      end
    endfunction
    function C30_t C24_30_dc (logic valid);
      begin
        C24_30_dc = 6'bx;
        C24_30_dc[0:0] = valid;
        C24_30_dc[5:1] = 5'd23;
      end
    endfunction
    function C30_t C25_30_dc (logic valid);
      begin
        C25_30_dc = 6'bx;
        C25_30_dc[0:0] = valid;
        C25_30_dc[5:1] = 5'd24;
      end
    endfunction
    function C30_t C26_30_dc (logic valid);
      begin
        C26_30_dc = 6'bx;
        C26_30_dc[0:0] = valid;
        C26_30_dc[5:1] = 5'd25;
      end
    endfunction
    function C30_t C27_30_dc (logic valid);
      begin
        C27_30_dc = 6'bx;
        C27_30_dc[0:0] = valid;
        C27_30_dc[5:1] = 5'd26;
      end
    endfunction
    function C30_t C28_30_dc (logic valid);
      begin
        C28_30_dc = 6'bx;
        C28_30_dc[0:0] = valid;
        C28_30_dc[5:1] = 5'd27;
      end
    endfunction
    function C30_t C29_30_dc (logic valid);
      begin
        C29_30_dc = 6'bx;
        C29_30_dc[0:0] = valid;
        C29_30_dc[5:1] = 5'd28;
      end
    endfunction
    function C30_t C30_30_dc (logic valid);
      begin
        C30_30_dc = 6'bx;
        C30_30_dc[0:0] = valid;
        C30_30_dc[5:1] = 5'd29;
      end
    endfunction
    typedef logic [0:0] Go_t;
    function Go_t Go_dc (logic valid);
      begin
        Go_dc = 1'bx;
        Go_dc[0:0] = valid;
      end
    endfunction
    typedef logic [16:0] Pointer_QTree_Bool_t;
    function Pointer_QTree_Bool_t Pointer_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_QTree_Bool_dc = 17'bx;
        Pointer_QTree_Bool_dc[0:0] = valid;
        Pointer_QTree_Bool_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [1:0] MyBool_t;
    function MyBool_t MyFalse_dc (logic valid, Go_t z1);
      begin
        MyFalse_dc = 2'bx;
        MyFalse_dc[0:0] = valid;
        MyFalse_dc[1:1] = 1'd0;
        ;
      end
    endfunction
    function MyBool_t MyTrue_dc (logic valid, Go_t z1);
      begin
        MyTrue_dc = 2'bx;
        MyTrue_dc[0:0] = valid;
        MyTrue_dc[1:1] = 1'd1;
        ;
      end
    endfunction
    typedef logic [66:0] QTree_Bool_t;
    function QTree_Bool_t QNone_Bool_dc (logic valid, Go_t z1);
      begin
        QNone_Bool_dc = 67'bx;
        QNone_Bool_dc[0:0] = valid;
        QNone_Bool_dc[2:1] = 2'd0;
        ;
      end
    endfunction
    function QTree_Bool_t QVal_Bool_dc (logic valid, MyBool_t z1);
      begin
        QVal_Bool_dc = 67'bx;
        QVal_Bool_dc[0:0] = valid;
        QVal_Bool_dc[2:1] = 2'd1;
        QVal_Bool_dc[3:3] = z1[1:1];
      end
    endfunction
    function QTree_Bool_t QNode_Bool_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        QNode_Bool_dc = 67'bx;
        QNode_Bool_dc[0:0] = valid;
        QNode_Bool_dc[2:1] = 2'd2;
        QNode_Bool_dc[18:3] = z1[16:1];
        QNode_Bool_dc[34:19] = z2[16:1];
        QNode_Bool_dc[50:35] = z3[16:1];
        QNode_Bool_dc[66:51] = z4[16:1];
      end
    endfunction
    function QTree_Bool_t QError_Bool_dc (logic valid, Go_t z1);
      begin
        QError_Bool_dc = 67'bx;
        QError_Bool_dc[0:0] = valid;
        QError_Bool_dc[2:1] = 2'd3;
        ;
      end
    endfunction
    typedef logic [83:0] MemIn_QTree_Bool_t;
    function MemIn_QTree_Bool_t ReadIn_QTree_Bool_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_QTree_Bool_dc = 84'bx;
        ReadIn_QTree_Bool_dc[0:0] = valid;
        ReadIn_QTree_Bool_dc[1:1] = 1'd0;
        ReadIn_QTree_Bool_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_QTree_Bool_t WriteIn_QTree_Bool_dc (logic valid, \Word16#_t  z1, QTree_Bool_t z2);
      begin
        WriteIn_QTree_Bool_dc = 84'bx;
        WriteIn_QTree_Bool_dc[0:0] = valid;
        WriteIn_QTree_Bool_dc[1:1] = 1'd1;
        WriteIn_QTree_Bool_dc[17:2] = z1[16:1];
        WriteIn_QTree_Bool_dc[83:18] = z2[66:1];
      end
    endfunction
    typedef logic [67:0] MemOut_QTree_Bool_t;
    function MemOut_QTree_Bool_t ReadOut_QTree_Bool_dc (logic valid, QTree_Bool_t z1);
      begin
        ReadOut_QTree_Bool_dc = 68'bx;
        ReadOut_QTree_Bool_dc[0:0] = valid;
        ReadOut_QTree_Bool_dc[1:1] = 1'd0;
        ReadOut_QTree_Bool_dc[67:2] = z1[66:1];
      end
    endfunction
    function MemOut_QTree_Bool_t ACK_QTree_Bool_dc (logic valid);
      begin
        ACK_QTree_Bool_dc = 68'bx;
        ACK_QTree_Bool_dc[0:0] = valid;
        ACK_QTree_Bool_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] Pointer_CTf_t;
    function Pointer_CTf_t Pointer_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_CTf_dc = 17'bx;
        Pointer_CTf_dc[0:0] = valid;
        Pointer_CTf_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [16:0] Pointer_MaskQTree_t;
    function Pointer_MaskQTree_t Pointer_MaskQTree_dc (logic valid, \Word16#_t  z1);
      begin
        Pointer_MaskQTree_dc = 17'bx;
        Pointer_MaskQTree_dc[0:0] = valid;
        Pointer_MaskQTree_dc[16:1] = z1[16:1];
      end
    endfunction
    typedef logic [163:0] CTf_t;
    function CTf_t Lfsbos_dc (logic valid, Go_t z1);
      begin
        Lfsbos_dc = 164'bx;
        Lfsbos_dc[0:0] = valid;
        Lfsbos_dc[3:1] = 3'd0;
        ;
      end
    endfunction
    function CTf_t Lcall_f3_dc (logic valid, Pointer_CTf_t z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_MaskQTree_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7, Pointer_MaskQTree_t z8, Pointer_QTree_Bool_t z9, Pointer_QTree_Bool_t z10);
      begin
        Lcall_f3_dc = 164'bx;
        Lcall_f3_dc[0:0] = valid;
        Lcall_f3_dc[3:1] = 3'd1;
        Lcall_f3_dc[19:4] = z1[16:1];
        Lcall_f3_dc[35:20] = z2[16:1];
        Lcall_f3_dc[51:36] = z3[16:1];
        Lcall_f3_dc[67:52] = z4[16:1];
        Lcall_f3_dc[83:68] = z5[16:1];
        Lcall_f3_dc[99:84] = z6[16:1];
        Lcall_f3_dc[115:100] = z7[16:1];
        Lcall_f3_dc[131:116] = z8[16:1];
        Lcall_f3_dc[147:132] = z9[16:1];
        Lcall_f3_dc[163:148] = z10[16:1];
      end
    endfunction
    function CTf_t Lcall_f2_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_CTf_t z2, Pointer_MaskQTree_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_MaskQTree_t z6, Pointer_QTree_Bool_t z7, Pointer_QTree_Bool_t z8);
      begin
        Lcall_f2_dc = 164'bx;
        Lcall_f2_dc[0:0] = valid;
        Lcall_f2_dc[3:1] = 3'd2;
        Lcall_f2_dc[19:4] = z1[16:1];
        Lcall_f2_dc[35:20] = z2[16:1];
        Lcall_f2_dc[51:36] = z3[16:1];
        Lcall_f2_dc[67:52] = z4[16:1];
        Lcall_f2_dc[83:68] = z5[16:1];
        Lcall_f2_dc[99:84] = z6[16:1];
        Lcall_f2_dc[115:100] = z7[16:1];
        Lcall_f2_dc[131:116] = z8[16:1];
      end
    endfunction
    function CTf_t Lcall_f1_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_CTf_t z3, Pointer_MaskQTree_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6);
      begin
        Lcall_f1_dc = 164'bx;
        Lcall_f1_dc[0:0] = valid;
        Lcall_f1_dc[3:1] = 3'd3;
        Lcall_f1_dc[19:4] = z1[16:1];
        Lcall_f1_dc[35:20] = z2[16:1];
        Lcall_f1_dc[51:36] = z3[16:1];
        Lcall_f1_dc[67:52] = z4[16:1];
        Lcall_f1_dc[83:68] = z5[16:1];
        Lcall_f1_dc[99:84] = z6[16:1];
      end
    endfunction
    function CTf_t Lcall_f0_dc (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_CTf_t z4);
      begin
        Lcall_f0_dc = 164'bx;
        Lcall_f0_dc[0:0] = valid;
        Lcall_f0_dc[3:1] = 3'd4;
        Lcall_f0_dc[19:4] = z1[16:1];
        Lcall_f0_dc[35:20] = z2[16:1];
        Lcall_f0_dc[51:36] = z3[16:1];
        Lcall_f0_dc[67:52] = z4[16:1];
      end
    endfunction
    typedef logic [180:0] MemIn_CTf_t;
    function MemIn_CTf_t ReadIn_CTf_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_CTf_dc = 181'bx;
        ReadIn_CTf_dc[0:0] = valid;
        ReadIn_CTf_dc[1:1] = 1'd0;
        ReadIn_CTf_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_CTf_t WriteIn_CTf_dc (logic valid, \Word16#_t  z1, CTf_t z2);
      begin
        WriteIn_CTf_dc = 181'bx;
        WriteIn_CTf_dc[0:0] = valid;
        WriteIn_CTf_dc[1:1] = 1'd1;
        WriteIn_CTf_dc[17:2] = z1[16:1];
        WriteIn_CTf_dc[180:18] = z2[163:1];
      end
    endfunction
    typedef logic [164:0] MemOut_CTf_t;
    function MemOut_CTf_t ReadOut_CTf_dc (logic valid, CTf_t z1);
      begin
        ReadOut_CTf_dc = 165'bx;
        ReadOut_CTf_dc[0:0] = valid;
        ReadOut_CTf_dc[1:1] = 1'd0;
        ReadOut_CTf_dc[164:2] = z1[163:1];
      end
    endfunction
    function MemOut_CTf_t ACK_CTf_dc (logic valid);
      begin
        ACK_CTf_dc = 165'bx;
        ACK_CTf_dc[0:0] = valid;
        ACK_CTf_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] \Pointer_CTf'_t ;
    function \Pointer_CTf'_t  \Pointer_CTf'_dc  (logic valid, \Word16#_t  z1);
      begin
        \Pointer_CTf'_dc  = 17'bx;
        \Pointer_CTf'_dc [0:0] = valid;
        \Pointer_CTf'_dc [16:1] = z1[16:1];
      end
    endfunction
    typedef logic [115:0] \CTf'_t ;
    function \CTf'_t  \Lf'sbos_dc  (logic valid, Go_t z1);
      begin
        \Lf'sbos_dc  = 116'bx;
        \Lf'sbos_dc [0:0] = valid;
        \Lf'sbos_dc [3:1] = 3'd0;
        ;
      end
    endfunction
    function \CTf'_t  \Lcall_f'3_dc  (logic valid, \Pointer_CTf'_t  z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6, Pointer_QTree_Bool_t z7);
      begin
        \Lcall_f'3_dc  = 116'bx;
        \Lcall_f'3_dc [0:0] = valid;
        \Lcall_f'3_dc [3:1] = 3'd1;
        \Lcall_f'3_dc [19:4] = z1[16:1];
        \Lcall_f'3_dc [35:20] = z2[16:1];
        \Lcall_f'3_dc [51:36] = z3[16:1];
        \Lcall_f'3_dc [67:52] = z4[16:1];
        \Lcall_f'3_dc [83:68] = z5[16:1];
        \Lcall_f'3_dc [99:84] = z6[16:1];
        \Lcall_f'3_dc [115:100] = z7[16:1];
      end
    endfunction
    function \CTf'_t  \Lcall_f'2_dc  (logic valid, Pointer_QTree_Bool_t z1, \Pointer_CTf'_t  z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5, Pointer_QTree_Bool_t z6);
      begin
        \Lcall_f'2_dc  = 116'bx;
        \Lcall_f'2_dc [0:0] = valid;
        \Lcall_f'2_dc [3:1] = 3'd2;
        \Lcall_f'2_dc [19:4] = z1[16:1];
        \Lcall_f'2_dc [35:20] = z2[16:1];
        \Lcall_f'2_dc [51:36] = z3[16:1];
        \Lcall_f'2_dc [67:52] = z4[16:1];
        \Lcall_f'2_dc [83:68] = z5[16:1];
        \Lcall_f'2_dc [99:84] = z6[16:1];
      end
    endfunction
    function \CTf'_t  \Lcall_f'1_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, \Pointer_CTf'_t  z3, Pointer_QTree_Bool_t z4, Pointer_QTree_Bool_t z5);
      begin
        \Lcall_f'1_dc  = 116'bx;
        \Lcall_f'1_dc [0:0] = valid;
        \Lcall_f'1_dc [3:1] = 3'd3;
        \Lcall_f'1_dc [19:4] = z1[16:1];
        \Lcall_f'1_dc [35:20] = z2[16:1];
        \Lcall_f'1_dc [51:36] = z3[16:1];
        \Lcall_f'1_dc [67:52] = z4[16:1];
        \Lcall_f'1_dc [83:68] = z5[16:1];
      end
    endfunction
    function \CTf'_t  \Lcall_f'0_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf'_t  z4);
      begin
        \Lcall_f'0_dc  = 116'bx;
        \Lcall_f'0_dc [0:0] = valid;
        \Lcall_f'0_dc [3:1] = 3'd4;
        \Lcall_f'0_dc [19:4] = z1[16:1];
        \Lcall_f'0_dc [35:20] = z2[16:1];
        \Lcall_f'0_dc [51:36] = z3[16:1];
        \Lcall_f'0_dc [67:52] = z4[16:1];
      end
    endfunction
    typedef logic [132:0] \MemIn_CTf'_t ;
    function \MemIn_CTf'_t  \ReadIn_CTf'_dc  (logic valid, \Word16#_t  z1);
      begin
        \ReadIn_CTf'_dc  = 133'bx;
        \ReadIn_CTf'_dc [0:0] = valid;
        \ReadIn_CTf'_dc [1:1] = 1'd0;
        \ReadIn_CTf'_dc [17:2] = z1[16:1];
      end
    endfunction
    function \MemIn_CTf'_t  \WriteIn_CTf'_dc  (logic valid, \Word16#_t  z1, \CTf'_t  z2);
      begin
        \WriteIn_CTf'_dc  = 133'bx;
        \WriteIn_CTf'_dc [0:0] = valid;
        \WriteIn_CTf'_dc [1:1] = 1'd1;
        \WriteIn_CTf'_dc [17:2] = z1[16:1];
        \WriteIn_CTf'_dc [132:18] = z2[115:1];
      end
    endfunction
    typedef logic [116:0] \MemOut_CTf'_t ;
    function \MemOut_CTf'_t  \ReadOut_CTf'_dc  (logic valid, \CTf'_t  z1);
      begin
        \ReadOut_CTf'_dc  = 117'bx;
        \ReadOut_CTf'_dc [0:0] = valid;
        \ReadOut_CTf'_dc [1:1] = 1'd0;
        \ReadOut_CTf'_dc [116:2] = z1[115:1];
      end
    endfunction
    function \MemOut_CTf'_t  \ACK_CTf'_dc  (logic valid);
      begin
        \ACK_CTf'_dc  = 117'bx;
        \ACK_CTf'_dc [0:0] = valid;
        \ACK_CTf'_dc [1:1] = 1'd1;
      end
    endfunction
    typedef logic [16:0] \Pointer_CTf'''''''''_f'''''''''_Bool_t ;
    function \Pointer_CTf'''''''''_f'''''''''_Bool_t  \Pointer_CTf'''''''''_f'''''''''_Bool_dc  (logic valid, \Word16#_t  z1);
      begin
        \Pointer_CTf'''''''''_f'''''''''_Bool_dc  = 17'bx;
        \Pointer_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        \Pointer_CTf'''''''''_f'''''''''_Bool_dc [16:1] = z1[16:1];
      end
    endfunction
    typedef logic [115:0] \CTf'''''''''_f'''''''''_Bool_t ;
    function \CTf'''''''''_f'''''''''_Bool_t  \Lf'''''''''_f'''''''''_Boolsbos_dc  (logic valid, Go_t z1);
      begin
        \Lf'''''''''_f'''''''''_Boolsbos_dc  = 116'bx;
        \Lf'''''''''_f'''''''''_Boolsbos_dc [0:0] = valid;
        \Lf'''''''''_f'''''''''_Boolsbos_dc [3:1] = 3'd0;
        ;
      end
    endfunction
    function \CTf'''''''''_f'''''''''_Bool_t  \Lcall_f'''''''''_f'''''''''_Bool3_dc  (logic valid, \Pointer_CTf'''''''''_f'''''''''_Bool_t  z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3, Pointer_MaskQTree_t z4, Pointer_QTree_Bool_t z5, Pointer_MaskQTree_t z6, Pointer_QTree_Bool_t z7);
      begin
        \Lcall_f'''''''''_f'''''''''_Bool3_dc  = 116'bx;
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [0:0] = valid;
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [3:1] = 3'd1;
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [19:4] = z1[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [35:20] = z2[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [51:36] = z3[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [67:52] = z4[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [83:68] = z5[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [99:84] = z6[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool3_dc [115:100] = z7[16:1];
      end
    endfunction
    function \CTf'''''''''_f'''''''''_Bool_t  \Lcall_f'''''''''_f'''''''''_Bool2_dc  (logic valid, Pointer_QTree_Bool_t z1, \Pointer_CTf'''''''''_f'''''''''_Bool_t  z2, Pointer_MaskQTree_t z3, Pointer_QTree_Bool_t z4, Pointer_MaskQTree_t z5, Pointer_QTree_Bool_t z6);
      begin
        \Lcall_f'''''''''_f'''''''''_Bool2_dc  = 116'bx;
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [0:0] = valid;
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [3:1] = 3'd2;
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [19:4] = z1[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [35:20] = z2[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [51:36] = z3[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [67:52] = z4[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [83:68] = z5[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool2_dc [99:84] = z6[16:1];
      end
    endfunction
    function \CTf'''''''''_f'''''''''_Bool_t  \Lcall_f'''''''''_f'''''''''_Bool1_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, \Pointer_CTf'''''''''_f'''''''''_Bool_t  z3, Pointer_MaskQTree_t z4, Pointer_QTree_Bool_t z5);
      begin
        \Lcall_f'''''''''_f'''''''''_Bool1_dc  = 116'bx;
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [0:0] = valid;
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [3:1] = 3'd3;
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [19:4] = z1[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [35:20] = z2[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [51:36] = z3[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [67:52] = z4[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool1_dc [83:68] = z5[16:1];
      end
    endfunction
    function \CTf'''''''''_f'''''''''_Bool_t  \Lcall_f'''''''''_f'''''''''_Bool0_dc  (logic valid, Pointer_QTree_Bool_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf'''''''''_f'''''''''_Bool_t  z4);
      begin
        \Lcall_f'''''''''_f'''''''''_Bool0_dc  = 116'bx;
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [0:0] = valid;
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [3:1] = 3'd4;
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [19:4] = z1[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [35:20] = z2[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [51:36] = z3[16:1];
        \Lcall_f'''''''''_f'''''''''_Bool0_dc [67:52] = z4[16:1];
      end
    endfunction
    typedef logic [132:0] \MemIn_CTf'''''''''_f'''''''''_Bool_t ;
    function \MemIn_CTf'''''''''_f'''''''''_Bool_t  \ReadIn_CTf'''''''''_f'''''''''_Bool_dc  (logic valid, \Word16#_t  z1);
      begin
        \ReadIn_CTf'''''''''_f'''''''''_Bool_dc  = 133'bx;
        \ReadIn_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        \ReadIn_CTf'''''''''_f'''''''''_Bool_dc [1:1] = 1'd0;
        \ReadIn_CTf'''''''''_f'''''''''_Bool_dc [17:2] = z1[16:1];
      end
    endfunction
    function \MemIn_CTf'''''''''_f'''''''''_Bool_t  \WriteIn_CTf'''''''''_f'''''''''_Bool_dc  (logic valid, \Word16#_t  z1, \CTf'''''''''_f'''''''''_Bool_t  z2);
      begin
        \WriteIn_CTf'''''''''_f'''''''''_Bool_dc  = 133'bx;
        \WriteIn_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        \WriteIn_CTf'''''''''_f'''''''''_Bool_dc [1:1] = 1'd1;
        \WriteIn_CTf'''''''''_f'''''''''_Bool_dc [17:2] = z1[16:1];
        \WriteIn_CTf'''''''''_f'''''''''_Bool_dc [132:18] = z2[115:1];
      end
    endfunction
    typedef logic [116:0] \MemOut_CTf'''''''''_f'''''''''_Bool_t ;
    function \MemOut_CTf'''''''''_f'''''''''_Bool_t  \ReadOut_CTf'''''''''_f'''''''''_Bool_dc  (logic valid, \CTf'''''''''_f'''''''''_Bool_t  z1);
      begin
        \ReadOut_CTf'''''''''_f'''''''''_Bool_dc  = 117'bx;
        \ReadOut_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        \ReadOut_CTf'''''''''_f'''''''''_Bool_dc [1:1] = 1'd0;
        \ReadOut_CTf'''''''''_f'''''''''_Bool_dc [116:2] = z1[115:1];
      end
    endfunction
    function \MemOut_CTf'''''''''_f'''''''''_Bool_t  \ACK_CTf'''''''''_f'''''''''_Bool_dc  (logic valid);
      begin
        \ACK_CTf'''''''''_f'''''''''_Bool_dc  = 117'bx;
        \ACK_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        \ACK_CTf'''''''''_f'''''''''_Bool_dc [1:1] = 1'd1;
      end
    endfunction
    typedef logic [66:0] MaskQTree_t;
    function MaskQTree_t MQNone_dc (logic valid, Go_t z1);
      begin
        MQNone_dc = 67'bx;
        MQNone_dc[0:0] = valid;
        MQNone_dc[2:1] = 2'd0;
        ;
      end
    endfunction
    function MaskQTree_t MQVal_dc (logic valid, Go_t z1);
      begin
        MQVal_dc = 67'bx;
        MQVal_dc[0:0] = valid;
        MQVal_dc[2:1] = 2'd1;
        ;
      end
    endfunction
    function MaskQTree_t MQNode_dc (logic valid, Pointer_MaskQTree_t z1, Pointer_MaskQTree_t z2, Pointer_MaskQTree_t z3, Pointer_MaskQTree_t z4);
      begin
        MQNode_dc = 67'bx;
        MQNode_dc[0:0] = valid;
        MQNode_dc[2:1] = 2'd2;
        MQNode_dc[18:3] = z1[16:1];
        MQNode_dc[34:19] = z2[16:1];
        MQNode_dc[50:35] = z3[16:1];
        MQNode_dc[66:51] = z4[16:1];
      end
    endfunction
    typedef logic [83:0] MemIn_MaskQTree_t;
    function MemIn_MaskQTree_t ReadIn_MaskQTree_dc (logic valid, \Word16#_t  z1);
      begin
        ReadIn_MaskQTree_dc = 84'bx;
        ReadIn_MaskQTree_dc[0:0] = valid;
        ReadIn_MaskQTree_dc[1:1] = 1'd0;
        ReadIn_MaskQTree_dc[17:2] = z1[16:1];
      end
    endfunction
    function MemIn_MaskQTree_t WriteIn_MaskQTree_dc (logic valid, \Word16#_t  z1, MaskQTree_t z2);
      begin
        WriteIn_MaskQTree_dc = 84'bx;
        WriteIn_MaskQTree_dc[0:0] = valid;
        WriteIn_MaskQTree_dc[1:1] = 1'd1;
        WriteIn_MaskQTree_dc[17:2] = z1[16:1];
        WriteIn_MaskQTree_dc[83:18] = z2[66:1];
      end
    endfunction
    typedef logic [67:0] MemOut_MaskQTree_t;
    function MemOut_MaskQTree_t ReadOut_MaskQTree_dc (logic valid, MaskQTree_t z1);
      begin
        ReadOut_MaskQTree_dc = 68'bx;
        ReadOut_MaskQTree_dc[0:0] = valid;
        ReadOut_MaskQTree_dc[1:1] = 1'd0;
        ReadOut_MaskQTree_dc[67:2] = z1[66:1];
      end
    endfunction
    function MemOut_MaskQTree_t ACK_MaskQTree_dc (logic valid);
      begin
        ACK_MaskQTree_dc = 68'bx;
        ACK_MaskQTree_dc[0:0] = valid;
        ACK_MaskQTree_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [3:0] C8_t;
    function C8_t C1_8_dc (logic valid);
      begin
        C1_8_dc = 4'bx;
        C1_8_dc[0:0] = valid;
        C1_8_dc[3:1] = 3'd0;
      end
    endfunction
    function C8_t C2_8_dc (logic valid);
      begin
        C2_8_dc = 4'bx;
        C2_8_dc[0:0] = valid;
        C2_8_dc[3:1] = 3'd1;
      end
    endfunction
    function C8_t C3_8_dc (logic valid);
      begin
        C3_8_dc = 4'bx;
        C3_8_dc[0:0] = valid;
        C3_8_dc[3:1] = 3'd2;
      end
    endfunction
    function C8_t C4_8_dc (logic valid);
      begin
        C4_8_dc = 4'bx;
        C4_8_dc[0:0] = valid;
        C4_8_dc[3:1] = 3'd3;
      end
    endfunction
    function C8_t C5_8_dc (logic valid);
      begin
        C5_8_dc = 4'bx;
        C5_8_dc[0:0] = valid;
        C5_8_dc[3:1] = 3'd4;
      end
    endfunction
    function C8_t C6_8_dc (logic valid);
      begin
        C6_8_dc = 4'bx;
        C6_8_dc[0:0] = valid;
        C6_8_dc[3:1] = 3'd5;
      end
    endfunction
    function C8_t C7_8_dc (logic valid);
      begin
        C7_8_dc = 4'bx;
        C7_8_dc[0:0] = valid;
        C7_8_dc[3:1] = 3'd6;
      end
    endfunction
    function C8_t C8_8_dc (logic valid);
      begin
        C8_8_dc = 4'bx;
        C8_8_dc[0:0] = valid;
        C8_8_dc[3:1] = 3'd7;
      end
    endfunction
    typedef logic [4:0] C12_t;
    function C12_t C1_12_dc (logic valid);
      begin
        C1_12_dc = 5'bx;
        C1_12_dc[0:0] = valid;
        C1_12_dc[4:1] = 4'd0;
      end
    endfunction
    function C12_t C2_12_dc (logic valid);
      begin
        C2_12_dc = 5'bx;
        C2_12_dc[0:0] = valid;
        C2_12_dc[4:1] = 4'd1;
      end
    endfunction
    function C12_t C3_12_dc (logic valid);
      begin
        C3_12_dc = 5'bx;
        C3_12_dc[0:0] = valid;
        C3_12_dc[4:1] = 4'd2;
      end
    endfunction
    function C12_t C4_12_dc (logic valid);
      begin
        C4_12_dc = 5'bx;
        C4_12_dc[0:0] = valid;
        C4_12_dc[4:1] = 4'd3;
      end
    endfunction
    function C12_t C5_12_dc (logic valid);
      begin
        C5_12_dc = 5'bx;
        C5_12_dc[0:0] = valid;
        C5_12_dc[4:1] = 4'd4;
      end
    endfunction
    function C12_t C6_12_dc (logic valid);
      begin
        C6_12_dc = 5'bx;
        C6_12_dc[0:0] = valid;
        C6_12_dc[4:1] = 4'd5;
      end
    endfunction
    function C12_t C7_12_dc (logic valid);
      begin
        C7_12_dc = 5'bx;
        C7_12_dc[0:0] = valid;
        C7_12_dc[4:1] = 4'd6;
      end
    endfunction
    function C12_t C8_12_dc (logic valid);
      begin
        C8_12_dc = 5'bx;
        C8_12_dc[0:0] = valid;
        C8_12_dc[4:1] = 4'd7;
      end
    endfunction
    function C12_t C9_12_dc (logic valid);
      begin
        C9_12_dc = 5'bx;
        C9_12_dc[0:0] = valid;
        C9_12_dc[4:1] = 4'd8;
      end
    endfunction
    function C12_t C10_12_dc (logic valid);
      begin
        C10_12_dc = 5'bx;
        C10_12_dc[0:0] = valid;
        C10_12_dc[4:1] = 4'd9;
      end
    endfunction
    function C12_t C11_12_dc (logic valid);
      begin
        C11_12_dc = 5'bx;
        C11_12_dc[0:0] = valid;
        C11_12_dc[4:1] = 4'd10;
      end
    endfunction
    function C12_t C12_12_dc (logic valid);
      begin
        C12_12_dc = 5'bx;
        C12_12_dc[0:0] = valid;
        C12_12_dc[4:1] = 4'd11;
      end
    endfunction
    typedef logic [3:0] C6_t;
    function C6_t C1_6_dc (logic valid);
      begin
        C1_6_dc = 4'bx;
        C1_6_dc[0:0] = valid;
        C1_6_dc[3:1] = 3'd0;
      end
    endfunction
    function C6_t C2_6_dc (logic valid);
      begin
        C2_6_dc = 4'bx;
        C2_6_dc[0:0] = valid;
        C2_6_dc[3:1] = 3'd1;
      end
    endfunction
    function C6_t C3_6_dc (logic valid);
      begin
        C3_6_dc = 4'bx;
        C3_6_dc[0:0] = valid;
        C3_6_dc[3:1] = 3'd2;
      end
    endfunction
    function C6_t C4_6_dc (logic valid);
      begin
        C4_6_dc = 4'bx;
        C4_6_dc[0:0] = valid;
        C4_6_dc[3:1] = 3'd3;
      end
    endfunction
    function C6_t C5_6_dc (logic valid);
      begin
        C5_6_dc = 4'bx;
        C5_6_dc[0:0] = valid;
        C5_6_dc[3:1] = 3'd4;
      end
    endfunction
    function C6_t C6_6_dc (logic valid);
      begin
        C6_6_dc = 4'bx;
        C6_6_dc[0:0] = valid;
        C6_6_dc[3:1] = 3'd5;
      end
    endfunction
    typedef logic [3:0] C5_t;
    function C5_t C1_5_dc (logic valid);
      begin
        C1_5_dc = 4'bx;
        C1_5_dc[0:0] = valid;
        C1_5_dc[3:1] = 3'd0;
      end
    endfunction
    function C5_t C2_5_dc (logic valid);
      begin
        C2_5_dc = 4'bx;
        C2_5_dc[0:0] = valid;
        C2_5_dc[3:1] = 3'd1;
      end
    endfunction
    function C5_t C3_5_dc (logic valid);
      begin
        C3_5_dc = 4'bx;
        C3_5_dc[0:0] = valid;
        C3_5_dc[3:1] = 3'd2;
      end
    endfunction
    function C5_t C4_5_dc (logic valid);
      begin
        C4_5_dc = 4'bx;
        C4_5_dc[0:0] = valid;
        C4_5_dc[3:1] = 3'd3;
      end
    endfunction
    function C5_t C5_5_dc (logic valid);
      begin
        C5_5_dc = 4'bx;
        C5_5_dc[0:0] = valid;
        C5_5_dc[3:1] = 3'd4;
      end
    endfunction
    typedef logic [5:0] C17_t;
    function C17_t C1_17_dc (logic valid);
      begin
        C1_17_dc = 6'bx;
        C1_17_dc[0:0] = valid;
        C1_17_dc[5:1] = 5'd0;
      end
    endfunction
    function C17_t C2_17_dc (logic valid);
      begin
        C2_17_dc = 6'bx;
        C2_17_dc[0:0] = valid;
        C2_17_dc[5:1] = 5'd1;
      end
    endfunction
    function C17_t C3_17_dc (logic valid);
      begin
        C3_17_dc = 6'bx;
        C3_17_dc[0:0] = valid;
        C3_17_dc[5:1] = 5'd2;
      end
    endfunction
    function C17_t C4_17_dc (logic valid);
      begin
        C4_17_dc = 6'bx;
        C4_17_dc[0:0] = valid;
        C4_17_dc[5:1] = 5'd3;
      end
    endfunction
    function C17_t C5_17_dc (logic valid);
      begin
        C5_17_dc = 6'bx;
        C5_17_dc[0:0] = valid;
        C5_17_dc[5:1] = 5'd4;
      end
    endfunction
    function C17_t C6_17_dc (logic valid);
      begin
        C6_17_dc = 6'bx;
        C6_17_dc[0:0] = valid;
        C6_17_dc[5:1] = 5'd5;
      end
    endfunction
    function C17_t C7_17_dc (logic valid);
      begin
        C7_17_dc = 6'bx;
        C7_17_dc[0:0] = valid;
        C7_17_dc[5:1] = 5'd6;
      end
    endfunction
    function C17_t C8_17_dc (logic valid);
      begin
        C8_17_dc = 6'bx;
        C8_17_dc[0:0] = valid;
        C8_17_dc[5:1] = 5'd7;
      end
    endfunction
    function C17_t C9_17_dc (logic valid);
      begin
        C9_17_dc = 6'bx;
        C9_17_dc[0:0] = valid;
        C9_17_dc[5:1] = 5'd8;
      end
    endfunction
    function C17_t C10_17_dc (logic valid);
      begin
        C10_17_dc = 6'bx;
        C10_17_dc[0:0] = valid;
        C10_17_dc[5:1] = 5'd9;
      end
    endfunction
    function C17_t C11_17_dc (logic valid);
      begin
        C11_17_dc = 6'bx;
        C11_17_dc[0:0] = valid;
        C11_17_dc[5:1] = 5'd10;
      end
    endfunction
    function C17_t C12_17_dc (logic valid);
      begin
        C12_17_dc = 6'bx;
        C12_17_dc[0:0] = valid;
        C12_17_dc[5:1] = 5'd11;
      end
    endfunction
    function C17_t C13_17_dc (logic valid);
      begin
        C13_17_dc = 6'bx;
        C13_17_dc[0:0] = valid;
        C13_17_dc[5:1] = 5'd12;
      end
    endfunction
    function C17_t C14_17_dc (logic valid);
      begin
        C14_17_dc = 6'bx;
        C14_17_dc[0:0] = valid;
        C14_17_dc[5:1] = 5'd13;
      end
    endfunction
    function C17_t C15_17_dc (logic valid);
      begin
        C15_17_dc = 6'bx;
        C15_17_dc[0:0] = valid;
        C15_17_dc[5:1] = 5'd14;
      end
    endfunction
    function C17_t C16_17_dc (logic valid);
      begin
        C16_17_dc = 6'bx;
        C16_17_dc[0:0] = valid;
        C16_17_dc[5:1] = 5'd15;
      end
    endfunction
    function C17_t C17_17_dc (logic valid);
      begin
        C17_17_dc = 6'bx;
        C17_17_dc[0:0] = valid;
        C17_17_dc[5:1] = 5'd16;
      end
    endfunction
    typedef logic [1:0] C2_t;
    function C2_t C1_2_dc (logic valid);
      begin
        C1_2_dc = 2'bx;
        C1_2_dc[0:0] = valid;
        C1_2_dc[1:1] = 1'd0;
      end
    endfunction
    function C2_t C2_2_dc (logic valid);
      begin
        C2_2_dc = 2'bx;
        C2_2_dc[0:0] = valid;
        C2_2_dc[1:1] = 1'd1;
      end
    endfunction
    typedef logic [48:0] \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_t ;
    function \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_t  \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc  (logic valid, Go_t z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf'''''''''_f'''''''''_Bool_t  z4);
      begin
        \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc  = 49'bx;
        \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc [0:0] = valid;
        ;
        \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc [16:1] = z2[16:1];
        \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc [32:17] = z3[16:1];
        \TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_CTf'''''''''_f'''''''''_Bool_dc [48:33] = z4[16:1];
      end
    endfunction
    typedef logic [48:0] \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_t ;
    function \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_t  \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc  (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3, \Pointer_CTf'_t  z4);
      begin
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc  = 49'bx;
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc [0:0] = valid;
        ;
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc [16:1] = z2[16:1];
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc [32:17] = z3[16:1];
        \TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf'_dc [48:33] = z4[16:1];
      end
    endfunction
    typedef logic [64:0] TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t;
    function TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_t TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc (logic valid, Go_t z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4, Pointer_CTf_t z5);
      begin
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc = 65'bx;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[0:0] = valid;
        ;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[16:1] = z2[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[32:17] = z3[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[48:33] = z4[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool___Pointer_CTf_dc[64:49] = z5[16:1];
      end
    endfunction
    typedef logic [32:0] TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t;
    function TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_t TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3);
      begin
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc = 33'bx;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
      end
    endfunction
    typedef logic [32:0] TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t;
    function TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_t TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_QTree_Bool_t z2, Pointer_QTree_Bool_t z3);
      begin
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc = 33'bx;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
      end
    endfunction
    typedef logic [48:0] TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_t;
    function TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_t TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc (logic valid, Go_t z1, Pointer_MaskQTree_t z2, Pointer_QTree_Bool_t z3, Pointer_QTree_Bool_t z4);
      begin
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc = 49'bx;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[0:0] = valid;
        ;
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[16:1] = z2[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[32:17] = z3[16:1];
        TupGo___Pointer_MaskQTree___Pointer_QTree_Bool___Pointer_QTree_Bool_dc[48:33] = z4[16:1];
      end
    endfunction
    typedef logic [0:0] TupGo_t;
    function TupGo_t TupGo_dc (logic valid, Go_t z1);
      begin
        TupGo_dc = 1'bx;
        TupGo_dc[0:0] = valid;
        ;
      end
    endfunction
endpackage