`timescale 1ns/1ns
import mMapKron_package::*;

module mMapKron(
  input logic clk,
  input logic reset,
  input Go_t \\QTree_Int_src_d ,
  output logic \\QTree_Int_src_r ,
  input QTree_Int_t dummy_write_QTree_Int_d,
  output logic dummy_write_QTree_Int_r,
  input Go_t sourceGo_d,
  output logic sourceGo_r,
  input Pointer_QTree_Int_t m1ahS_0_d,
  output logic m1ahS_0_r,
  input Pointer_QTree_Int_t m2ahT_1_d,
  output logic m2ahT_1_r,
  output \Word16#_t  forkHP1_QTree_Int_snk_dout,
  input logic forkHP1_QTree_Int_snk_rout,
  output Pointer_QTree_Int_t dummy_write_QTree_Int_sink_dout,
  input logic dummy_write_QTree_Int_sink_rout,
  output Int_t \es_7_1I#_dout ,
  input logic \es_7_1I#_rout 
  );
  /* --define=INPUTS=((__05CQTree_Int_src, 0, 1, Go), (dummy_write_QTree_Int, 66, 73786976294838206464, QTree_Int), (sourceGo, 0, 1, Go), (m1ahS_0, 16, 65536, Pointer_QTree_Int), (m2ahT_1, 16, 65536, Pointer_QTree_Int)) */
  /* --define=TAPS=() */
  /* --define=OUTPUTS=((forkHP1_QTree_Int_snk, 16, 65536, Word16__023), (dummy_write_QTree_Int_sink, 16, 65536, Pointer_QTree_Int), (es_7_1I__023, 32, 4294967296, Int)) */
  /* TYPE_START
CT__024wnnz_Int 16 3 (0,[0]) (1,[16p,16p,16p,16p]) (2,[32,16p,16p,16p]) (3,[32,32,16p,16p]) (4,[32,32,32,16p])
QTree_Int 16 2 (0,[0]) (1,[32]) (2,[16p,16p,16p,16p]) (3,[0])
CTf__027_f__027_Int_Int_Int_Int 16 3 (0,[0]) (1,[16p,16p,0,0,32,0,0,16p,16p]) (2,[16p,16p,16p,0,0,32,0,0,16p]) (3,[16p,16p,16p,16p,0,0,32,0,0]) (4,[16p,16p,16p,16p])
CTf_f_Int_Int_Int_Int 16 3 (0,[0]) (1,[16p,16p,16p,0,0,0,0,16p,16p]) (2,[16p,16p,16p,16p,0,0,0,0,16p]) (3,[16p,16p,16p,16p,16p,0,0,0,0]) (4,[16p,16p,16p,16p])
TupGo___Pointer_QTree_Int 16 0 (0,[0,16p])
TupGo___Pointer_QTree_Int___Pointer_CT__024wnnz_Int 16 0 (0,[0,16p,16p])
TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf__027_f__027_Int_Int_Int_Int 16 0 (0,[0,16p,0,0,32,0,0,16p])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int 16 0 (0,[0,16p,16p,0,0,0,0,16p])
TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int 16 0 (0,[0,16p,0,0,32,0,0])
TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int 16 0 (0,[0,16p,16p,0,0,0,0])
TYPE_END */
  /*  */
  /*  */
  Go_t go_1_d;
  logic go_1_r;
  Go_t go_2_d;
  logic go_2_r;
  Go_t go_3_d;
  logic go_3_r;
  Go_t go_4_d;
  logic go_4_r;
  Go_t go_5_d;
  logic go_5_r;
  Go_t go_6_d;
  logic go_6_r;
  Go_t go__7_d;
  logic go__7_r;
  Go_t go__8_d;
  logic go__8_r;
  Go_t go__9_d;
  logic go__9_r;
  Go_t go__10_d;
  logic go__10_r;
  Go_t go__11_d;
  logic go__11_r;
  Go_t go__12_d;
  logic go__12_r;
  \Word16#_t  initHP_CT$wnnz_Int_d;
  logic initHP_CT$wnnz_Int_r;
  \Word16#_t  incrHP_CT$wnnz_Int_d;
  logic incrHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_d;
  logic incrHP_mergeCT$wnnz_Int_r;
  Go_t incrHP_CT$wnnz_Int1_d;
  logic incrHP_CT$wnnz_Int1_r;
  Go_t incrHP_CT$wnnz_Int2_d;
  logic incrHP_CT$wnnz_Int2_r;
  \Word16#_t  addHP_CT$wnnz_Int_d;
  logic addHP_CT$wnnz_Int_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_d;
  logic mergeHP_CT$wnnz_Int_r;
  Go_t incrHP_mergeCT$wnnz_Int_buf_d;
  logic incrHP_mergeCT$wnnz_Int_buf_r;
  \Word16#_t  mergeHP_CT$wnnz_Int_buf_d;
  logic mergeHP_CT$wnnz_Int_buf_r;
  \Word16#_t  forkHP1_CT$wnnz_Int_d;
  logic forkHP1_CT$wnnz_Int_r;
  \Word16#_t  forkHP1_CT$wnnz_In2_d;
  logic forkHP1_CT$wnnz_In2_r;
  \Word16#_t  forkHP1_CT$wnnz_In3_d;
  logic forkHP1_CT$wnnz_In3_r;
  C2_t memMergeChoice_CT$wnnz_Int_d;
  logic memMergeChoice_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_d;
  logic memMergeIn_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_d;
  logic memOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memReadOut_CT$wnnz_Int_d;
  logic memReadOut_CT$wnnz_Int_r;
  MemOut_CT$wnnz_Int_t memWriteOut_CT$wnnz_Int_d;
  logic memWriteOut_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_dbuf_d;
  logic memMergeIn_CT$wnnz_Int_dbuf_r;
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_rbuf_d;
  logic memMergeIn_CT$wnnz_Int_rbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_dbuf_d;
  logic memOut_CT$wnnz_Int_dbuf_r;
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_rbuf_d;
  logic memOut_CT$wnnz_Int_rbuf_r;
  \Word16#_t  destructReadIn_CT$wnnz_Int_d;
  logic destructReadIn_CT$wnnz_Int_r;
  MemIn_CT$wnnz_Int_t dconReadIn_CT$wnnz_Int_d;
  logic dconReadIn_CT$wnnz_Int_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  C5_t writeMerge_choice_CT$wnnz_Int_d;
  logic writeMerge_choice_CT$wnnz_Int_r;
  CT$wnnz_Int_t writeMerge_data_CT$wnnz_Int_d;
  logic writeMerge_data_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet20_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet21_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet22_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_r;
  MemIn_CT$wnnz_Int_t dconWriteIn_CT$wnnz_Int_d;
  logic dconWriteIn_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t dconPtr_CT$wnnz_Int_d;
  logic dconPtr_CT$wnnz_Int_r;
  Pointer_CT$wnnz_Int_t _45_d;
  logic _45_r;
  assign _45_r = 1'd1;
  Pointer_CT$wnnz_Int_t demuxWriteResult_CT$wnnz_Int_d;
  logic demuxWriteResult_CT$wnnz_Int_r;
  \Word16#_t  initHP_QTree_Int_d;
  logic initHP_QTree_Int_r;
  \Word16#_t  incrHP_QTree_Int_d;
  logic incrHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_d;
  logic incrHP_mergeQTree_Int_r;
  Go_t incrHP_QTree_Int1_d;
  logic incrHP_QTree_Int1_r;
  Go_t incrHP_QTree_Int2_d;
  logic incrHP_QTree_Int2_r;
  \Word16#_t  addHP_QTree_Int_d;
  logic addHP_QTree_Int_r;
  \Word16#_t  mergeHP_QTree_Int_d;
  logic mergeHP_QTree_Int_r;
  Go_t incrHP_mergeQTree_Int_buf_d;
  logic incrHP_mergeQTree_Int_buf_r;
  \Word16#_t  mergeHP_QTree_Int_buf_d;
  logic mergeHP_QTree_Int_buf_r;
  Go_t go_1_dummy_write_QTree_Int_d;
  logic go_1_dummy_write_QTree_Int_r;
  Go_t go_2_dummy_write_QTree_Int_d;
  logic go_2_dummy_write_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_d;
  logic forkHP1_QTree_Int_r;
  \Word16#_t  forkHP1_QTree_Int_snk_d;
  logic forkHP1_QTree_Int_snk_r;
  \Word16#_t  forkHP1_QTree_In3_d;
  logic forkHP1_QTree_In3_r;
  \Word16#_t  forkHP1_QTree_In4_d;
  logic forkHP1_QTree_In4_r;
  C2_t memMergeChoice_QTree_Int_d;
  logic memMergeChoice_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_d;
  logic memMergeIn_QTree_Int_r;
  MemOut_QTree_Int_t memOut_QTree_Int_d;
  logic memOut_QTree_Int_r;
  MemOut_QTree_Int_t memReadOut_QTree_Int_d;
  logic memReadOut_QTree_Int_r;
  MemOut_QTree_Int_t memWriteOut_QTree_Int_d;
  logic memWriteOut_QTree_Int_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_dbuf_d;
  logic memMergeIn_QTree_Int_dbuf_r;
  MemIn_QTree_Int_t memMergeIn_QTree_Int_rbuf_d;
  logic memMergeIn_QTree_Int_rbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_dbuf_d;
  logic memOut_QTree_Int_dbuf_r;
  MemOut_QTree_Int_t memOut_QTree_Int_rbuf_d;
  logic memOut_QTree_Int_rbuf_r;
  C3_t readMerge_choice_QTree_Int_d;
  logic readMerge_choice_QTree_Int_r;
  Pointer_QTree_Int_t readMerge_data_QTree_Int_d;
  logic readMerge_data_QTree_Int_r;
  QTree_Int_t readPointer_QTree_Intm1ahU_1_argbuf_d;
  logic readPointer_QTree_Intm1ahU_1_argbuf_r;
  QTree_Int_t readPointer_QTree_Intm2ai5_1_argbuf_d;
  logic readPointer_QTree_Intm2ai5_1_argbuf_r;
  QTree_Int_t readPointer_QTree_IntwstH_1_1_argbuf_d;
  logic readPointer_QTree_IntwstH_1_1_argbuf_r;
  \Word16#_t  destructReadIn_QTree_Int_d;
  logic destructReadIn_QTree_Int_r;
  MemIn_QTree_Int_t dconReadIn_QTree_Int_d;
  logic dconReadIn_QTree_Int_r;
  QTree_Int_t destructReadOut_QTree_Int_d;
  logic destructReadOut_QTree_Int_r;
  C10_t writeMerge_choice_QTree_Int_d;
  logic writeMerge_choice_QTree_Int_r;
  QTree_Int_t writeMerge_data_QTree_Int_d;
  logic writeMerge_data_QTree_Int_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_r;
  Pointer_QTree_Int_t dummy_write_QTree_Int_sink_d;
  logic dummy_write_QTree_Int_sink_r;
  MemIn_QTree_Int_t dconWriteIn_QTree_Int_d;
  logic dconWriteIn_QTree_Int_r;
  Pointer_QTree_Int_t dconPtr_QTree_Int_d;
  logic dconPtr_QTree_Int_r;
  Pointer_QTree_Int_t _44_d;
  logic _44_r;
  assign _44_r = 1'd1;
  Pointer_QTree_Int_t demuxWriteResult_QTree_Int_d;
  logic demuxWriteResult_QTree_Int_r;
  \Word16#_t  \initHP_CTf'_f'_Int_Int_Int_Int_d ;
  logic \initHP_CTf'_f'_Int_Int_Int_Int_r ;
  \Word16#_t  \incrHP_CTf'_f'_Int_Int_Int_Int_d ;
  logic \incrHP_CTf'_f'_Int_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTf'_f'_Int_Int_Int_Int_d ;
  logic \incrHP_mergeCTf'_f'_Int_Int_Int_Int_r ;
  Go_t \incrHP_CTf'_f'_Int_Int_Int_Int1_d ;
  logic \incrHP_CTf'_f'_Int_Int_Int_Int1_r ;
  Go_t \incrHP_CTf'_f'_Int_Int_Int_Int2_d ;
  logic \incrHP_CTf'_f'_Int_Int_Int_Int2_r ;
  \Word16#_t  \addHP_CTf'_f'_Int_Int_Int_Int_d ;
  logic \addHP_CTf'_f'_Int_Int_Int_Int_r ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_Int_Int_Int_d ;
  logic \mergeHP_CTf'_f'_Int_Int_Int_Int_r ;
  Go_t \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_d ;
  logic \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_r ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d ;
  logic \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_r ;
  \Word16#_t  \forkHP1_CTf'_f'_Int_Int_Int_Int_d ;
  logic \forkHP1_CTf'_f'_Int_Int_Int_Int_r ;
  \Word16#_t  \forkHP1_CTf'_f'_Int_Int_Int_In2_d ;
  logic \forkHP1_CTf'_f'_Int_Int_Int_In2_r ;
  \Word16#_t  \forkHP1_CTf'_f'_Int_Int_Int_In3_d ;
  logic \forkHP1_CTf'_f'_Int_Int_Int_In3_r ;
  C2_t \memMergeChoice_CTf'_f'_Int_Int_Int_Int_d ;
  logic \memMergeChoice_CTf'_f'_Int_Int_Int_Int_r ;
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \memMergeIn_CTf'_f'_Int_Int_Int_Int_d ;
  logic \memMergeIn_CTf'_f'_Int_Int_Int_Int_r ;
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memOut_CTf'_f'_Int_Int_Int_Int_d ;
  logic \memOut_CTf'_f'_Int_Int_Int_Int_r ;
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memReadOut_CTf'_f'_Int_Int_Int_Int_d ;
  logic \memReadOut_CTf'_f'_Int_Int_Int_Int_r ;
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memWriteOut_CTf'_f'_Int_Int_Int_Int_d ;
  logic \memWriteOut_CTf'_f'_Int_Int_Int_Int_r ;
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d ;
  logic \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_r ;
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_d ;
  logic \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_r ;
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d ;
  logic \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_r ;
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_d ;
  logic \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_r ;
  \Word16#_t  \destructReadIn_CTf'_f'_Int_Int_Int_Int_d ;
  logic \destructReadIn_CTf'_f'_Int_Int_Int_Int_r ;
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \dconReadIn_CTf'_f'_Int_Int_Int_Int_d ;
  logic \dconReadIn_CTf'_f'_Int_Int_Int_Int_r ;
  \CTf'_f'_Int_Int_Int_Int_t  \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_d ;
  logic \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_r ;
  C5_t \writeMerge_choice_CTf'_f'_Int_Int_Int_Int_d ;
  logic \writeMerge_choice_CTf'_f'_Int_Int_Int_Int_r ;
  \CTf'_f'_Int_Int_Int_Int_t  \writeMerge_data_CTf'_f'_Int_Int_Int_Int_d ;
  logic \writeMerge_data_CTf'_f'_Int_Int_Int_Int_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_r ;
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \dconWriteIn_CTf'_f'_Int_Int_Int_Int_d ;
  logic \dconWriteIn_CTf'_f'_Int_Int_Int_Int_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \dconPtr_CTf'_f'_Int_Int_Int_Int_d ;
  logic \dconPtr_CTf'_f'_Int_Int_Int_Int_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  _43_d;
  logic _43_r;
  assign _43_r = 1'd1;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d ;
  logic \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_r ;
  \Word16#_t  initHP_CTf_f_Int_Int_Int_Int_d;
  logic initHP_CTf_f_Int_Int_Int_Int_r;
  \Word16#_t  incrHP_CTf_f_Int_Int_Int_Int_d;
  logic incrHP_CTf_f_Int_Int_Int_Int_r;
  Go_t incrHP_mergeCTf_f_Int_Int_Int_Int_d;
  logic incrHP_mergeCTf_f_Int_Int_Int_Int_r;
  Go_t incrHP_CTf_f_Int_Int_Int_Int1_d;
  logic incrHP_CTf_f_Int_Int_Int_Int1_r;
  Go_t incrHP_CTf_f_Int_Int_Int_Int2_d;
  logic incrHP_CTf_f_Int_Int_Int_Int2_r;
  \Word16#_t  addHP_CTf_f_Int_Int_Int_Int_d;
  logic addHP_CTf_f_Int_Int_Int_Int_r;
  \Word16#_t  mergeHP_CTf_f_Int_Int_Int_Int_d;
  logic mergeHP_CTf_f_Int_Int_Int_Int_r;
  Go_t incrHP_mergeCTf_f_Int_Int_Int_Int_buf_d;
  logic incrHP_mergeCTf_f_Int_Int_Int_Int_buf_r;
  \Word16#_t  mergeHP_CTf_f_Int_Int_Int_Int_buf_d;
  logic mergeHP_CTf_f_Int_Int_Int_Int_buf_r;
  \Word16#_t  forkHP1_CTf_f_Int_Int_Int_Int_d;
  logic forkHP1_CTf_f_Int_Int_Int_Int_r;
  \Word16#_t  forkHP1_CTf_f_Int_Int_Int_In2_d;
  logic forkHP1_CTf_f_Int_Int_Int_In2_r;
  \Word16#_t  forkHP1_CTf_f_Int_Int_Int_In3_d;
  logic forkHP1_CTf_f_Int_Int_Int_In3_r;
  C2_t memMergeChoice_CTf_f_Int_Int_Int_Int_d;
  logic memMergeChoice_CTf_f_Int_Int_Int_Int_r;
  MemIn_CTf_f_Int_Int_Int_Int_t memMergeIn_CTf_f_Int_Int_Int_Int_d;
  logic memMergeIn_CTf_f_Int_Int_Int_Int_r;
  MemOut_CTf_f_Int_Int_Int_Int_t memOut_CTf_f_Int_Int_Int_Int_d;
  logic memOut_CTf_f_Int_Int_Int_Int_r;
  MemOut_CTf_f_Int_Int_Int_Int_t memReadOut_CTf_f_Int_Int_Int_Int_d;
  logic memReadOut_CTf_f_Int_Int_Int_Int_r;
  MemOut_CTf_f_Int_Int_Int_Int_t memWriteOut_CTf_f_Int_Int_Int_Int_d;
  logic memWriteOut_CTf_f_Int_Int_Int_Int_r;
  MemIn_CTf_f_Int_Int_Int_Int_t memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d;
  logic memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_r;
  MemIn_CTf_f_Int_Int_Int_Int_t memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_d;
  logic memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_r;
  MemOut_CTf_f_Int_Int_Int_Int_t memOut_CTf_f_Int_Int_Int_Int_dbuf_d;
  logic memOut_CTf_f_Int_Int_Int_Int_dbuf_r;
  MemOut_CTf_f_Int_Int_Int_Int_t memOut_CTf_f_Int_Int_Int_Int_rbuf_d;
  logic memOut_CTf_f_Int_Int_Int_Int_rbuf_r;
  \Word16#_t  destructReadIn_CTf_f_Int_Int_Int_Int_d;
  logic destructReadIn_CTf_f_Int_Int_Int_Int_r;
  MemIn_CTf_f_Int_Int_Int_Int_t dconReadIn_CTf_f_Int_Int_Int_Int_d;
  logic dconReadIn_CTf_f_Int_Int_Int_Int_r;
  CTf_f_Int_Int_Int_Int_t readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_d;
  logic readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_r;
  C5_t writeMerge_choice_CTf_f_Int_Int_Int_Int_d;
  logic writeMerge_choice_CTf_f_Int_Int_Int_Int_r;
  CTf_f_Int_Int_Int_Int_t writeMerge_data_CTf_f_Int_Int_Int_Int_d;
  logic writeMerge_data_CTf_f_Int_Int_Int_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_r;
  MemIn_CTf_f_Int_Int_Int_Int_t dconWriteIn_CTf_f_Int_Int_Int_Int_d;
  logic dconWriteIn_CTf_f_Int_Int_Int_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t dconPtr_CTf_f_Int_Int_Int_Int_d;
  logic dconPtr_CTf_f_Int_Int_Int_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t _42_d;
  logic _42_r;
  assign _42_r = 1'd1;
  Pointer_CTf_f_Int_Int_Int_Int_t demuxWriteResult_CTf_f_Int_Int_Int_Int_d;
  logic demuxWriteResult_CTf_f_Int_Int_Int_Int_r;
  Go_t \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_r ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwstH_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_IntwstH_r ;
  Go_t go_7_1_d;
  logic go_7_1_r;
  Go_t go_7_2_d;
  logic go_7_2_r;
  Pointer_QTree_Int_t wstH_1_argbuf_d;
  logic wstH_1_argbuf_r;
  Int_t \es_7_1I#_d ;
  logic \es_7_1I#_r ;
  C2_t applyfnInt_Bool_5_choice_d;
  logic applyfnInt_Bool_5_choice_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5_data_d;
  logic applyfnInt_Bool_5_data_r;
  MyDTInt_Bool_t arg0_1_d;
  logic arg0_1_r;
  MyDTInt_Bool_t arg0_2_d;
  logic arg0_2_r;
  MyDTInt_Bool_t arg0_3_d;
  logic arg0_3_r;
  MyBool_t applyfnInt_Bool_5_resbuf_d;
  logic applyfnInt_Bool_5_resbuf_r;
  MyBool_t applyfnInt_Bool_5_2_argbuf_d;
  logic applyfnInt_Bool_5_2_argbuf_r;
  MyBool_t es_7_1_1_d;
  logic es_7_1_1_r;
  MyBool_t es_7_1_2_d;
  logic es_7_1_2_r;
  MyBool_t es_7_1_3_d;
  logic es_7_1_3_r;
  MyBool_t es_7_1_4_d;
  logic es_7_1_4_r;
  MyBool_t es_7_1_5_d;
  logic es_7_1_5_r;
  MyBool_t es_7_1_6_d;
  logic es_7_1_6_r;
  MyBool_t applyfnInt_Bool_5_1_d;
  logic applyfnInt_Bool_5_1_r;
  MyBool_t applyfnInt_Bool_5_2_d;
  logic applyfnInt_Bool_5_2_r;
  Go_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r;
  MyDTInt_Bool_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r;
  Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r;
  MyBool_t es_2_1_d;
  logic es_2_1_r;
  MyBool_t es_2_2_d;
  logic es_2_2_r;
  MyBool_t es_2_3_d;
  logic es_2_3_r;
  MyBool_t es_2_4_d;
  logic es_2_4_r;
  MyBool_t es_2_5_d;
  logic es_2_5_r;
  MyBool_t es_2_6_d;
  logic es_2_6_r;
  MyBool_t es_2_7_d;
  logic es_2_7_r;
  C2_t applyfnInt_Int_5_choice_d;
  logic applyfnInt_Int_5_choice_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5_data_d;
  logic applyfnInt_Int_5_data_r;
  MyDTInt_Int_t arg0_2_1_d;
  logic arg0_2_1_r;
  MyDTInt_Int_t arg0_2_2_d;
  logic arg0_2_2_r;
  MyDTInt_Int_t arg0_2_3_d;
  logic arg0_2_3_r;
  Int_t applyfnInt_Int_5_resbuf_d;
  logic applyfnInt_Int_5_resbuf_r;
  Int_t applyfnInt_Int_5_2_argbuf_d;
  logic applyfnInt_Int_5_2_argbuf_r;
  QTree_Int_t es_8_1QVal_Int_d;
  logic es_8_1QVal_Int_r;
  Int_t applyfnInt_Int_5_1_d;
  logic applyfnInt_Int_5_1_r;
  Int_t applyfnInt_Int_5_2_d;
  logic applyfnInt_Int_5_2_r;
  Go_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r;
  MyDTInt_Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r;
  Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r;
  Int_t es_4_1_1_argbuf_d;
  logic es_4_1_1_argbuf_r;
  C3_t applyfnInt_Int_Int_5_choice_d;
  logic applyfnInt_Int_Int_5_choice_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5_data_d;
  logic applyfnInt_Int_Int_5_data_r;
  MyDTInt_Int_Int_t arg0_4_1_d;
  logic arg0_4_1_r;
  MyDTInt_Int_Int_t arg0_4_2_d;
  logic arg0_4_2_r;
  MyDTInt_Int_Int_t arg0_4_3_d;
  logic arg0_4_3_r;
  Int_t applyfnInt_Int_Int_5_resbuf_d;
  logic applyfnInt_Int_Int_5_resbuf_r;
  Int_t applyfnInt_Int_Int_5_2_argbuf_d;
  logic applyfnInt_Int_Int_5_2_argbuf_r;
  Int_t es_6_1_1_argbuf_d;
  logic es_6_1_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_3_argbuf_d;
  logic applyfnInt_Int_Int_5_3_argbuf_r;
  Int_t es_10_1_argbuf_d;
  logic es_10_1_argbuf_r;
  Int_t applyfnInt_Int_Int_5_1_d;
  logic applyfnInt_Int_Int_5_1_r;
  Int_t applyfnInt_Int_Int_5_2_d;
  logic applyfnInt_Int_Int_5_2_r;
  Int_t applyfnInt_Int_Int_5_3_d;
  logic applyfnInt_Int_Int_5_3_r;
  MyDTInt_Int_Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r;
  Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r;
  Int_t es_1_1_argbuf_d;
  logic es_1_1_argbuf_r;
  Int_t arg0_1Dcon_eqZero_d;
  logic arg0_1Dcon_eqZero_r;
  Int_t arg0_1Dcon_eqZero_1_d;
  logic arg0_1Dcon_eqZero_1_r;
  Int_t arg0_1Dcon_eqZero_2_d;
  logic arg0_1Dcon_eqZero_2_r;
  Int_t arg0_1Dcon_eqZero_3_d;
  logic arg0_1Dcon_eqZero_3_r;
  Int_t arg0_1Dcon_eqZero_4_d;
  logic arg0_1Dcon_eqZero_4_r;
  \Int#_t  x1aph_destruct_d;
  logic x1aph_destruct_r;
  Int_t \arg0_1Dcon_eqZero_1I#_d ;
  logic \arg0_1Dcon_eqZero_1I#_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_d ;
  logic \arg0_1Dcon_eqZero_3I#_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_2_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_3_d ;
  logic \arg0_1Dcon_eqZero_3I#_3_r ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_argbuf_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_argbuf_r ;
  \Int#_t  \arg0_1Dcon_eqZero_3I#_1_argbuf_0_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ;
  Bool_t lizzieLet1_1wild1X19_1_Eq_d;
  logic lizzieLet1_1wild1X19_1_Eq_r;
  Go_t \arg0_1Dcon_eqZero_3I#_2_argbuf_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_argbuf_r ;
  TupGo___Bool_t boolConvert_1TupGo___Bool_1_d;
  logic boolConvert_1TupGo___Bool_1_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r;
  Go_t arg0_2Dcon_eqZero_d;
  logic arg0_2Dcon_eqZero_r;
  Int_t arg0_2_1Dcon_main1_d;
  logic arg0_2_1Dcon_main1_r;
  Int_t arg0_2_1Dcon_main1_1_d;
  logic arg0_2_1Dcon_main1_1_r;
  Int_t arg0_2_1Dcon_main1_2_d;
  logic arg0_2_1Dcon_main1_2_r;
  Int_t arg0_2_1Dcon_main1_3_d;
  logic arg0_2_1Dcon_main1_3_r;
  Int_t arg0_2_1Dcon_main1_4_d;
  logic arg0_2_1Dcon_main1_4_r;
  \Int#_t  xap7_destruct_d;
  logic xap7_destruct_r;
  Int_t \arg0_2_1Dcon_main1_1I#_d ;
  logic \arg0_2_1Dcon_main1_1I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_d ;
  logic \arg0_2_1Dcon_main1_3I#_r ;
  Go_t \arg0_2_1Dcon_main1_3I#_1_argbuf_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_r ;
  \Int#_t  \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d ;
  logic \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  Int_t \es_0_1_1I#_mux_d ;
  logic \es_0_1_1I#_mux_r ;
  Go_t arg0_2_2Dcon_main1_d;
  logic arg0_2_2Dcon_main1_r;
  Int_t \es_0_1_1I#_mux_mux_d ;
  logic \es_0_1_1I#_mux_mux_r ;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  Int_t \arg0_4_1Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_4_1Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_4_r ;
  \Int#_t  xa1m0_destruct_d;
  logic xa1m0_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r ;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r ;
  \Int#_t  ya1m1_destruct_d;
  logic ya1m1_destruct_r;
  Int_t \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ;
  \Int#_t  \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d ;
  logic \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r ;
  Int_t \es_0_2_1I#_d ;
  logic \es_0_2_1I#_r ;
  Int_t \es_0_2_1I#_mux_d ;
  logic \es_0_2_1I#_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_r ;
  Int_t \es_0_2_1I#_mux_mux_mux_d ;
  logic \es_0_2_1I#_mux_mux_mux_r ;
  Go_t boolConvert_1TupGo___Boolgo_1_d;
  logic boolConvert_1TupGo___Boolgo_1_r;
  Bool_t boolConvert_1TupGo___Boolbool_d;
  logic boolConvert_1TupGo___Boolbool_r;
  Bool_t bool_1_d;
  logic bool_1_r;
  Bool_t bool_2_d;
  logic bool_2_r;
  MyBool_t lizzieLet3_1_d;
  logic lizzieLet3_1_r;
  MyBool_t lizzieLet3_2_d;
  logic lizzieLet3_2_r;
  Go_t bool_1False_d;
  logic bool_1False_r;
  Go_t bool_1True_d;
  logic bool_1True_r;
  MyBool_t bool_1False_1MyFalse_d;
  logic bool_1False_1MyFalse_r;
  MyBool_t boolConvert_1_resbuf_d;
  logic boolConvert_1_resbuf_r;
  MyBool_t bool_1True_1MyTrue_d;
  logic bool_1True_1MyTrue_r;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_r;
  Go_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_r;
  Pointer_QTree_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r;
  Go_t call_$wnnz_Int_initBufi_d;
  logic call_$wnnz_Int_initBufi_r;
  C5_t go_10_goMux_choice_d;
  logic go_10_goMux_choice_r;
  Go_t go_10_goMux_data_d;
  logic go_10_goMux_data_r;
  Go_t call_$wnnz_Int_unlockFork1_d;
  logic call_$wnnz_Int_unlockFork1_r;
  Go_t call_$wnnz_Int_unlockFork2_d;
  logic call_$wnnz_Int_unlockFork2_r;
  Go_t call_$wnnz_Int_unlockFork3_d;
  logic call_$wnnz_Int_unlockFork3_r;
  Go_t call_$wnnz_Int_initBuf_d;
  logic call_$wnnz_Int_initBuf_r;
  Go_t call_$wnnz_Int_goMux1_d;
  logic call_$wnnz_Int_goMux1_r;
  Pointer_QTree_Int_t call_$wnnz_Int_goMux2_d;
  logic call_$wnnz_Int_goMux2_r;
  Pointer_CT$wnnz_Int_t call_$wnnz_Int_goMux3_d;
  logic call_$wnnz_Int_goMux3_r;
  Go_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_r ;
  Pointer_QTree_Int_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_r ;
  MyDTInt_Bool_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_r ;
  MyDTInt_Int_Int_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_r ;
  Int_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_r ;
  MyDTInt_Bool_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_r ;
  MyDTInt_Int_t \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_initBufi_d ;
  logic \call_f'_f'_Int_Int_Int_Int_initBufi_r ;
  C5_t go_11_goMux_choice_d;
  logic go_11_goMux_choice_r;
  Go_t go_11_goMux_data_d;
  logic go_11_goMux_data_r;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork1_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork1_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork2_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork2_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork3_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork3_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork4_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork4_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork5_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork5_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork6_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork6_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork7_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork7_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_unlockFork8_d ;
  logic \call_f'_f'_Int_Int_Int_Int_unlockFork8_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_initBuf_d ;
  logic \call_f'_f'_Int_Int_Int_Int_initBuf_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_goMux1_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux1_r ;
  Pointer_QTree_Int_t \call_f'_f'_Int_Int_Int_Int_goMux2_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux2_r ;
  MyDTInt_Bool_t \call_f'_f'_Int_Int_Int_Int_goMux3_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux3_r ;
  MyDTInt_Int_Int_t \call_f'_f'_Int_Int_Int_Int_goMux4_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux4_r ;
  Int_t \call_f'_f'_Int_Int_Int_Int_goMux5_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux5_r ;
  MyDTInt_Bool_t \call_f'_f'_Int_Int_Int_Int_goMux6_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux6_r ;
  MyDTInt_Int_t \call_f'_f'_Int_Int_Int_Int_goMux7_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux7_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \call_f'_f'_Int_Int_Int_Int_goMux8_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goMux8_r ;
  Go_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_r;
  MyDTInt_Bool_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_r;
  MyDTInt_Int_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_r;
  MyDTInt_Bool_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_r;
  MyDTInt_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_r;
  Pointer_CTf_f_Int_Int_Int_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_r;
  Go_t call_f_f_Int_Int_Int_Int_initBufi_d;
  logic call_f_f_Int_Int_Int_Int_initBufi_r;
  C5_t go_12_goMux_choice_d;
  logic go_12_goMux_choice_r;
  Go_t go_12_goMux_data_d;
  logic go_12_goMux_data_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork1_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork1_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork2_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork2_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork3_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork3_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork4_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork4_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork5_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork5_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork6_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork6_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork7_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork7_r;
  Go_t call_f_f_Int_Int_Int_Int_unlockFork8_d;
  logic call_f_f_Int_Int_Int_Int_unlockFork8_r;
  Go_t call_f_f_Int_Int_Int_Int_initBuf_d;
  logic call_f_f_Int_Int_Int_Int_initBuf_r;
  Go_t call_f_f_Int_Int_Int_Int_goMux1_d;
  logic call_f_f_Int_Int_Int_Int_goMux1_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_Int_Int_goMux2_d;
  logic call_f_f_Int_Int_Int_Int_goMux2_r;
  Pointer_QTree_Int_t call_f_f_Int_Int_Int_Int_goMux3_d;
  logic call_f_f_Int_Int_Int_Int_goMux3_r;
  MyDTInt_Bool_t call_f_f_Int_Int_Int_Int_goMux4_d;
  logic call_f_f_Int_Int_Int_Int_goMux4_r;
  MyDTInt_Int_Int_t call_f_f_Int_Int_Int_Int_goMux5_d;
  logic call_f_f_Int_Int_Int_Int_goMux5_r;
  MyDTInt_Bool_t call_f_f_Int_Int_Int_Int_goMux6_d;
  logic call_f_f_Int_Int_Int_Int_goMux6_r;
  MyDTInt_Int_t call_f_f_Int_Int_Int_Int_goMux7_d;
  logic call_f_f_Int_Int_Int_Int_goMux7_r;
  Pointer_CTf_f_Int_Int_Int_Int_t call_f_f_Int_Int_Int_Int_goMux8_d;
  logic call_f_f_Int_Int_Int_Int_goMux8_r;
  MyDTInt_Int_t es_2_1MyFalse_d;
  logic es_2_1MyFalse_r;
  MyDTInt_Int_t _41_d;
  logic _41_r;
  assign _41_r = 1'd1;
  MyDTInt_Int_t es_2_1MyFalse_1_d;
  logic es_2_1MyFalse_1_r;
  MyDTInt_Int_t es_2_1MyFalse_2_d;
  logic es_2_1MyFalse_2_r;
  MyDTInt_Int_t es_2_1MyFalse_1_argbuf_d;
  logic es_2_1MyFalse_1_argbuf_r;
  Go_t es_2_2MyFalse_d;
  logic es_2_2MyFalse_r;
  Go_t es_2_2MyTrue_d;
  logic es_2_2MyTrue_r;
  Go_t es_2_2MyFalse_1_d;
  logic es_2_2MyFalse_1_r;
  Go_t es_2_2MyFalse_2_d;
  logic es_2_2MyFalse_2_r;
  Go_t es_2_2MyFalse_3_d;
  logic es_2_2MyFalse_3_r;
  Go_t es_2_2MyFalse_1_argbuf_d;
  logic es_2_2MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r;
  Go_t es_2_2MyFalse_2_argbuf_d;
  logic es_2_2MyFalse_2_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r;
  Go_t es_2_2MyTrue_1_d;
  logic es_2_2MyTrue_1_r;
  Go_t es_2_2MyTrue_2_d;
  logic es_2_2MyTrue_2_r;
  QTree_Int_t es_2_2MyTrue_1QNone_Int_d;
  logic es_2_2MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet10_1_argbuf_d;
  logic lizzieLet10_1_argbuf_r;
  Go_t es_2_2MyTrue_2_argbuf_d;
  logic es_2_2MyTrue_2_argbuf_r;
  MyDTInt_Bool_t es_2_3MyFalse_d;
  logic es_2_3MyFalse_r;
  MyDTInt_Bool_t _40_d;
  logic _40_r;
  assign _40_r = 1'd1;
  MyDTInt_Bool_t es_2_3MyFalse_1_argbuf_d;
  logic es_2_3MyFalse_1_argbuf_r;
  MyDTInt_Int_Int_t es_2_4MyFalse_d;
  logic es_2_4MyFalse_r;
  MyDTInt_Int_Int_t _39_d;
  logic _39_r;
  assign _39_r = 1'd1;
  MyDTInt_Int_Int_t es_2_4MyFalse_1_d;
  logic es_2_4MyFalse_1_r;
  MyDTInt_Int_Int_t es_2_4MyFalse_2_d;
  logic es_2_4MyFalse_2_r;
  MyDTInt_Int_Int_t es_2_4MyFalse_1_argbuf_d;
  logic es_2_4MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_2_5MyFalse_d;
  logic es_2_5MyFalse_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_2_5MyTrue_d;
  logic es_2_5MyTrue_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_2_5MyTrue_1_argbuf_d;
  logic es_2_5MyTrue_1_argbuf_r;
  Int_t es_2_6MyFalse_d;
  logic es_2_6MyFalse_r;
  Int_t _38_d;
  logic _38_r;
  assign _38_r = 1'd1;
  Int_t es_2_6MyFalse_1_d;
  logic es_2_6MyFalse_1_r;
  Int_t es_2_6MyFalse_2_d;
  logic es_2_6MyFalse_2_r;
  Int_t es_2_6MyFalse_1_argbuf_d;
  logic es_2_6MyFalse_1_argbuf_r;
  Int_t es_2_7MyFalse_d;
  logic es_2_7MyFalse_r;
  Int_t _37_d;
  logic _37_r;
  assign _37_r = 1'd1;
  Int_t es_2_7MyFalse_1_d;
  logic es_2_7MyFalse_1_r;
  Int_t es_2_7MyFalse_2_d;
  logic es_2_7MyFalse_2_r;
  Int_t es_2_7MyFalse_1_argbuf_d;
  logic es_2_7MyFalse_1_argbuf_r;
  \Int#_t  contRet_0_1_argbuf_d;
  logic contRet_0_1_argbuf_r;
  \Int#_t  es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_d;
  logic es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_r;
  MyDTInt_Int_t es_7_1_1MyFalse_d;
  logic es_7_1_1MyFalse_r;
  MyDTInt_Int_t _36_d;
  logic _36_r;
  assign _36_r = 1'd1;
  MyDTInt_Int_t es_7_1_1MyFalse_1_argbuf_d;
  logic es_7_1_1MyFalse_1_argbuf_r;
  Go_t es_7_1_2MyFalse_d;
  logic es_7_1_2MyFalse_r;
  Go_t es_7_1_2MyTrue_d;
  logic es_7_1_2MyTrue_r;
  Go_t es_7_1_2MyFalse_1_d;
  logic es_7_1_2MyFalse_1_r;
  Go_t es_7_1_2MyFalse_2_d;
  logic es_7_1_2MyFalse_2_r;
  Go_t es_7_1_2MyFalse_1_argbuf_d;
  logic es_7_1_2MyFalse_1_argbuf_r;
  TupGo___MyDTInt_Int___Int_t applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d;
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r;
  Go_t es_7_1_2MyFalse_2_argbuf_d;
  logic es_7_1_2MyFalse_2_argbuf_r;
  Go_t es_7_1_2MyTrue_1_d;
  logic es_7_1_2MyTrue_1_r;
  Go_t es_7_1_2MyTrue_2_d;
  logic es_7_1_2MyTrue_2_r;
  QTree_Int_t es_7_1_2MyTrue_1QNone_Int_d;
  logic es_7_1_2MyTrue_1QNone_Int_r;
  QTree_Int_t lizzieLet9_1_argbuf_d;
  logic lizzieLet9_1_argbuf_r;
  Go_t es_7_1_2MyTrue_2_argbuf_d;
  logic es_7_1_2MyTrue_2_argbuf_r;
  MyDTInt_Int_Int_t es_7_1_3MyFalse_d;
  logic es_7_1_3MyFalse_r;
  MyDTInt_Int_Int_t _35_d;
  logic _35_r;
  assign _35_r = 1'd1;
  MyDTInt_Int_Int_t es_7_1_3MyFalse_1_argbuf_d;
  logic es_7_1_3MyFalse_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyFalse_d;
  logic es_7_1_4MyFalse_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyTrue_d;
  logic es_7_1_4MyTrue_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyFalse_1_argbuf_d;
  logic es_7_1_4MyFalse_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyTrue_1_argbuf_d;
  logic es_7_1_4MyTrue_1_argbuf_r;
  Int_t es_7_1_5MyFalse_d;
  logic es_7_1_5MyFalse_r;
  Int_t _34_d;
  logic _34_r;
  assign _34_r = 1'd1;
  Int_t es_7_1_5MyFalse_1_argbuf_d;
  logic es_7_1_5MyFalse_1_argbuf_r;
  Int_t es_7_1_6MyFalse_d;
  logic es_7_1_6MyFalse_r;
  Int_t _33_d;
  logic _33_r;
  assign _33_r = 1'd1;
  Int_t es_7_1_6MyFalse_1_argbuf_d;
  logic es_7_1_6MyFalse_1_argbuf_r;
  QTree_Int_t lizzieLet8_1_argbuf_d;
  logic lizzieLet8_1_argbuf_r;
  Go_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_r ;
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_r ;
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_r ;
  MyDTInt_Int_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_r ;
  Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_r ;
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_r ;
  MyDTInt_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_r ;
  MyDTInt_Int_t f_mapaia_1_1_argbuf_d;
  logic f_mapaia_1_1_argbuf_r;
  Go_t go_13_1_d;
  logic go_13_1_r;
  Go_t go_13_2_d;
  logic go_13_2_r;
  MyDTInt_Bool_t is_z_kronai6_1_1_argbuf_d;
  logic is_z_kronai6_1_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapai9_1_1_argbuf_d;
  logic is_z_mapai9_1_1_argbuf_r;
  Pointer_QTree_Int_t m2ai5_1_1_argbuf_d;
  logic m2ai5_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_kronai7_1_1_argbuf_d;
  logic op_kronai7_1_1_argbuf_r;
  Int_t vai8_1_1_argbuf_d;
  logic vai8_1_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet8_1_1_argbuf_d;
  logic lizzieLet8_1_1_argbuf_r;
  Go_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_r;
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_r;
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_r;
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_r;
  MyDTInt_Int_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_r;
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_r;
  MyDTInt_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_r;
  MyDTInt_Int_t f_mapahZ_1_1_argbuf_d;
  logic f_mapahZ_1_1_argbuf_r;
  Go_t go_14_1_d;
  logic go_14_1_r;
  Go_t go_14_2_d;
  logic go_14_2_r;
  MyDTInt_Bool_t is_z_kronahW_1_1_argbuf_d;
  logic is_z_kronahW_1_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapahY_1_1_argbuf_d;
  logic is_z_mapahY_1_1_argbuf_r;
  Pointer_QTree_Int_t m1ahU_1_1_argbuf_d;
  logic m1ahU_1_1_argbuf_r;
  Pointer_QTree_Int_t m2ahV_1_1_argbuf_d;
  logic m2ahV_1_1_argbuf_r;
  MyDTInt_Int_Int_t op_kronahX_1_1_argbuf_d;
  logic op_kronahX_1_1_argbuf_r;
  Pointer_QTree_Int_t es_0_1_argbuf_d;
  logic es_0_1_argbuf_r;
  MyDTInt_Int_t f_mapahZ_2_2_argbuf_d;
  logic f_mapahZ_2_2_argbuf_r;
  MyDTInt_Int_t f_mapahZ_2_1_d;
  logic f_mapahZ_2_1_r;
  MyDTInt_Int_t f_mapahZ_2_2_d;
  logic f_mapahZ_2_2_r;
  MyDTInt_Int_t f_mapahZ_3_2_argbuf_d;
  logic f_mapahZ_3_2_argbuf_r;
  MyDTInt_Int_t f_mapahZ_3_1_d;
  logic f_mapahZ_3_1_r;
  MyDTInt_Int_t f_mapahZ_3_2_d;
  logic f_mapahZ_3_2_r;
  MyDTInt_Int_t f_mapahZ_4_1_argbuf_d;
  logic f_mapahZ_4_1_argbuf_r;
  MyDTInt_Int_t f_mapaia_2_2_argbuf_d;
  logic f_mapaia_2_2_argbuf_r;
  MyDTInt_Int_t f_mapaia_2_1_d;
  logic f_mapaia_2_1_r;
  MyDTInt_Int_t f_mapaia_2_2_d;
  logic f_mapaia_2_2_r;
  MyDTInt_Int_t f_mapaia_3_2_argbuf_d;
  logic f_mapaia_3_2_argbuf_r;
  MyDTInt_Int_t f_mapaia_3_1_d;
  logic f_mapaia_3_1_r;
  MyDTInt_Int_t f_mapaia_3_2_d;
  logic f_mapaia_3_2_r;
  MyDTInt_Int_t f_mapaia_4_1_argbuf_d;
  logic f_mapaia_4_1_argbuf_r;
  MyDTInt_Int_t go_1Dcon_main1_d;
  logic go_1Dcon_main1_r;
  C5_t go_10_goMux_choice_1_d;
  logic go_10_goMux_choice_1_r;
  C5_t go_10_goMux_choice_2_d;
  logic go_10_goMux_choice_2_r;
  Pointer_QTree_Int_t wstH_1_goMux_mux_d;
  logic wstH_1_goMux_mux_r;
  Pointer_CT$wnnz_Int_t sc_0_goMux_mux_d;
  logic sc_0_goMux_mux_r;
  C5_t go_11_goMux_choice_1_d;
  logic go_11_goMux_choice_1_r;
  C5_t go_11_goMux_choice_2_d;
  logic go_11_goMux_choice_2_r;
  C5_t go_11_goMux_choice_3_d;
  logic go_11_goMux_choice_3_r;
  C5_t go_11_goMux_choice_4_d;
  logic go_11_goMux_choice_4_r;
  C5_t go_11_goMux_choice_5_d;
  logic go_11_goMux_choice_5_r;
  C5_t go_11_goMux_choice_6_d;
  logic go_11_goMux_choice_6_r;
  C5_t go_11_goMux_choice_7_d;
  logic go_11_goMux_choice_7_r;
  Pointer_QTree_Int_t m2ai5_goMux_mux_d;
  logic m2ai5_goMux_mux_r;
  MyDTInt_Bool_t is_z_kronai6_goMux_mux_d;
  logic is_z_kronai6_goMux_mux_r;
  MyDTInt_Int_Int_t op_kronai7_goMux_mux_d;
  logic op_kronai7_goMux_mux_r;
  Int_t vai8_goMux_mux_d;
  logic vai8_goMux_mux_r;
  MyDTInt_Bool_t is_z_mapai9_goMux_mux_d;
  logic is_z_mapai9_goMux_mux_r;
  MyDTInt_Int_t f_mapaia_goMux_mux_d;
  logic f_mapaia_goMux_mux_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_1_goMux_mux_d;
  logic sc_0_1_goMux_mux_r;
  C5_t go_12_goMux_choice_1_d;
  logic go_12_goMux_choice_1_r;
  C5_t go_12_goMux_choice_2_d;
  logic go_12_goMux_choice_2_r;
  C5_t go_12_goMux_choice_3_d;
  logic go_12_goMux_choice_3_r;
  C5_t go_12_goMux_choice_4_d;
  logic go_12_goMux_choice_4_r;
  C5_t go_12_goMux_choice_5_d;
  logic go_12_goMux_choice_5_r;
  C5_t go_12_goMux_choice_6_d;
  logic go_12_goMux_choice_6_r;
  C5_t go_12_goMux_choice_7_d;
  logic go_12_goMux_choice_7_r;
  Pointer_QTree_Int_t m1ahU_goMux_mux_d;
  logic m1ahU_goMux_mux_r;
  Pointer_QTree_Int_t m2ahV_goMux_mux_d;
  logic m2ahV_goMux_mux_r;
  MyDTInt_Bool_t is_z_kronahW_goMux_mux_d;
  logic is_z_kronahW_goMux_mux_r;
  MyDTInt_Int_Int_t op_kronahX_goMux_mux_d;
  logic op_kronahX_goMux_mux_r;
  MyDTInt_Bool_t is_z_mapahY_goMux_mux_d;
  logic is_z_mapahY_goMux_mux_r;
  MyDTInt_Int_t f_mapahZ_goMux_mux_d;
  logic f_mapahZ_goMux_mux_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_2_goMux_mux_d;
  logic sc_0_2_goMux_mux_r;
  \CTf'_f'_Int_Int_Int_Int_t  \go_13_1Lf'_f'_Int_Int_Int_Intsbos_d ;
  logic \go_13_1Lf'_f'_Int_Int_Int_Intsbos_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet17_1_argbuf_d;
  logic lizzieLet17_1_argbuf_r;
  Go_t go_13_2_argbuf_d;
  logic go_13_2_argbuf_r;
  \TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_t  \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d ;
  logic \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_r ;
  CTf_f_Int_Int_Int_Int_t go_14_1Lf_f_Int_Int_Int_Intsbos_d;
  logic go_14_1Lf_f_Int_Int_Int_Intsbos_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet18_1_argbuf_d;
  logic lizzieLet18_1_argbuf_r;
  Go_t go_14_2_argbuf_d;
  logic go_14_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_t call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d;
  logic call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_r;
  C4_t go_15_goMux_choice_1_d;
  logic go_15_goMux_choice_1_r;
  C4_t go_15_goMux_choice_2_d;
  logic go_15_goMux_choice_2_r;
  \Int#_t  srtarg_0_goMux_mux_d;
  logic srtarg_0_goMux_mux_r;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_d;
  logic scfarg_0_goMux_mux_r;
  C6_t go_16_goMux_choice_1_d;
  logic go_16_goMux_choice_1_r;
  C6_t go_16_goMux_choice_2_d;
  logic go_16_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_1_goMux_mux_d;
  logic srtarg_0_1_goMux_mux_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  scfarg_0_1_goMux_mux_d;
  logic scfarg_0_1_goMux_mux_r;
  C4_t go_17_goMux_choice_1_d;
  logic go_17_goMux_choice_1_r;
  C4_t go_17_goMux_choice_2_d;
  logic go_17_goMux_choice_2_r;
  Pointer_QTree_Int_t srtarg_0_2_goMux_mux_d;
  logic srtarg_0_2_goMux_mux_r;
  Pointer_CTf_f_Int_Int_Int_Int_t scfarg_0_2_goMux_mux_d;
  logic scfarg_0_2_goMux_mux_r;
  MyDTInt_Int_t es_6_1_argbuf_d;
  logic es_6_1_argbuf_r;
  MyDTInt_Bool_t go_2Dcon_eqZero_d;
  logic go_2Dcon_eqZero_r;
  MyDTInt_Bool_t es_5_1_argbuf_d;
  logic es_5_1_argbuf_r;
  MyDTInt_Int_Int_t \go_3Dcon_$fNumInt_$ctimes_d ;
  logic \go_3Dcon_$fNumInt_$ctimes_r ;
  MyDTInt_Int_Int_t es_4_1_argbuf_d;
  logic es_4_1_argbuf_r;
  MyDTInt_Bool_t go_4Dcon_eqZero_d;
  logic go_4Dcon_eqZero_r;
  MyDTInt_Bool_t es_3_1_argbuf_d;
  logic es_3_1_argbuf_r;
  Go_t go_5_argbuf_d;
  logic go_5_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_r;
  Go_t go_6_argbuf_d;
  logic go_6_argbuf_r;
  TupGo___Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_Int_1_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_Int_1_r ;
  CT$wnnz_Int_t go_7_1L$wnnz_Intsbos_d;
  logic go_7_1L$wnnz_Intsbos_r;
  CT$wnnz_Int_t lizzieLet0_1_argbuf_d;
  logic lizzieLet0_1_argbuf_r;
  Go_t go_7_2_argbuf_d;
  logic go_7_2_argbuf_r;
  TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_t call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d;
  logic call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r;
  MyDTInt_Bool_t is_z_kronahW_2_2_argbuf_d;
  logic is_z_kronahW_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_kronahW_2_1_d;
  logic is_z_kronahW_2_1_r;
  MyDTInt_Bool_t is_z_kronahW_2_2_d;
  logic is_z_kronahW_2_2_r;
  MyDTInt_Bool_t is_z_kronahW_3_2_argbuf_d;
  logic is_z_kronahW_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_kronahW_3_1_d;
  logic is_z_kronahW_3_1_r;
  MyDTInt_Bool_t is_z_kronahW_3_2_d;
  logic is_z_kronahW_3_2_r;
  MyDTInt_Bool_t is_z_kronahW_4_1_argbuf_d;
  logic is_z_kronahW_4_1_argbuf_r;
  MyDTInt_Bool_t is_z_kronai6_2_2_argbuf_d;
  logic is_z_kronai6_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_kronai6_2_1_d;
  logic is_z_kronai6_2_1_r;
  MyDTInt_Bool_t is_z_kronai6_2_2_d;
  logic is_z_kronai6_2_2_r;
  MyDTInt_Bool_t is_z_kronai6_3_2_argbuf_d;
  logic is_z_kronai6_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_kronai6_3_1_d;
  logic is_z_kronai6_3_1_r;
  MyDTInt_Bool_t is_z_kronai6_3_2_d;
  logic is_z_kronai6_3_2_r;
  MyDTInt_Bool_t is_z_kronai6_4_1_argbuf_d;
  logic is_z_kronai6_4_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapahY_2_2_argbuf_d;
  logic is_z_mapahY_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapahY_2_1_d;
  logic is_z_mapahY_2_1_r;
  MyDTInt_Bool_t is_z_mapahY_2_2_d;
  logic is_z_mapahY_2_2_r;
  MyDTInt_Bool_t is_z_mapahY_3_2_argbuf_d;
  logic is_z_mapahY_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapahY_3_1_d;
  logic is_z_mapahY_3_1_r;
  MyDTInt_Bool_t is_z_mapahY_3_2_d;
  logic is_z_mapahY_3_2_r;
  MyDTInt_Bool_t is_z_mapahY_4_1_argbuf_d;
  logic is_z_mapahY_4_1_argbuf_r;
  MyDTInt_Bool_t is_z_mapai9_2_2_argbuf_d;
  logic is_z_mapai9_2_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapai9_2_1_d;
  logic is_z_mapai9_2_1_r;
  MyDTInt_Bool_t is_z_mapai9_2_2_d;
  logic is_z_mapai9_2_2_r;
  MyDTInt_Bool_t is_z_mapai9_3_2_argbuf_d;
  logic is_z_mapai9_3_2_argbuf_r;
  MyDTInt_Bool_t is_z_mapai9_3_1_d;
  logic is_z_mapai9_3_1_r;
  MyDTInt_Bool_t is_z_mapai9_3_2_d;
  logic is_z_mapai9_3_2_r;
  MyDTInt_Bool_t is_z_mapai9_4_1_argbuf_d;
  logic is_z_mapai9_4_1_argbuf_r;
  Pointer_QTree_Int_t q1ai1_destruct_d;
  logic q1ai1_destruct_r;
  Pointer_QTree_Int_t q2ai2_destruct_d;
  logic q2ai2_destruct_r;
  Pointer_QTree_Int_t q3ai3_destruct_d;
  logic q3ai3_destruct_r;
  Pointer_QTree_Int_t q4ai4_destruct_d;
  logic q4ai4_destruct_r;
  Int_t vai0_destruct_d;
  logic vai0_destruct_r;
  QTree_Int_t _32_d;
  logic _32_r;
  assign _32_r = 1'd1;
  QTree_Int_t lizzieLet13_1_1QVal_Int_d;
  logic lizzieLet13_1_1QVal_Int_r;
  QTree_Int_t lizzieLet13_1_1QNode_Int_d;
  logic lizzieLet13_1_1QNode_Int_r;
  QTree_Int_t _31_d;
  logic _31_r;
  assign _31_r = 1'd1;
  MyDTInt_Int_t _30_d;
  logic _30_r;
  assign _30_r = 1'd1;
  MyDTInt_Int_t lizzieLet13_1_3QVal_Int_d;
  logic lizzieLet13_1_3QVal_Int_r;
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_d;
  logic lizzieLet13_1_3QNode_Int_r;
  MyDTInt_Int_t _29_d;
  logic _29_r;
  assign _29_r = 1'd1;
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_1_d;
  logic lizzieLet13_1_3QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_2_d;
  logic lizzieLet13_1_3QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_2_argbuf_d;
  logic lizzieLet13_1_3QNode_Int_2_argbuf_r;
  MyDTInt_Int_t lizzieLet13_1_3QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_3QVal_Int_1_argbuf_r;
  Go_t lizzieLet13_1_4QNone_Int_d;
  logic lizzieLet13_1_4QNone_Int_r;
  Go_t lizzieLet13_1_4QVal_Int_d;
  logic lizzieLet13_1_4QVal_Int_r;
  Go_t lizzieLet13_1_4QNode_Int_d;
  logic lizzieLet13_1_4QNode_Int_r;
  Go_t lizzieLet13_1_4QError_Int_d;
  logic lizzieLet13_1_4QError_Int_r;
  Go_t lizzieLet13_1_4QError_Int_1_d;
  logic lizzieLet13_1_4QError_Int_1_r;
  Go_t lizzieLet13_1_4QError_Int_2_d;
  logic lizzieLet13_1_4QError_Int_2_r;
  QTree_Int_t lizzieLet13_1_4QError_Int_1QError_Int_d;
  logic lizzieLet13_1_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet16_1_argbuf_d;
  logic lizzieLet16_1_argbuf_r;
  Go_t lizzieLet13_1_4QError_Int_2_argbuf_d;
  logic lizzieLet13_1_4QError_Int_2_argbuf_r;
  Go_t lizzieLet13_1_4QNode_Int_1_argbuf_d;
  logic lizzieLet13_1_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet13_1_4QNone_Int_1_d;
  logic lizzieLet13_1_4QNone_Int_1_r;
  Go_t lizzieLet13_1_4QNone_Int_2_d;
  logic lizzieLet13_1_4QNone_Int_2_r;
  QTree_Int_t lizzieLet13_1_4QNone_Int_1QNone_Int_d;
  logic lizzieLet13_1_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet14_1_argbuf_d;
  logic lizzieLet14_1_argbuf_r;
  Go_t lizzieLet13_1_4QNone_Int_2_argbuf_d;
  logic lizzieLet13_1_4QNone_Int_2_argbuf_r;
  C4_t go_17_goMux_choice_d;
  logic go_17_goMux_choice_r;
  Go_t go_17_goMux_data_d;
  logic go_17_goMux_data_r;
  Go_t lizzieLet13_1_4QVal_Int_1_d;
  logic lizzieLet13_1_4QVal_Int_1_r;
  Go_t lizzieLet13_1_4QVal_Int_2_d;
  logic lizzieLet13_1_4QVal_Int_2_r;
  Go_t lizzieLet13_1_4QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_4QVal_Int_1_argbuf_r;
  TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_r ;
  Go_t lizzieLet13_1_4QVal_Int_2_argbuf_d;
  logic lizzieLet13_1_4QVal_Int_2_argbuf_r;
  MyDTInt_Bool_t _28_d;
  logic _28_r;
  assign _28_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_1_5QVal_Int_d;
  logic lizzieLet13_1_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_d;
  logic lizzieLet13_1_5QNode_Int_r;
  MyDTInt_Bool_t _27_d;
  logic _27_r;
  assign _27_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_1_d;
  logic lizzieLet13_1_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_2_d;
  logic lizzieLet13_1_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_2_argbuf_d;
  logic lizzieLet13_1_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet13_1_5QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_5QVal_Int_1_argbuf_r;
  MyDTInt_Bool_t _26_d;
  logic _26_r;
  assign _26_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_1_6QVal_Int_d;
  logic lizzieLet13_1_6QVal_Int_r;
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_d;
  logic lizzieLet13_1_6QNode_Int_r;
  MyDTInt_Bool_t _25_d;
  logic _25_r;
  assign _25_r = 1'd1;
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_1_d;
  logic lizzieLet13_1_6QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_2_d;
  logic lizzieLet13_1_6QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_2_argbuf_d;
  logic lizzieLet13_1_6QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet13_1_6QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_6QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t _24_d;
  logic _24_r;
  assign _24_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_1_7QVal_Int_d;
  logic lizzieLet13_1_7QVal_Int_r;
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_d;
  logic lizzieLet13_1_7QNode_Int_r;
  Pointer_QTree_Int_t _23_d;
  logic _23_r;
  assign _23_r = 1'd1;
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_1_d;
  logic lizzieLet13_1_7QNode_Int_1_r;
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_2_d;
  logic lizzieLet13_1_7QNode_Int_2_r;
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_2_argbuf_d;
  logic lizzieLet13_1_7QNode_Int_2_argbuf_r;
  Pointer_QTree_Int_t lizzieLet13_1_7QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_7QVal_Int_1_argbuf_r;
  MyDTInt_Int_Int_t _22_d;
  logic _22_r;
  assign _22_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_1_8QVal_Int_d;
  logic lizzieLet13_1_8QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_d;
  logic lizzieLet13_1_8QNode_Int_r;
  MyDTInt_Int_Int_t _21_d;
  logic _21_r;
  assign _21_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_1_d;
  logic lizzieLet13_1_8QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_2_d;
  logic lizzieLet13_1_8QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_2_argbuf_d;
  logic lizzieLet13_1_8QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet13_1_8QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_8QVal_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNone_Int_d;
  logic lizzieLet13_1_9QNone_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QVal_Int_d;
  logic lizzieLet13_1_9QVal_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNode_Int_d;
  logic lizzieLet13_1_9QNode_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QError_Int_d;
  logic lizzieLet13_1_9QError_Int_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QError_Int_1_argbuf_d;
  logic lizzieLet13_1_9QError_Int_1_argbuf_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_d;
  logic lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet15_1_argbuf_d;
  logic lizzieLet15_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNone_Int_1_argbuf_d;
  logic lizzieLet13_1_9QNone_Int_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QVal_Int_1_argbuf_d;
  logic lizzieLet13_1_9QVal_Int_1_argbuf_r;
  \Int#_t  wwstK_4_destruct_d;
  logic wwstK_4_destruct_r;
  \Int#_t  ww1XuL_2_destruct_d;
  logic ww1XuL_2_destruct_r;
  \Int#_t  ww2XuO_1_destruct_d;
  logic ww2XuO_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_d;
  logic sc_0_6_destruct_r;
  \Int#_t  wwstK_3_destruct_d;
  logic wwstK_3_destruct_r;
  \Int#_t  ww1XuL_1_destruct_d;
  logic ww1XuL_1_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_5_destruct_d;
  logic sc_0_5_destruct_r;
  Pointer_QTree_Int_t q4abZ_3_destruct_d;
  logic q4abZ_3_destruct_r;
  \Int#_t  wwstK_2_destruct_d;
  logic wwstK_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_4_destruct_d;
  logic sc_0_4_destruct_r;
  Pointer_QTree_Int_t q4abZ_2_destruct_d;
  logic q4abZ_2_destruct_r;
  Pointer_QTree_Int_t q3abY_2_destruct_d;
  logic q3abY_2_destruct_r;
  Pointer_CT$wnnz_Int_t sc_0_3_destruct_d;
  logic sc_0_3_destruct_r;
  Pointer_QTree_Int_t q4abZ_1_destruct_d;
  logic q4abZ_1_destruct_r;
  Pointer_QTree_Int_t q3abY_1_destruct_d;
  logic q3abY_1_destruct_r;
  Pointer_QTree_Int_t q2abX_1_destruct_d;
  logic q2abX_1_destruct_r;
  CT$wnnz_Int_t _20_d;
  logic _20_r;
  assign _20_r = 1'd1;
  CT$wnnz_Int_t lizzieLet19_1Lcall_$wnnz_Int3_d;
  logic lizzieLet19_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet19_1Lcall_$wnnz_Int2_d;
  logic lizzieLet19_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet19_1Lcall_$wnnz_Int1_d;
  logic lizzieLet19_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet19_1Lcall_$wnnz_Int0_d;
  logic lizzieLet19_1Lcall_$wnnz_Int0_r;
  Go_t _19_d;
  logic _19_r;
  assign _19_r = 1'd1;
  Go_t lizzieLet19_3Lcall_$wnnz_Int3_d;
  logic lizzieLet19_3Lcall_$wnnz_Int3_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int2_d;
  logic lizzieLet19_3Lcall_$wnnz_Int2_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int1_d;
  logic lizzieLet19_3Lcall_$wnnz_Int1_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int0_d;
  logic lizzieLet19_3Lcall_$wnnz_Int0_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_r;
  Go_t lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_d;
  logic lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_r;
  \Int#_t  lizzieLet19_4L$wnnz_Intsbos_d;
  logic lizzieLet19_4L$wnnz_Intsbos_r;
  \Int#_t  lizzieLet19_4Lcall_$wnnz_Int3_d;
  logic lizzieLet19_4Lcall_$wnnz_Int3_r;
  \Int#_t  lizzieLet19_4Lcall_$wnnz_Int2_d;
  logic lizzieLet19_4Lcall_$wnnz_Int2_r;
  \Int#_t  lizzieLet19_4Lcall_$wnnz_Int1_d;
  logic lizzieLet19_4Lcall_$wnnz_Int1_r;
  \Int#_t  lizzieLet19_4Lcall_$wnnz_Int0_d;
  logic lizzieLet19_4Lcall_$wnnz_Int0_r;
  \Int#_t  lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_r;
  \Int#_t  lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_$wnnz_Int_goConst_d;
  logic call_$wnnz_Int_goConst_r;
  \Int#_t  \$wnnz_Int_resbuf_d ;
  logic \$wnnz_Int_resbuf_r ;
  CT$wnnz_Int_t lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_d;
  logic lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_r;
  CT$wnnz_Int_t lizzieLet20_1_argbuf_d;
  logic lizzieLet20_1_argbuf_r;
  Bool_t lizzieLet2_1_argbuf_d;
  logic lizzieLet2_1_argbuf_r;
  Pointer_QTree_Int_t es_12_destruct_d;
  logic es_12_destruct_r;
  Pointer_QTree_Int_t es_13_1_destruct_d;
  logic es_13_1_destruct_r;
  Pointer_QTree_Int_t es_14_2_destruct_d;
  logic es_14_2_destruct_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_10_destruct_d;
  logic sc_0_10_destruct_r;
  Pointer_QTree_Int_t es_13_destruct_d;
  logic es_13_destruct_r;
  Pointer_QTree_Int_t es_14_1_destruct_d;
  logic es_14_1_destruct_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_9_destruct_d;
  logic sc_0_9_destruct_r;
  Pointer_QTree_Int_t q1aic_3_destruct_d;
  logic q1aic_3_destruct_r;
  MyDTInt_Bool_t is_z_kronai6_4_destruct_d;
  logic is_z_kronai6_4_destruct_r;
  MyDTInt_Int_Int_t op_kronai7_4_destruct_d;
  logic op_kronai7_4_destruct_r;
  Int_t vai8_4_destruct_d;
  logic vai8_4_destruct_r;
  MyDTInt_Bool_t is_z_mapai9_4_destruct_d;
  logic is_z_mapai9_4_destruct_r;
  MyDTInt_Int_t f_mapaia_4_destruct_d;
  logic f_mapaia_4_destruct_r;
  Pointer_QTree_Int_t es_14_destruct_d;
  logic es_14_destruct_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_8_destruct_d;
  logic sc_0_8_destruct_r;
  Pointer_QTree_Int_t q1aic_2_destruct_d;
  logic q1aic_2_destruct_r;
  MyDTInt_Bool_t is_z_kronai6_3_destruct_d;
  logic is_z_kronai6_3_destruct_r;
  MyDTInt_Int_Int_t op_kronai7_3_destruct_d;
  logic op_kronai7_3_destruct_r;
  Int_t vai8_3_destruct_d;
  logic vai8_3_destruct_r;
  MyDTInt_Bool_t is_z_mapai9_3_destruct_d;
  logic is_z_mapai9_3_destruct_r;
  MyDTInt_Int_t f_mapaia_3_destruct_d;
  logic f_mapaia_3_destruct_r;
  Pointer_QTree_Int_t q2aid_2_destruct_d;
  logic q2aid_2_destruct_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_7_destruct_d;
  logic sc_0_7_destruct_r;
  Pointer_QTree_Int_t q1aic_1_destruct_d;
  logic q1aic_1_destruct_r;
  MyDTInt_Bool_t is_z_kronai6_2_destruct_d;
  logic is_z_kronai6_2_destruct_r;
  MyDTInt_Int_Int_t op_kronai7_2_destruct_d;
  logic op_kronai7_2_destruct_r;
  Int_t vai8_2_destruct_d;
  logic vai8_2_destruct_r;
  MyDTInt_Bool_t is_z_mapai9_2_destruct_d;
  logic is_z_mapai9_2_destruct_r;
  MyDTInt_Int_t f_mapaia_2_destruct_d;
  logic f_mapaia_2_destruct_r;
  Pointer_QTree_Int_t q2aid_1_destruct_d;
  logic q2aid_1_destruct_r;
  Pointer_QTree_Int_t q3aie_1_destruct_d;
  logic q3aie_1_destruct_r;
  \CTf'_f'_Int_Int_Int_Int_t  _18_d;
  logic _18_r;
  assign _18_r = 1'd1;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d ;
  logic \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_r ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d ;
  logic \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_r ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d ;
  logic \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_r ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d ;
  logic \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_r ;
  Go_t _17_d;
  logic _17_r;
  assign _17_r = 1'd1;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_r ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d ;
  logic \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_r ;
  QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r ;
  QTree_Int_t lizzieLet27_1_argbuf_d;
  logic lizzieLet27_1_argbuf_r;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet26_1_argbuf_d;
  logic lizzieLet26_1_argbuf_r;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet25_1_argbuf_d;
  logic lizzieLet25_1_argbuf_r;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet24_1_argbuf_d;
  logic lizzieLet24_1_argbuf_r;
  Pointer_QTree_Int_t \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d ;
  logic \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r ;
  Pointer_QTree_Int_t \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  logic \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r ;
  Go_t \call_f'_f'_Int_Int_Int_Int_goConst_d ;
  logic \call_f'_f'_Int_Int_Int_Int_goConst_r ;
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_Int_resbuf_d ;
  logic \f'_f'_Int_Int_Int_Int_resbuf_r ;
  Pointer_QTree_Int_t es_1_1_destruct_d;
  logic es_1_1_destruct_r;
  Pointer_QTree_Int_t es_2_2_destruct_d;
  logic es_2_2_destruct_r;
  Pointer_QTree_Int_t es_3_3_destruct_d;
  logic es_3_3_destruct_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_14_destruct_d;
  logic sc_0_14_destruct_r;
  Pointer_QTree_Int_t es_2_1_destruct_d;
  logic es_2_1_destruct_r;
  Pointer_QTree_Int_t es_3_2_destruct_d;
  logic es_3_2_destruct_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_13_destruct_d;
  logic sc_0_13_destruct_r;
  Pointer_QTree_Int_t q1ai1_3_destruct_d;
  logic q1ai1_3_destruct_r;
  Pointer_QTree_Int_t m2ahV_4_destruct_d;
  logic m2ahV_4_destruct_r;
  MyDTInt_Bool_t is_z_kronahW_4_destruct_d;
  logic is_z_kronahW_4_destruct_r;
  MyDTInt_Int_Int_t op_kronahX_4_destruct_d;
  logic op_kronahX_4_destruct_r;
  MyDTInt_Bool_t is_z_mapahY_4_destruct_d;
  logic is_z_mapahY_4_destruct_r;
  MyDTInt_Int_t f_mapahZ_4_destruct_d;
  logic f_mapahZ_4_destruct_r;
  Pointer_QTree_Int_t es_3_1_destruct_d;
  logic es_3_1_destruct_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_12_destruct_d;
  logic sc_0_12_destruct_r;
  Pointer_QTree_Int_t q1ai1_2_destruct_d;
  logic q1ai1_2_destruct_r;
  Pointer_QTree_Int_t m2ahV_3_destruct_d;
  logic m2ahV_3_destruct_r;
  MyDTInt_Bool_t is_z_kronahW_3_destruct_d;
  logic is_z_kronahW_3_destruct_r;
  MyDTInt_Int_Int_t op_kronahX_3_destruct_d;
  logic op_kronahX_3_destruct_r;
  MyDTInt_Bool_t is_z_mapahY_3_destruct_d;
  logic is_z_mapahY_3_destruct_r;
  MyDTInt_Int_t f_mapahZ_3_destruct_d;
  logic f_mapahZ_3_destruct_r;
  Pointer_QTree_Int_t q2ai2_2_destruct_d;
  logic q2ai2_2_destruct_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_11_destruct_d;
  logic sc_0_11_destruct_r;
  Pointer_QTree_Int_t q1ai1_1_destruct_d;
  logic q1ai1_1_destruct_r;
  Pointer_QTree_Int_t m2ahV_2_destruct_d;
  logic m2ahV_2_destruct_r;
  MyDTInt_Bool_t is_z_kronahW_2_destruct_d;
  logic is_z_kronahW_2_destruct_r;
  MyDTInt_Int_Int_t op_kronahX_2_destruct_d;
  logic op_kronahX_2_destruct_r;
  MyDTInt_Bool_t is_z_mapahY_2_destruct_d;
  logic is_z_mapahY_2_destruct_r;
  MyDTInt_Int_t f_mapahZ_2_destruct_d;
  logic f_mapahZ_2_destruct_r;
  Pointer_QTree_Int_t q2ai2_1_destruct_d;
  logic q2ai2_1_destruct_r;
  Pointer_QTree_Int_t q3ai3_1_destruct_d;
  logic q3ai3_1_destruct_r;
  CTf_f_Int_Int_Int_Int_t _16_d;
  logic _16_r;
  assign _16_r = 1'd1;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d;
  logic lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d;
  logic lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d;
  logic lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d;
  logic lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_r;
  Go_t _15_d;
  logic _15_r;
  assign _15_r = 1'd1;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_r;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d;
  logic lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_r;
  Pointer_QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_r;
  Pointer_QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_r;
  Pointer_QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_r;
  Pointer_QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_r;
  QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r;
  QTree_Int_t lizzieLet32_1_argbuf_d;
  logic lizzieLet32_1_argbuf_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet31_1_argbuf_d;
  logic lizzieLet31_1_argbuf_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet30_1_argbuf_d;
  logic lizzieLet30_1_argbuf_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet29_1_argbuf_d;
  logic lizzieLet29_1_argbuf_r;
  Pointer_QTree_Int_t lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d;
  logic lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r;
  Pointer_QTree_Int_t lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  logic lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r;
  Go_t call_f_f_Int_Int_Int_Int_goConst_d;
  logic call_f_f_Int_Int_Int_Int_goConst_r;
  Pointer_QTree_Int_t f_f_Int_Int_Int_Int_resbuf_d;
  logic f_f_Int_Int_Int_Int_resbuf_r;
  Go_t lizzieLet3_1MyFalse_d;
  logic lizzieLet3_1MyFalse_r;
  Go_t lizzieLet3_1MyTrue_d;
  logic lizzieLet3_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalse_d;
  logic lizzieLet3_1MyFalse_1MyFalse_r;
  MyBool_t lizzieLet3_1MyTrue_1MyTrue_d;
  logic lizzieLet3_1MyTrue_1MyTrue_r;
  MyBool_t lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d;
  logic lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r;
  Pointer_QTree_Int_t q1abW_destruct_d;
  logic q1abW_destruct_r;
  Pointer_QTree_Int_t q2abX_destruct_d;
  logic q2abX_destruct_r;
  Pointer_QTree_Int_t q3abY_destruct_d;
  logic q3abY_destruct_r;
  Pointer_QTree_Int_t q4abZ_destruct_d;
  logic q4abZ_destruct_r;
  QTree_Int_t _14_d;
  logic _14_r;
  assign _14_r = 1'd1;
  QTree_Int_t _13_d;
  logic _13_r;
  assign _13_r = 1'd1;
  QTree_Int_t lizzieLet4_1QNode_Int_d;
  logic lizzieLet4_1QNode_Int_r;
  QTree_Int_t _12_d;
  logic _12_r;
  assign _12_r = 1'd1;
  Go_t lizzieLet4_3QNone_Int_d;
  logic lizzieLet4_3QNone_Int_r;
  Go_t lizzieLet4_3QVal_Int_d;
  logic lizzieLet4_3QVal_Int_r;
  Go_t lizzieLet4_3QNode_Int_d;
  logic lizzieLet4_3QNode_Int_r;
  Go_t lizzieLet4_3QError_Int_d;
  logic lizzieLet4_3QError_Int_r;
  Go_t lizzieLet4_3QError_Int_1_d;
  logic lizzieLet4_3QError_Int_1_r;
  Go_t lizzieLet4_3QError_Int_2_d;
  logic lizzieLet4_3QError_Int_2_r;
  Go_t lizzieLet4_3QError_Int_1_argbuf_d;
  logic lizzieLet4_3QError_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet11_1_1_argbuf_d;
  logic lizzieLet11_1_1_argbuf_r;
  Go_t lizzieLet4_3QError_Int_2_argbuf_d;
  logic lizzieLet4_3QError_Int_2_argbuf_r;
  Go_t lizzieLet4_3QNode_Int_1_argbuf_d;
  logic lizzieLet4_3QNode_Int_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_1_d;
  logic lizzieLet4_3QNone_Int_1_r;
  Go_t lizzieLet4_3QNone_Int_2_d;
  logic lizzieLet4_3QNone_Int_2_r;
  Go_t lizzieLet4_3QNone_Int_1_argbuf_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_r;
  \Int#_t  lizzieLet11_1_argbuf_d;
  logic lizzieLet11_1_argbuf_r;
  Go_t lizzieLet4_3QNone_Int_2_argbuf_d;
  logic lizzieLet4_3QNone_Int_2_argbuf_r;
  C4_t go_15_goMux_choice_d;
  logic go_15_goMux_choice_r;
  Go_t go_15_goMux_data_d;
  logic go_15_goMux_data_r;
  Go_t lizzieLet4_3QVal_Int_1_d;
  logic lizzieLet4_3QVal_Int_1_r;
  Go_t lizzieLet4_3QVal_Int_2_d;
  logic lizzieLet4_3QVal_Int_2_r;
  Go_t lizzieLet4_3QVal_Int_1_argbuf_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_r;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_r;
  \Int#_t  lizzieLet12_1_argbuf_d;
  logic lizzieLet12_1_argbuf_r;
  Go_t lizzieLet4_3QVal_Int_2_argbuf_d;
  logic lizzieLet4_3QVal_Int_2_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_d;
  logic lizzieLet4_4QNone_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_d;
  logic lizzieLet4_4QVal_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNode_Int_d;
  logic lizzieLet4_4QNode_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_d;
  logic lizzieLet4_4QError_Int_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_1_argbuf_d;
  logic lizzieLet4_4QError_Int_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_d;
  logic lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_r;
  CT$wnnz_Int_t lizzieLet5_1_argbuf_d;
  logic lizzieLet5_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_1_argbuf_d;
  logic lizzieLet4_4QNone_Int_1_argbuf_r;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_1_argbuf_d;
  logic lizzieLet4_4QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t q1aic_destruct_d;
  logic q1aic_destruct_r;
  Pointer_QTree_Int_t q2aid_destruct_d;
  logic q2aid_destruct_r;
  Pointer_QTree_Int_t q3aie_destruct_d;
  logic q3aie_destruct_r;
  Pointer_QTree_Int_t q4aif_destruct_d;
  logic q4aif_destruct_r;
  Int_t \v'aib_destruct_d ;
  logic \v'aib_destruct_r ;
  QTree_Int_t _11_d;
  logic _11_r;
  assign _11_r = 1'd1;
  QTree_Int_t lizzieLet6_1QVal_Int_d;
  logic lizzieLet6_1QVal_Int_r;
  QTree_Int_t lizzieLet6_1QNode_Int_d;
  logic lizzieLet6_1QNode_Int_r;
  QTree_Int_t _10_d;
  logic _10_r;
  assign _10_r = 1'd1;
  MyDTInt_Int_t _9_d;
  logic _9_r;
  assign _9_r = 1'd1;
  MyDTInt_Int_t lizzieLet6_3QVal_Int_d;
  logic lizzieLet6_3QVal_Int_r;
  MyDTInt_Int_t lizzieLet6_3QNode_Int_d;
  logic lizzieLet6_3QNode_Int_r;
  MyDTInt_Int_t _8_d;
  logic _8_r;
  assign _8_r = 1'd1;
  MyDTInt_Int_t lizzieLet6_3QNode_Int_1_d;
  logic lizzieLet6_3QNode_Int_1_r;
  MyDTInt_Int_t lizzieLet6_3QNode_Int_2_d;
  logic lizzieLet6_3QNode_Int_2_r;
  MyDTInt_Int_t lizzieLet6_3QNode_Int_2_argbuf_d;
  logic lizzieLet6_3QNode_Int_2_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_d;
  logic lizzieLet6_4QNone_Int_r;
  Go_t lizzieLet6_4QVal_Int_d;
  logic lizzieLet6_4QVal_Int_r;
  Go_t lizzieLet6_4QNode_Int_d;
  logic lizzieLet6_4QNode_Int_r;
  Go_t lizzieLet6_4QError_Int_d;
  logic lizzieLet6_4QError_Int_r;
  Go_t lizzieLet6_4QError_Int_1_d;
  logic lizzieLet6_4QError_Int_1_r;
  Go_t lizzieLet6_4QError_Int_2_d;
  logic lizzieLet6_4QError_Int_2_r;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_d;
  logic lizzieLet6_4QError_Int_1QError_Int_r;
  QTree_Int_t lizzieLet12_1_1_argbuf_d;
  logic lizzieLet12_1_1_argbuf_r;
  Go_t lizzieLet6_4QError_Int_2_argbuf_d;
  logic lizzieLet6_4QError_Int_2_argbuf_r;
  Go_t lizzieLet6_4QNode_Int_1_argbuf_d;
  logic lizzieLet6_4QNode_Int_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_1_d;
  logic lizzieLet6_4QNone_Int_1_r;
  Go_t lizzieLet6_4QNone_Int_2_d;
  logic lizzieLet6_4QNone_Int_2_r;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_r;
  QTree_Int_t lizzieLet7_1_argbuf_d;
  logic lizzieLet7_1_argbuf_r;
  Go_t lizzieLet6_4QNone_Int_2_argbuf_d;
  logic lizzieLet6_4QNone_Int_2_argbuf_r;
  C6_t go_16_goMux_choice_d;
  logic go_16_goMux_choice_r;
  Go_t go_16_goMux_data_d;
  logic go_16_goMux_data_r;
  Go_t lizzieLet6_4QVal_Int_1_d;
  logic lizzieLet6_4QVal_Int_1_r;
  Go_t lizzieLet6_4QVal_Int_2_d;
  logic lizzieLet6_4QVal_Int_2_r;
  Go_t lizzieLet6_4QVal_Int_1_argbuf_d;
  logic lizzieLet6_4QVal_Int_1_argbuf_r;
  TupGo___MyDTInt_Bool___Int_t applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d;
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r;
  MyDTInt_Bool_t _7_d;
  logic _7_r;
  assign _7_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_d;
  logic lizzieLet6_5QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_d;
  logic lizzieLet6_5QNode_Int_r;
  MyDTInt_Bool_t _6_d;
  logic _6_r;
  assign _6_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_1_d;
  logic lizzieLet6_5QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_d;
  logic lizzieLet6_5QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_argbuf_d;
  logic lizzieLet6_5QNode_Int_2_argbuf_r;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_1_argbuf_d;
  logic lizzieLet6_5QVal_Int_1_argbuf_r;
  MyDTInt_Bool_t _5_d;
  logic _5_r;
  assign _5_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_6QVal_Int_d;
  logic lizzieLet6_6QVal_Int_r;
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_d;
  logic lizzieLet6_6QNode_Int_r;
  MyDTInt_Bool_t _4_d;
  logic _4_r;
  assign _4_r = 1'd1;
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_1_d;
  logic lizzieLet6_6QNode_Int_1_r;
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_2_d;
  logic lizzieLet6_6QNode_Int_2_r;
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_2_argbuf_d;
  logic lizzieLet6_6QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t _3_d;
  logic _3_r;
  assign _3_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_d;
  logic lizzieLet6_7QVal_Int_r;
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_d;
  logic lizzieLet6_7QNode_Int_r;
  MyDTInt_Int_Int_t _2_d;
  logic _2_r;
  assign _2_r = 1'd1;
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_1_d;
  logic lizzieLet6_7QNode_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_2_d;
  logic lizzieLet6_7QNode_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_2_argbuf_d;
  logic lizzieLet6_7QNode_Int_2_argbuf_r;
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_1_d;
  logic lizzieLet6_7QVal_Int_1_r;
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_2_d;
  logic lizzieLet6_7QVal_Int_2_r;
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_1_argbuf_d;
  logic lizzieLet6_7QVal_Int_1_argbuf_r;
  TupMyDTInt_Int_Int___Int___Int_t applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d;
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QNone_Int_d;
  logic lizzieLet6_8QNone_Int_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QVal_Int_d;
  logic lizzieLet6_8QVal_Int_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QNode_Int_d;
  logic lizzieLet6_8QNode_Int_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QError_Int_d;
  logic lizzieLet6_8QError_Int_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QError_Int_1_argbuf_d;
  logic lizzieLet6_8QError_Int_1_argbuf_r;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_d ;
  logic \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet11_2_1_argbuf_d;
  logic lizzieLet11_2_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QNone_Int_1_argbuf_d;
  logic lizzieLet6_8QNone_Int_1_argbuf_r;
  Int_t _1_d;
  logic _1_r;
  assign _1_r = 1'd1;
  Int_t lizzieLet6_9QVal_Int_d;
  logic lizzieLet6_9QVal_Int_r;
  Int_t lizzieLet6_9QNode_Int_d;
  logic lizzieLet6_9QNode_Int_r;
  Int_t _0_d;
  logic _0_r;
  assign _0_r = 1'd1;
  Int_t lizzieLet6_9QNode_Int_1_d;
  logic lizzieLet6_9QNode_Int_1_r;
  Int_t lizzieLet6_9QNode_Int_2_d;
  logic lizzieLet6_9QNode_Int_2_r;
  Int_t lizzieLet6_9QNode_Int_2_argbuf_d;
  logic lizzieLet6_9QNode_Int_2_argbuf_r;
  Int_t lizzieLet6_9QVal_Int_1_d;
  logic lizzieLet6_9QVal_Int_1_r;
  Int_t lizzieLet6_9QVal_Int_2_d;
  logic lizzieLet6_9QVal_Int_2_r;
  Int_t lizzieLet6_9QVal_Int_1_argbuf_d;
  logic lizzieLet6_9QVal_Int_1_argbuf_r;
  Pointer_QTree_Int_t m1ahU_1_argbuf_d;
  logic m1ahU_1_argbuf_r;
  Pointer_QTree_Int_t m2ahV_2_2_argbuf_d;
  logic m2ahV_2_2_argbuf_r;
  Pointer_QTree_Int_t m2ahV_2_1_d;
  logic m2ahV_2_1_r;
  Pointer_QTree_Int_t m2ahV_2_2_d;
  logic m2ahV_2_2_r;
  Pointer_QTree_Int_t m2ahV_3_2_argbuf_d;
  logic m2ahV_3_2_argbuf_r;
  Pointer_QTree_Int_t m2ahV_3_1_d;
  logic m2ahV_3_1_r;
  Pointer_QTree_Int_t m2ahV_3_2_d;
  logic m2ahV_3_2_r;
  Pointer_QTree_Int_t m2ahV_4_1_argbuf_d;
  logic m2ahV_4_1_argbuf_r;
  Pointer_QTree_Int_t m2ai5_1_argbuf_d;
  logic m2ai5_1_argbuf_r;
  MyDTInt_Int_Int_t op_kronahX_2_2_argbuf_d;
  logic op_kronahX_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_kronahX_2_1_d;
  logic op_kronahX_2_1_r;
  MyDTInt_Int_Int_t op_kronahX_2_2_d;
  logic op_kronahX_2_2_r;
  MyDTInt_Int_Int_t op_kronahX_3_2_argbuf_d;
  logic op_kronahX_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_kronahX_3_1_d;
  logic op_kronahX_3_1_r;
  MyDTInt_Int_Int_t op_kronahX_3_2_d;
  logic op_kronahX_3_2_r;
  MyDTInt_Int_Int_t op_kronahX_4_1_argbuf_d;
  logic op_kronahX_4_1_argbuf_r;
  MyDTInt_Int_Int_t op_kronai7_2_2_argbuf_d;
  logic op_kronai7_2_2_argbuf_r;
  MyDTInt_Int_Int_t op_kronai7_2_1_d;
  logic op_kronai7_2_1_r;
  MyDTInt_Int_Int_t op_kronai7_2_2_d;
  logic op_kronai7_2_2_r;
  MyDTInt_Int_Int_t op_kronai7_3_2_argbuf_d;
  logic op_kronai7_3_2_argbuf_r;
  MyDTInt_Int_Int_t op_kronai7_3_1_d;
  logic op_kronai7_3_1_r;
  MyDTInt_Int_Int_t op_kronai7_3_2_d;
  logic op_kronai7_3_2_r;
  MyDTInt_Int_Int_t op_kronai7_4_1_argbuf_d;
  logic op_kronai7_4_1_argbuf_r;
  Pointer_QTree_Int_t q1abW_1_argbuf_d;
  logic q1abW_1_argbuf_r;
  Pointer_QTree_Int_t q1ai1_3_1_argbuf_d;
  logic q1ai1_3_1_argbuf_r;
  Pointer_QTree_Int_t q1aic_3_1_argbuf_d;
  logic q1aic_3_1_argbuf_r;
  Pointer_QTree_Int_t q2abX_1_1_argbuf_d;
  logic q2abX_1_1_argbuf_r;
  Pointer_QTree_Int_t q2ai2_2_1_argbuf_d;
  logic q2ai2_2_1_argbuf_r;
  Pointer_QTree_Int_t q2aid_2_1_argbuf_d;
  logic q2aid_2_1_argbuf_r;
  Pointer_QTree_Int_t q3abY_2_1_argbuf_d;
  logic q3abY_2_1_argbuf_r;
  Pointer_QTree_Int_t q3ai3_1_1_argbuf_d;
  logic q3ai3_1_1_argbuf_r;
  Pointer_QTree_Int_t q3aie_1_1_argbuf_d;
  logic q3aie_1_1_argbuf_r;
  Pointer_QTree_Int_t q4abZ_3_1_argbuf_d;
  logic q4abZ_3_1_argbuf_r;
  Pointer_QTree_Int_t q4ai4_1_argbuf_d;
  logic q4ai4_1_argbuf_r;
  Pointer_QTree_Int_t q4aif_1_argbuf_d;
  logic q4aif_1_argbuf_r;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r;
  CT$wnnz_Int_t lizzieLet19_1_d;
  logic lizzieLet19_1_r;
  CT$wnnz_Int_t lizzieLet19_2_d;
  logic lizzieLet19_2_r;
  CT$wnnz_Int_t lizzieLet19_3_d;
  logic lizzieLet19_3_r;
  CT$wnnz_Int_t lizzieLet19_4_d;
  logic lizzieLet19_4_r;
  \CTf'_f'_Int_Int_Int_Int_t  \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d ;
  logic \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r ;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet23_1_d;
  logic lizzieLet23_1_r;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet23_2_d;
  logic lizzieLet23_2_r;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet23_3_d;
  logic lizzieLet23_3_r;
  \CTf'_f'_Int_Int_Int_Int_t  lizzieLet23_4_d;
  logic lizzieLet23_4_r;
  CTf_f_Int_Int_Int_Int_t readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d;
  logic readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_1_d;
  logic lizzieLet28_1_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_2_d;
  logic lizzieLet28_2_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_3_d;
  logic lizzieLet28_3_r;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4_d;
  logic lizzieLet28_4_r;
  QTree_Int_t readPointer_QTree_Intm1ahU_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm1ahU_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet13_1_1_d;
  logic lizzieLet13_1_1_r;
  QTree_Int_t lizzieLet13_1_2_d;
  logic lizzieLet13_1_2_r;
  QTree_Int_t lizzieLet13_1_3_d;
  logic lizzieLet13_1_3_r;
  QTree_Int_t lizzieLet13_1_4_d;
  logic lizzieLet13_1_4_r;
  QTree_Int_t lizzieLet13_1_5_d;
  logic lizzieLet13_1_5_r;
  QTree_Int_t lizzieLet13_1_6_d;
  logic lizzieLet13_1_6_r;
  QTree_Int_t lizzieLet13_1_7_d;
  logic lizzieLet13_1_7_r;
  QTree_Int_t lizzieLet13_1_8_d;
  logic lizzieLet13_1_8_r;
  QTree_Int_t lizzieLet13_1_9_d;
  logic lizzieLet13_1_9_r;
  QTree_Int_t readPointer_QTree_Intm2ai5_1_argbuf_rwb_d;
  logic readPointer_QTree_Intm2ai5_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet6_1_d;
  logic lizzieLet6_1_r;
  QTree_Int_t lizzieLet6_2_d;
  logic lizzieLet6_2_r;
  QTree_Int_t lizzieLet6_3_d;
  logic lizzieLet6_3_r;
  QTree_Int_t lizzieLet6_4_d;
  logic lizzieLet6_4_r;
  QTree_Int_t lizzieLet6_5_d;
  logic lizzieLet6_5_r;
  QTree_Int_t lizzieLet6_6_d;
  logic lizzieLet6_6_r;
  QTree_Int_t lizzieLet6_7_d;
  logic lizzieLet6_7_r;
  QTree_Int_t lizzieLet6_8_d;
  logic lizzieLet6_8_r;
  QTree_Int_t lizzieLet6_9_d;
  logic lizzieLet6_9_r;
  QTree_Int_t readPointer_QTree_IntwstH_1_1_argbuf_rwb_d;
  logic readPointer_QTree_IntwstH_1_1_argbuf_rwb_r;
  QTree_Int_t lizzieLet4_1_d;
  logic lizzieLet4_1_r;
  QTree_Int_t lizzieLet4_2_d;
  logic lizzieLet4_2_r;
  QTree_Int_t lizzieLet4_3_d;
  logic lizzieLet4_3_r;
  QTree_Int_t lizzieLet4_4_d;
  logic lizzieLet4_4_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_10_1_argbuf_d;
  logic sc_0_10_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_14_1_argbuf_d;
  logic sc_0_14_1_argbuf_r;
  Pointer_CT$wnnz_Int_t sc_0_6_1_argbuf_d;
  logic sc_0_6_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  scfarg_0_1_1_argbuf_d;
  logic scfarg_0_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t scfarg_0_2_1_argbuf_d;
  logic scfarg_0_2_1_argbuf_r;
  Pointer_CT$wnnz_Int_t scfarg_0_1_argbuf_d;
  logic scfarg_0_1_argbuf_r;
  Int_t \v'aib_1_argbuf_d ;
  logic \v'aib_1_argbuf_r ;
  Int_t \v'aib_1_d ;
  logic \v'aib_1_r ;
  Int_t \v'aib_2_d ;
  logic \v'aib_2_r ;
  Int_t vai0_1_argbuf_d;
  logic vai0_1_argbuf_r;
  Int_t vai8_2_2_argbuf_d;
  logic vai8_2_2_argbuf_r;
  Int_t vai8_2_1_d;
  logic vai8_2_1_r;
  Int_t vai8_2_2_d;
  logic vai8_2_2_r;
  Int_t vai8_3_2_argbuf_d;
  logic vai8_3_2_argbuf_r;
  Int_t vai8_3_1_d;
  logic vai8_3_1_r;
  Int_t vai8_3_2_d;
  logic vai8_3_2_r;
  Int_t vai8_4_1_argbuf_d;
  logic vai8_4_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t lizzieLet13_1_argbuf_d;
  logic lizzieLet13_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca2_1_argbuf_d;
  logic sca2_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca1_1_argbuf_d;
  logic sca1_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca0_1_argbuf_d;
  logic sca0_1_argbuf_r;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r;
  Pointer_CT$wnnz_Int_t sca3_1_argbuf_d;
  logic sca3_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sca3_1_1_argbuf_d;
  logic sca3_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_1_1_argbuf_d;
  logic lizzieLet6_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sca2_1_1_argbuf_d;
  logic sca2_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sca1_1_1_argbuf_d;
  logic sca1_1_1_argbuf_r;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_r ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sca0_1_1_argbuf_d;
  logic sca0_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sca3_2_1_argbuf_d;
  logic sca3_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet10_1_1_argbuf_d;
  logic lizzieLet10_1_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sca2_2_1_argbuf_d;
  logic sca2_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sca1_2_1_argbuf_d;
  logic sca1_2_1_argbuf_r;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_r;
  Pointer_CTf_f_Int_Int_Int_Int_t sca0_2_1_argbuf_d;
  logic sca0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet4_1_1_argbuf_d;
  logic lizzieLet4_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet5_1_1_argbuf_d;
  logic lizzieLet5_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet7_1_1_argbuf_d;
  logic lizzieLet7_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet9_1_1_argbuf_d;
  logic lizzieLet9_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_1_1_argbuf_d;
  logic contRet_0_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_r;
  Pointer_QTree_Int_t contRet_0_2_1_argbuf_d;
  logic contRet_0_2_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet1_1_1_argbuf_d;
  logic lizzieLet1_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet2_1_1_argbuf_d;
  logic lizzieLet2_1_1_argbuf_r;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_r;
  Pointer_QTree_Int_t lizzieLet3_1_1_argbuf_d;
  logic lizzieLet3_1_1_argbuf_r;
  Pointer_QTree_Int_t wstH_1_1_argbuf_d;
  logic wstH_1_1_argbuf_r;
  CT$wnnz_Int_t lizzieLet21_1_argbuf_d;
  logic lizzieLet21_1_argbuf_r;
  CT$wnnz_Int_t wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_d;
  logic wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_r;
  CT$wnnz_Int_t lizzieLet22_1_argbuf_d;
  logic lizzieLet22_1_argbuf_r;
  CT$wnnz_Int_t wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_d;
  logic wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_r;
  \Int#_t  es_6_2_1ww2XuO_1_1_Add32_d;
  logic es_6_2_1ww2XuO_1_1_Add32_r;
  \Int#_t  wwstK_4_1ww1XuL_2_1_Add32_d;
  logic wwstK_4_1ww1XuL_2_1_Add32_r;
  Int_t \es_0_1_1I#_d ;
  logic \es_0_1_1I#_r ;
  \Int#_t  xap7_1lizzieLet0_1_1_Add32_d;
  logic xap7_1lizzieLet0_1_1_Add32_r;
  
  /* fork (Ty Go) : (sourceGo,Go) > [(go_1,Go),
                                (go_2,Go),
                                (go_3,Go),
                                (go_4,Go),
                                (go_5,Go),
                                (go_6,Go),
                                (go__7,Go),
                                (go__8,Go),
                                (go__9,Go),
                                (go__10,Go),
                                (go__11,Go),
                                (go__12,Go)] */
  logic [11:0] sourceGo_emitted;
  logic [11:0] sourceGo_done;
  assign go_1_d = (sourceGo_d[0] && (! sourceGo_emitted[0]));
  assign go_2_d = (sourceGo_d[0] && (! sourceGo_emitted[1]));
  assign go_3_d = (sourceGo_d[0] && (! sourceGo_emitted[2]));
  assign go_4_d = (sourceGo_d[0] && (! sourceGo_emitted[3]));
  assign go_5_d = (sourceGo_d[0] && (! sourceGo_emitted[4]));
  assign go_6_d = (sourceGo_d[0] && (! sourceGo_emitted[5]));
  assign go__7_d = (sourceGo_d[0] && (! sourceGo_emitted[6]));
  assign go__8_d = (sourceGo_d[0] && (! sourceGo_emitted[7]));
  assign go__9_d = (sourceGo_d[0] && (! sourceGo_emitted[8]));
  assign go__10_d = (sourceGo_d[0] && (! sourceGo_emitted[9]));
  assign go__11_d = (sourceGo_d[0] && (! sourceGo_emitted[10]));
  assign go__12_d = (sourceGo_d[0] && (! sourceGo_emitted[11]));
  assign sourceGo_done = (sourceGo_emitted | ({go__12_d[0],
                                               go__11_d[0],
                                               go__10_d[0],
                                               go__9_d[0],
                                               go__8_d[0],
                                               go__7_d[0],
                                               go_6_d[0],
                                               go_5_d[0],
                                               go_4_d[0],
                                               go_3_d[0],
                                               go_2_d[0],
                                               go_1_d[0]} & {go__12_r,
                                                             go__11_r,
                                                             go__10_r,
                                                             go__9_r,
                                                             go__8_r,
                                                             go__7_r,
                                                             go_6_r,
                                                             go_5_r,
                                                             go_4_r,
                                                             go_3_r,
                                                             go_2_r,
                                                             go_1_r}));
  assign sourceGo_r = (& sourceGo_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sourceGo_emitted <= 12'd0;
    else
      sourceGo_emitted <= (sourceGo_r ? 12'd0 :
                           sourceGo_done);
  
  /* const (Ty Word16#,
       Lit 0) : (go__7,Go) > (initHP_CT$wnnz_Int,Word16#) */
  assign initHP_CT$wnnz_Int_d = {16'd0, go__7_d[0]};
  assign go__7_r = initHP_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CT$wnnz_Int1,Go) > (incrHP_CT$wnnz_Int,Word16#) */
  assign incrHP_CT$wnnz_Int_d = {16'd1, incrHP_CT$wnnz_Int1_d[0]};
  assign incrHP_CT$wnnz_Int1_r = incrHP_CT$wnnz_Int_r;
  
  /* merge (Ty Go) : [(go__8,Go),
                 (incrHP_CT$wnnz_Int2,Go)] > (incrHP_mergeCT$wnnz_Int,Go) */
  logic [1:0] incrHP_mergeCT$wnnz_Int_selected;
  logic [1:0] incrHP_mergeCT$wnnz_Int_select;
  always_comb
    begin
      incrHP_mergeCT$wnnz_Int_selected = 2'd0;
      if ((| incrHP_mergeCT$wnnz_Int_select))
        incrHP_mergeCT$wnnz_Int_selected = incrHP_mergeCT$wnnz_Int_select;
      else
        if (go__8_d[0]) incrHP_mergeCT$wnnz_Int_selected[0] = 1'd1;
        else if (incrHP_CT$wnnz_Int2_d[0])
          incrHP_mergeCT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_select <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_select <= (incrHP_mergeCT$wnnz_Int_r ? 2'd0 :
                                         incrHP_mergeCT$wnnz_Int_selected);
  always_comb
    if (incrHP_mergeCT$wnnz_Int_selected[0])
      incrHP_mergeCT$wnnz_Int_d = go__8_d;
    else if (incrHP_mergeCT$wnnz_Int_selected[1])
      incrHP_mergeCT$wnnz_Int_d = incrHP_CT$wnnz_Int2_d;
    else incrHP_mergeCT$wnnz_Int_d = 1'd0;
  assign {incrHP_CT$wnnz_Int2_r,
          go__8_r} = (incrHP_mergeCT$wnnz_Int_r ? incrHP_mergeCT$wnnz_Int_selected :
                      2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCT$wnnz_Int_buf,Go) > [(incrHP_CT$wnnz_Int1,Go),
                                                   (incrHP_CT$wnnz_Int2,Go)] */
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_emitted;
  logic [1:0] incrHP_mergeCT$wnnz_Int_buf_done;
  assign incrHP_CT$wnnz_Int1_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[0]));
  assign incrHP_CT$wnnz_Int2_d = (incrHP_mergeCT$wnnz_Int_buf_d[0] && (! incrHP_mergeCT$wnnz_Int_buf_emitted[1]));
  assign incrHP_mergeCT$wnnz_Int_buf_done = (incrHP_mergeCT$wnnz_Int_buf_emitted | ({incrHP_CT$wnnz_Int2_d[0],
                                                                                     incrHP_CT$wnnz_Int1_d[0]} & {incrHP_CT$wnnz_Int2_r,
                                                                                                                  incrHP_CT$wnnz_Int1_r}));
  assign incrHP_mergeCT$wnnz_Int_buf_r = (& incrHP_mergeCT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCT$wnnz_Int_buf_emitted <= (incrHP_mergeCT$wnnz_Int_buf_r ? 2'd0 :
                                              incrHP_mergeCT$wnnz_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CT$wnnz_Int,Word16#) (forkHP1_CT$wnnz_Int,Word16#) > (addHP_CT$wnnz_Int,Word16#) */
  assign addHP_CT$wnnz_Int_d = {(incrHP_CT$wnnz_Int_d[16:1] + forkHP1_CT$wnnz_Int_d[16:1]),
                                (incrHP_CT$wnnz_Int_d[0] && forkHP1_CT$wnnz_Int_d[0])};
  assign {incrHP_CT$wnnz_Int_r,
          forkHP1_CT$wnnz_Int_r} = {2 {(addHP_CT$wnnz_Int_r && addHP_CT$wnnz_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CT$wnnz_Int,Word16#),
                      (addHP_CT$wnnz_Int,Word16#)] > (mergeHP_CT$wnnz_Int,Word16#) */
  logic [1:0] mergeHP_CT$wnnz_Int_selected;
  logic [1:0] mergeHP_CT$wnnz_Int_select;
  always_comb
    begin
      mergeHP_CT$wnnz_Int_selected = 2'd0;
      if ((| mergeHP_CT$wnnz_Int_select))
        mergeHP_CT$wnnz_Int_selected = mergeHP_CT$wnnz_Int_select;
      else
        if (initHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[0] = 1'd1;
        else if (addHP_CT$wnnz_Int_d[0])
          mergeHP_CT$wnnz_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_select <= 2'd0;
    else
      mergeHP_CT$wnnz_Int_select <= (mergeHP_CT$wnnz_Int_r ? 2'd0 :
                                     mergeHP_CT$wnnz_Int_selected);
  always_comb
    if (mergeHP_CT$wnnz_Int_selected[0])
      mergeHP_CT$wnnz_Int_d = initHP_CT$wnnz_Int_d;
    else if (mergeHP_CT$wnnz_Int_selected[1])
      mergeHP_CT$wnnz_Int_d = addHP_CT$wnnz_Int_d;
    else mergeHP_CT$wnnz_Int_d = {16'd0, 1'd0};
  assign {addHP_CT$wnnz_Int_r,
          initHP_CT$wnnz_Int_r} = (mergeHP_CT$wnnz_Int_r ? mergeHP_CT$wnnz_Int_selected :
                                   2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCT$wnnz_Int,Go) > (incrHP_mergeCT$wnnz_Int_buf,Go) */
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_d;
  logic incrHP_mergeCT$wnnz_Int_bufchan_r;
  assign incrHP_mergeCT$wnnz_Int_r = ((! incrHP_mergeCT$wnnz_Int_bufchan_d[0]) || incrHP_mergeCT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCT$wnnz_Int_r)
        incrHP_mergeCT$wnnz_Int_bufchan_d <= incrHP_mergeCT$wnnz_Int_d;
  Go_t incrHP_mergeCT$wnnz_Int_bufchan_buf;
  assign incrHP_mergeCT$wnnz_Int_bufchan_r = (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0]);
  assign incrHP_mergeCT$wnnz_Int_buf_d = (incrHP_mergeCT$wnnz_Int_bufchan_buf[0] ? incrHP_mergeCT$wnnz_Int_bufchan_buf :
                                          incrHP_mergeCT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCT$wnnz_Int_buf_r && incrHP_mergeCT$wnnz_Int_bufchan_buf[0]))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCT$wnnz_Int_buf_r) && (! incrHP_mergeCT$wnnz_Int_bufchan_buf[0])))
        incrHP_mergeCT$wnnz_Int_bufchan_buf <= incrHP_mergeCT$wnnz_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CT$wnnz_Int,Word16#) > (mergeHP_CT$wnnz_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_d;
  logic mergeHP_CT$wnnz_Int_bufchan_r;
  assign mergeHP_CT$wnnz_Int_r = ((! mergeHP_CT$wnnz_Int_bufchan_d[0]) || mergeHP_CT$wnnz_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CT$wnnz_Int_r)
        mergeHP_CT$wnnz_Int_bufchan_d <= mergeHP_CT$wnnz_Int_d;
  \Word16#_t  mergeHP_CT$wnnz_Int_bufchan_buf;
  assign mergeHP_CT$wnnz_Int_bufchan_r = (! mergeHP_CT$wnnz_Int_bufchan_buf[0]);
  assign mergeHP_CT$wnnz_Int_buf_d = (mergeHP_CT$wnnz_Int_bufchan_buf[0] ? mergeHP_CT$wnnz_Int_bufchan_buf :
                                      mergeHP_CT$wnnz_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CT$wnnz_Int_buf_r && mergeHP_CT$wnnz_Int_bufchan_buf[0]))
        mergeHP_CT$wnnz_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CT$wnnz_Int_buf_r) && (! mergeHP_CT$wnnz_Int_bufchan_buf[0])))
        mergeHP_CT$wnnz_Int_bufchan_buf <= mergeHP_CT$wnnz_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CT$wnnz_Int_buf,Word16#) > [(forkHP1_CT$wnnz_Int,Word16#),
                                                         (forkHP1_CT$wnnz_In2,Word16#),
                                                         (forkHP1_CT$wnnz_In3,Word16#)] */
  logic [2:0] mergeHP_CT$wnnz_Int_buf_emitted;
  logic [2:0] mergeHP_CT$wnnz_Int_buf_done;
  assign forkHP1_CT$wnnz_Int_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[0]))};
  assign forkHP1_CT$wnnz_In2_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[1]))};
  assign forkHP1_CT$wnnz_In3_d = {mergeHP_CT$wnnz_Int_buf_d[16:1],
                                  (mergeHP_CT$wnnz_Int_buf_d[0] && (! mergeHP_CT$wnnz_Int_buf_emitted[2]))};
  assign mergeHP_CT$wnnz_Int_buf_done = (mergeHP_CT$wnnz_Int_buf_emitted | ({forkHP1_CT$wnnz_In3_d[0],
                                                                             forkHP1_CT$wnnz_In2_d[0],
                                                                             forkHP1_CT$wnnz_Int_d[0]} & {forkHP1_CT$wnnz_In3_r,
                                                                                                          forkHP1_CT$wnnz_In2_r,
                                                                                                          forkHP1_CT$wnnz_Int_r}));
  assign mergeHP_CT$wnnz_Int_buf_r = (& mergeHP_CT$wnnz_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CT$wnnz_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CT$wnnz_Int_buf_emitted <= (mergeHP_CT$wnnz_Int_buf_r ? 3'd0 :
                                          mergeHP_CT$wnnz_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CT$wnnz_Int) : [(dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int),
                                    (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int)] > (memMergeChoice_CT$wnnz_Int,C2) (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  logic [1:0] dconReadIn_CT$wnnz_Int_select_d;
  assign dconReadIn_CT$wnnz_Int_select_d = ((| dconReadIn_CT$wnnz_Int_select_q) ? dconReadIn_CT$wnnz_Int_select_q :
                                            (dconReadIn_CT$wnnz_Int_d[0] ? 2'd1 :
                                             (dconWriteIn_CT$wnnz_Int_d[0] ? 2'd2 :
                                              2'd0)));
  logic [1:0] dconReadIn_CT$wnnz_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_select_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_select_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                          dconReadIn_CT$wnnz_Int_select_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_CT$wnnz_Int_emit_q <= 2'd0;
    else
      dconReadIn_CT$wnnz_Int_emit_q <= (dconReadIn_CT$wnnz_Int_done ? 2'd0 :
                                        dconReadIn_CT$wnnz_Int_emit_d);
  logic [1:0] dconReadIn_CT$wnnz_Int_emit_d;
  assign dconReadIn_CT$wnnz_Int_emit_d = (dconReadIn_CT$wnnz_Int_emit_q | ({memMergeChoice_CT$wnnz_Int_d[0],
                                                                            memMergeIn_CT$wnnz_Int_d[0]} & {memMergeChoice_CT$wnnz_Int_r,
                                                                                                            memMergeIn_CT$wnnz_Int_r}));
  logic dconReadIn_CT$wnnz_Int_done;
  assign dconReadIn_CT$wnnz_Int_done = (& dconReadIn_CT$wnnz_Int_emit_d);
  assign {dconWriteIn_CT$wnnz_Int_r,
          dconReadIn_CT$wnnz_Int_r} = (dconReadIn_CT$wnnz_Int_done ? dconReadIn_CT$wnnz_Int_select_d :
                                       2'd0);
  assign memMergeIn_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconReadIn_CT$wnnz_Int_d :
                                     ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[0])) ? dconWriteIn_CT$wnnz_Int_d :
                                      {132'd0, 1'd0}));
  assign memMergeChoice_CT$wnnz_Int_d = ((dconReadIn_CT$wnnz_Int_select_d[0] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                         ((dconReadIn_CT$wnnz_Int_select_d[1] && (! dconReadIn_CT$wnnz_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                          {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CT$wnnz_Int,
      Ty MemOut_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) > (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) */
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CT$wnnz_Int_dbuf_address;
  logic [114:0] memMergeIn_CT$wnnz_Int_dbuf_din;
  logic [114:0] memOut_CT$wnnz_Int_q;
  logic memOut_CT$wnnz_Int_valid;
  logic memMergeIn_CT$wnnz_Int_dbuf_we;
  logic memOut_CT$wnnz_Int_we;
  assign memMergeIn_CT$wnnz_Int_dbuf_din = memMergeIn_CT$wnnz_Int_dbuf_d[132:18];
  assign memMergeIn_CT$wnnz_Int_dbuf_address = memMergeIn_CT$wnnz_Int_dbuf_d[17:2];
  assign memMergeIn_CT$wnnz_Int_dbuf_we = (memMergeIn_CT$wnnz_Int_dbuf_d[1:1] && memMergeIn_CT$wnnz_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CT$wnnz_Int_we <= 1'd0;
        memOut_CT$wnnz_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CT$wnnz_Int_we <= memMergeIn_CT$wnnz_Int_dbuf_we;
        memOut_CT$wnnz_Int_valid <= memMergeIn_CT$wnnz_Int_dbuf_d[0];
        if (memMergeIn_CT$wnnz_Int_dbuf_we)
          begin
            memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address] <= memMergeIn_CT$wnnz_Int_dbuf_din;
            memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_din;
          end
        else
          memOut_CT$wnnz_Int_q <= memMergeIn_CT$wnnz_Int_dbuf_mem[memMergeIn_CT$wnnz_Int_dbuf_address];
      end
  assign memOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_q,
                                 memOut_CT$wnnz_Int_we,
                                 memOut_CT$wnnz_Int_valid};
  assign memMergeIn_CT$wnnz_Int_dbuf_r = ((! memOut_CT$wnnz_Int_valid) || memOut_CT$wnnz_Int_r);
  logic [31:0] profiling_MemIn_CT$wnnz_Int_read;
  logic [31:0] profiling_MemIn_CT$wnnz_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CT$wnnz_Int_write <= 0;
        profiling_MemIn_CT$wnnz_Int_read <= 0;
      end
    else
      if ((memMergeIn_CT$wnnz_Int_dbuf_we == 1'd1))
        profiling_MemIn_CT$wnnz_Int_write <= (profiling_MemIn_CT$wnnz_Int_write + 1);
      else
        if ((memOut_CT$wnnz_Int_valid == 1'd1))
          profiling_MemIn_CT$wnnz_Int_read <= (profiling_MemIn_CT$wnnz_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CT$wnnz_Int) : (memMergeChoice_CT$wnnz_Int,C2) (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) > [(memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int),
                                                                                                                (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int)] */
  logic [1:0] memOut_CT$wnnz_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CT$wnnz_Int_d[0] && memOut_CT$wnnz_Int_dbuf_d[0]))
      unique case (memMergeChoice_CT$wnnz_Int_d[1:1])
        1'd0: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd2;
        default: memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CT$wnnz_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                     memOut_CT$wnnz_Int_dbuf_onehotd[0]};
  assign memWriteOut_CT$wnnz_Int_d = {memOut_CT$wnnz_Int_dbuf_d[116:1],
                                      memOut_CT$wnnz_Int_dbuf_onehotd[1]};
  assign memOut_CT$wnnz_Int_dbuf_r = (| (memOut_CT$wnnz_Int_dbuf_onehotd & {memWriteOut_CT$wnnz_Int_r,
                                                                            memReadOut_CT$wnnz_Int_r}));
  assign memMergeChoice_CT$wnnz_Int_r = memOut_CT$wnnz_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_dbuf,MemIn_CT$wnnz_Int) */
  assign memMergeIn_CT$wnnz_Int_rbuf_r = ((! memMergeIn_CT$wnnz_Int_dbuf_d[0]) || memMergeIn_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CT$wnnz_Int_dbuf_d <= {132'd0, 1'd0};
    else
      if (memMergeIn_CT$wnnz_Int_rbuf_r)
        memMergeIn_CT$wnnz_Int_dbuf_d <= memMergeIn_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CT$wnnz_Int) : (memMergeIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) > (memMergeIn_CT$wnnz_Int_rbuf,MemIn_CT$wnnz_Int) */
  MemIn_CT$wnnz_Int_t memMergeIn_CT$wnnz_Int_buf;
  assign memMergeIn_CT$wnnz_Int_r = (! memMergeIn_CT$wnnz_Int_buf[0]);
  assign memMergeIn_CT$wnnz_Int_rbuf_d = (memMergeIn_CT$wnnz_Int_buf[0] ? memMergeIn_CT$wnnz_Int_buf :
                                          memMergeIn_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
    else
      if ((memMergeIn_CT$wnnz_Int_rbuf_r && memMergeIn_CT$wnnz_Int_buf[0]))
        memMergeIn_CT$wnnz_Int_buf <= {132'd0, 1'd0};
      else if (((! memMergeIn_CT$wnnz_Int_rbuf_r) && (! memMergeIn_CT$wnnz_Int_buf[0])))
        memMergeIn_CT$wnnz_Int_buf <= memMergeIn_CT$wnnz_Int_d;
  
  /* dbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_dbuf,MemOut_CT$wnnz_Int) */
  assign memOut_CT$wnnz_Int_rbuf_r = ((! memOut_CT$wnnz_Int_dbuf_d[0]) || memOut_CT$wnnz_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_dbuf_d <= {116'd0, 1'd0};
    else
      if (memOut_CT$wnnz_Int_rbuf_r)
        memOut_CT$wnnz_Int_dbuf_d <= memOut_CT$wnnz_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CT$wnnz_Int) : (memOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > (memOut_CT$wnnz_Int_rbuf,MemOut_CT$wnnz_Int) */
  MemOut_CT$wnnz_Int_t memOut_CT$wnnz_Int_buf;
  assign memOut_CT$wnnz_Int_r = (! memOut_CT$wnnz_Int_buf[0]);
  assign memOut_CT$wnnz_Int_rbuf_d = (memOut_CT$wnnz_Int_buf[0] ? memOut_CT$wnnz_Int_buf :
                                      memOut_CT$wnnz_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
    else
      if ((memOut_CT$wnnz_Int_rbuf_r && memOut_CT$wnnz_Int_buf[0]))
        memOut_CT$wnnz_Int_buf <= {116'd0, 1'd0};
      else if (((! memOut_CT$wnnz_Int_rbuf_r) && (! memOut_CT$wnnz_Int_buf[0])))
        memOut_CT$wnnz_Int_buf <= memOut_CT$wnnz_Int_d;
  
  /* destruct (Ty Pointer_CT$wnnz_Int,
          Dcon Pointer_CT$wnnz_Int) : (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) > [(destructReadIn_CT$wnnz_Int,Word16#)] */
  assign destructReadIn_CT$wnnz_Int_d = {scfarg_0_1_argbuf_d[16:1],
                                         scfarg_0_1_argbuf_d[0]};
  assign scfarg_0_1_argbuf_r = destructReadIn_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon ReadIn_CT$wnnz_Int) : [(destructReadIn_CT$wnnz_Int,Word16#)] > (dconReadIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconReadIn_CT$wnnz_Int_d = ReadIn_CT$wnnz_Int_dc((& {destructReadIn_CT$wnnz_Int_d[0]}), destructReadIn_CT$wnnz_Int_d);
  assign {destructReadIn_CT$wnnz_Int_r} = {1 {(dconReadIn_CT$wnnz_Int_r && dconReadIn_CT$wnnz_Int_d[0])}};
  
  /* destruct (Ty MemOut_CT$wnnz_Int,
          Dcon ReadOut_CT$wnnz_Int) : (memReadOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) > [(readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int)] */
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d = {memReadOut_CT$wnnz_Int_d[116:2],
                                                       memReadOut_CT$wnnz_Int_d[0]};
  assign memReadOut_CT$wnnz_Int_r = readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CT$wnnz_Int) : [(lizzieLet0_1_argbuf,CT$wnnz_Int),
                              (lizzieLet20_1_argbuf,CT$wnnz_Int),
                              (lizzieLet21_1_argbuf,CT$wnnz_Int),
                              (lizzieLet22_1_argbuf,CT$wnnz_Int),
                              (lizzieLet5_1_argbuf,CT$wnnz_Int)] > (writeMerge_choice_CT$wnnz_Int,C5) (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int) */
  logic [4:0] lizzieLet0_1_argbuf_select_d;
  assign lizzieLet0_1_argbuf_select_d = ((| lizzieLet0_1_argbuf_select_q) ? lizzieLet0_1_argbuf_select_q :
                                         (lizzieLet0_1_argbuf_d[0] ? 5'd1 :
                                          (lizzieLet20_1_argbuf_d[0] ? 5'd2 :
                                           (lizzieLet21_1_argbuf_d[0] ? 5'd4 :
                                            (lizzieLet22_1_argbuf_d[0] ? 5'd8 :
                                             (lizzieLet5_1_argbuf_d[0] ? 5'd16 :
                                              5'd0))))));
  logic [4:0] lizzieLet0_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet0_1_argbuf_select_q <= (lizzieLet0_1_argbuf_done ? 5'd0 :
                                       lizzieLet0_1_argbuf_select_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet0_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet0_1_argbuf_emit_q <= (lizzieLet0_1_argbuf_done ? 2'd0 :
                                     lizzieLet0_1_argbuf_emit_d);
  logic [1:0] lizzieLet0_1_argbuf_emit_d;
  assign lizzieLet0_1_argbuf_emit_d = (lizzieLet0_1_argbuf_emit_q | ({writeMerge_choice_CT$wnnz_Int_d[0],
                                                                      writeMerge_data_CT$wnnz_Int_d[0]} & {writeMerge_choice_CT$wnnz_Int_r,
                                                                                                           writeMerge_data_CT$wnnz_Int_r}));
  logic lizzieLet0_1_argbuf_done;
  assign lizzieLet0_1_argbuf_done = (& lizzieLet0_1_argbuf_emit_d);
  assign {lizzieLet5_1_argbuf_r,
          lizzieLet22_1_argbuf_r,
          lizzieLet21_1_argbuf_r,
          lizzieLet20_1_argbuf_r,
          lizzieLet0_1_argbuf_r} = (lizzieLet0_1_argbuf_done ? lizzieLet0_1_argbuf_select_d :
                                    5'd0);
  assign writeMerge_data_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet0_1_argbuf_d :
                                          ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet20_1_argbuf_d :
                                           ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet21_1_argbuf_d :
                                            ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet22_1_argbuf_d :
                                             ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[0])) ? lizzieLet5_1_argbuf_d :
                                              {115'd0, 1'd0})))));
  assign writeMerge_choice_CT$wnnz_Int_d = ((lizzieLet0_1_argbuf_select_d[0] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                            ((lizzieLet0_1_argbuf_select_d[1] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                             ((lizzieLet0_1_argbuf_select_d[2] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                              ((lizzieLet0_1_argbuf_select_d[3] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                               ((lizzieLet0_1_argbuf_select_d[4] && (! lizzieLet0_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CT$wnnz_Int) : (writeMerge_choice_CT$wnnz_Int,C5) (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet20_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet21_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet22_1_argbuf,Pointer_CT$wnnz_Int),
                                                                                                                          (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int)] */
  logic [4:0] demuxWriteResult_CT$wnnz_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CT$wnnz_Int_d[0] && demuxWriteResult_CT$wnnz_Int_d[0]))
      unique case (writeMerge_choice_CT$wnnz_Int_d[3:1])
        3'd0: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd16;
        default: demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CT$wnnz_Int_onehotd = 5'd0;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[0]};
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[1]};
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[2]};
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                   demuxWriteResult_CT$wnnz_Int_onehotd[3]};
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_d = {demuxWriteResult_CT$wnnz_Int_d[16:1],
                                                  demuxWriteResult_CT$wnnz_Int_onehotd[4]};
  assign demuxWriteResult_CT$wnnz_Int_r = (| (demuxWriteResult_CT$wnnz_Int_onehotd & {writeCT$wnnz_IntlizzieLet5_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet22_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet21_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet20_1_argbuf_r,
                                                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_r}));
  assign writeMerge_choice_CT$wnnz_Int_r = demuxWriteResult_CT$wnnz_Int_r;
  
  /* dcon (Ty MemIn_CT$wnnz_Int,
      Dcon WriteIn_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In2,Word16#),
                                   (writeMerge_data_CT$wnnz_Int,CT$wnnz_Int)] > (dconWriteIn_CT$wnnz_Int,MemIn_CT$wnnz_Int) */
  assign dconWriteIn_CT$wnnz_Int_d = WriteIn_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In2_d[0],
                                                                writeMerge_data_CT$wnnz_Int_d[0]}), forkHP1_CT$wnnz_In2_d, writeMerge_data_CT$wnnz_Int_d);
  assign {forkHP1_CT$wnnz_In2_r,
          writeMerge_data_CT$wnnz_Int_r} = {2 {(dconWriteIn_CT$wnnz_Int_r && dconWriteIn_CT$wnnz_Int_d[0])}};
  
  /* dcon (Ty Pointer_CT$wnnz_Int,
      Dcon Pointer_CT$wnnz_Int) : [(forkHP1_CT$wnnz_In3,Word16#)] > (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) */
  assign dconPtr_CT$wnnz_Int_d = Pointer_CT$wnnz_Int_dc((& {forkHP1_CT$wnnz_In3_d[0]}), forkHP1_CT$wnnz_In3_d);
  assign {forkHP1_CT$wnnz_In3_r} = {1 {(dconPtr_CT$wnnz_Int_r && dconPtr_CT$wnnz_Int_d[0])}};
  
  /* demux (Ty MemOut_CT$wnnz_Int,
       Ty Pointer_CT$wnnz_Int) : (memWriteOut_CT$wnnz_Int,MemOut_CT$wnnz_Int) (dconPtr_CT$wnnz_Int,Pointer_CT$wnnz_Int) > [(_45,Pointer_CT$wnnz_Int),
                                                                                                                           (demuxWriteResult_CT$wnnz_Int,Pointer_CT$wnnz_Int)] */
  logic [1:0] dconPtr_CT$wnnz_Int_onehotd;
  always_comb
    if ((memWriteOut_CT$wnnz_Int_d[0] && dconPtr_CT$wnnz_Int_d[0]))
      unique case (memWriteOut_CT$wnnz_Int_d[1:1])
        1'd0: dconPtr_CT$wnnz_Int_onehotd = 2'd1;
        1'd1: dconPtr_CT$wnnz_Int_onehotd = 2'd2;
        default: dconPtr_CT$wnnz_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CT$wnnz_Int_onehotd = 2'd0;
  assign _45_d = {dconPtr_CT$wnnz_Int_d[16:1],
                  dconPtr_CT$wnnz_Int_onehotd[0]};
  assign demuxWriteResult_CT$wnnz_Int_d = {dconPtr_CT$wnnz_Int_d[16:1],
                                           dconPtr_CT$wnnz_Int_onehotd[1]};
  assign dconPtr_CT$wnnz_Int_r = (| (dconPtr_CT$wnnz_Int_onehotd & {demuxWriteResult_CT$wnnz_Int_r,
                                                                    _45_r}));
  assign memWriteOut_CT$wnnz_Int_r = dconPtr_CT$wnnz_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go_1_dummy_write_QTree_Int,Go) > (initHP_QTree_Int,Word16#) */
  assign initHP_QTree_Int_d = {16'd0,
                               go_1_dummy_write_QTree_Int_d[0]};
  assign go_1_dummy_write_QTree_Int_r = initHP_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_QTree_Int1,Go) > (incrHP_QTree_Int,Word16#) */
  assign incrHP_QTree_Int_d = {16'd1, incrHP_QTree_Int1_d[0]};
  assign incrHP_QTree_Int1_r = incrHP_QTree_Int_r;
  
  /* merge (Ty Go) : [(go_2_dummy_write_QTree_Int,Go),
                 (incrHP_QTree_Int2,Go)] > (incrHP_mergeQTree_Int,Go) */
  logic [1:0] incrHP_mergeQTree_Int_selected;
  logic [1:0] incrHP_mergeQTree_Int_select;
  always_comb
    begin
      incrHP_mergeQTree_Int_selected = 2'd0;
      if ((| incrHP_mergeQTree_Int_select))
        incrHP_mergeQTree_Int_selected = incrHP_mergeQTree_Int_select;
      else
        if (go_2_dummy_write_QTree_Int_d[0])
          incrHP_mergeQTree_Int_selected[0] = 1'd1;
        else if (incrHP_QTree_Int2_d[0])
          incrHP_mergeQTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_select <= 2'd0;
    else
      incrHP_mergeQTree_Int_select <= (incrHP_mergeQTree_Int_r ? 2'd0 :
                                       incrHP_mergeQTree_Int_selected);
  always_comb
    if (incrHP_mergeQTree_Int_selected[0])
      incrHP_mergeQTree_Int_d = go_2_dummy_write_QTree_Int_d;
    else if (incrHP_mergeQTree_Int_selected[1])
      incrHP_mergeQTree_Int_d = incrHP_QTree_Int2_d;
    else incrHP_mergeQTree_Int_d = 1'd0;
  assign {incrHP_QTree_Int2_r,
          go_2_dummy_write_QTree_Int_r} = (incrHP_mergeQTree_Int_r ? incrHP_mergeQTree_Int_selected :
                                           2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeQTree_Int_buf,Go) > [(incrHP_QTree_Int1,Go),
                                                 (incrHP_QTree_Int2,Go)] */
  logic [1:0] incrHP_mergeQTree_Int_buf_emitted;
  logic [1:0] incrHP_mergeQTree_Int_buf_done;
  assign incrHP_QTree_Int1_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[0]));
  assign incrHP_QTree_Int2_d = (incrHP_mergeQTree_Int_buf_d[0] && (! incrHP_mergeQTree_Int_buf_emitted[1]));
  assign incrHP_mergeQTree_Int_buf_done = (incrHP_mergeQTree_Int_buf_emitted | ({incrHP_QTree_Int2_d[0],
                                                                                 incrHP_QTree_Int1_d[0]} & {incrHP_QTree_Int2_r,
                                                                                                            incrHP_QTree_Int1_r}));
  assign incrHP_mergeQTree_Int_buf_r = (& incrHP_mergeQTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeQTree_Int_buf_emitted <= (incrHP_mergeQTree_Int_buf_r ? 2'd0 :
                                            incrHP_mergeQTree_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_QTree_Int,Word16#) (forkHP1_QTree_Int,Word16#) > (addHP_QTree_Int,Word16#) */
  assign addHP_QTree_Int_d = {(incrHP_QTree_Int_d[16:1] + forkHP1_QTree_Int_d[16:1]),
                              (incrHP_QTree_Int_d[0] && forkHP1_QTree_Int_d[0])};
  assign {incrHP_QTree_Int_r,
          forkHP1_QTree_Int_r} = {2 {(addHP_QTree_Int_r && addHP_QTree_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_QTree_Int,Word16#),
                      (addHP_QTree_Int,Word16#)] > (mergeHP_QTree_Int,Word16#) */
  logic [1:0] mergeHP_QTree_Int_selected;
  logic [1:0] mergeHP_QTree_Int_select;
  always_comb
    begin
      mergeHP_QTree_Int_selected = 2'd0;
      if ((| mergeHP_QTree_Int_select))
        mergeHP_QTree_Int_selected = mergeHP_QTree_Int_select;
      else
        if (initHP_QTree_Int_d[0]) mergeHP_QTree_Int_selected[0] = 1'd1;
        else if (addHP_QTree_Int_d[0])
          mergeHP_QTree_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_select <= 2'd0;
    else
      mergeHP_QTree_Int_select <= (mergeHP_QTree_Int_r ? 2'd0 :
                                   mergeHP_QTree_Int_selected);
  always_comb
    if (mergeHP_QTree_Int_selected[0])
      mergeHP_QTree_Int_d = initHP_QTree_Int_d;
    else if (mergeHP_QTree_Int_selected[1])
      mergeHP_QTree_Int_d = addHP_QTree_Int_d;
    else mergeHP_QTree_Int_d = {16'd0, 1'd0};
  assign {addHP_QTree_Int_r,
          initHP_QTree_Int_r} = (mergeHP_QTree_Int_r ? mergeHP_QTree_Int_selected :
                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeQTree_Int,Go) > (incrHP_mergeQTree_Int_buf,Go) */
  Go_t incrHP_mergeQTree_Int_bufchan_d;
  logic incrHP_mergeQTree_Int_bufchan_r;
  assign incrHP_mergeQTree_Int_r = ((! incrHP_mergeQTree_Int_bufchan_d[0]) || incrHP_mergeQTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeQTree_Int_r)
        incrHP_mergeQTree_Int_bufchan_d <= incrHP_mergeQTree_Int_d;
  Go_t incrHP_mergeQTree_Int_bufchan_buf;
  assign incrHP_mergeQTree_Int_bufchan_r = (! incrHP_mergeQTree_Int_bufchan_buf[0]);
  assign incrHP_mergeQTree_Int_buf_d = (incrHP_mergeQTree_Int_bufchan_buf[0] ? incrHP_mergeQTree_Int_bufchan_buf :
                                        incrHP_mergeQTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeQTree_Int_buf_r && incrHP_mergeQTree_Int_bufchan_buf[0]))
        incrHP_mergeQTree_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeQTree_Int_buf_r) && (! incrHP_mergeQTree_Int_bufchan_buf[0])))
        incrHP_mergeQTree_Int_bufchan_buf <= incrHP_mergeQTree_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_QTree_Int,Word16#) > (mergeHP_QTree_Int_buf,Word16#) */
  \Word16#_t  mergeHP_QTree_Int_bufchan_d;
  logic mergeHP_QTree_Int_bufchan_r;
  assign mergeHP_QTree_Int_r = ((! mergeHP_QTree_Int_bufchan_d[0]) || mergeHP_QTree_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_QTree_Int_r)
        mergeHP_QTree_Int_bufchan_d <= mergeHP_QTree_Int_d;
  \Word16#_t  mergeHP_QTree_Int_bufchan_buf;
  assign mergeHP_QTree_Int_bufchan_r = (! mergeHP_QTree_Int_bufchan_buf[0]);
  assign mergeHP_QTree_Int_buf_d = (mergeHP_QTree_Int_bufchan_buf[0] ? mergeHP_QTree_Int_bufchan_buf :
                                    mergeHP_QTree_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_QTree_Int_buf_r && mergeHP_QTree_Int_bufchan_buf[0]))
        mergeHP_QTree_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_QTree_Int_buf_r) && (! mergeHP_QTree_Int_bufchan_buf[0])))
        mergeHP_QTree_Int_bufchan_buf <= mergeHP_QTree_Int_bufchan_d;
  
  /* sink (Ty Word16#) : (forkHP1_QTree_Int_snk,Word16#) > */
  assign {forkHP1_QTree_Int_snk_r,
          forkHP1_QTree_Int_snk_dout} = {forkHP1_QTree_Int_snk_rout,
                                         forkHP1_QTree_Int_snk_d};
  
  /* source (Ty Go) : > (\QTree_Int_src,Go) */
  
  /* fork (Ty Go) : (\QTree_Int_src,Go) > [(go_1_dummy_write_QTree_Int,Go),
                                      (go_2_dummy_write_QTree_Int,Go)] */
  logic [1:0] \\QTree_Int_src_emitted ;
  logic [1:0] \\QTree_Int_src_done ;
  assign go_1_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [0]));
  assign go_2_dummy_write_QTree_Int_d = (\\QTree_Int_src_d [0] && (! \\QTree_Int_src_emitted [1]));
  assign \\QTree_Int_src_done  = (\\QTree_Int_src_emitted  | ({go_2_dummy_write_QTree_Int_d[0],
                                                               go_1_dummy_write_QTree_Int_d[0]} & {go_2_dummy_write_QTree_Int_r,
                                                                                                   go_1_dummy_write_QTree_Int_r}));
  assign \\QTree_Int_src_r  = (& \\QTree_Int_src_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \\QTree_Int_src_emitted  <= 2'd0;
    else
      \\QTree_Int_src_emitted  <= (\\QTree_Int_src_r  ? 2'd0 :
                                   \\QTree_Int_src_done );
  
  /* source (Ty QTree_Int) : > (dummy_write_QTree_Int,QTree_Int) */
  
  /* sink (Ty Pointer_QTree_Int) : (dummy_write_QTree_Int_sink,Pointer_QTree_Int) > */
  assign {dummy_write_QTree_Int_sink_r,
          dummy_write_QTree_Int_sink_dout} = {dummy_write_QTree_Int_sink_rout,
                                              dummy_write_QTree_Int_sink_d};
  
  /* fork (Ty Word16#) : (mergeHP_QTree_Int_buf,Word16#) > [(forkHP1_QTree_Int,Word16#),
                                                       (forkHP1_QTree_Int_snk,Word16#),
                                                       (forkHP1_QTree_In3,Word16#),
                                                       (forkHP1_QTree_In4,Word16#)] */
  logic [3:0] mergeHP_QTree_Int_buf_emitted;
  logic [3:0] mergeHP_QTree_Int_buf_done;
  assign forkHP1_QTree_Int_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[0]))};
  assign forkHP1_QTree_Int_snk_d = {mergeHP_QTree_Int_buf_d[16:1],
                                    (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[1]))};
  assign forkHP1_QTree_In3_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[2]))};
  assign forkHP1_QTree_In4_d = {mergeHP_QTree_Int_buf_d[16:1],
                                (mergeHP_QTree_Int_buf_d[0] && (! mergeHP_QTree_Int_buf_emitted[3]))};
  assign mergeHP_QTree_Int_buf_done = (mergeHP_QTree_Int_buf_emitted | ({forkHP1_QTree_In4_d[0],
                                                                         forkHP1_QTree_In3_d[0],
                                                                         forkHP1_QTree_Int_snk_d[0],
                                                                         forkHP1_QTree_Int_d[0]} & {forkHP1_QTree_In4_r,
                                                                                                    forkHP1_QTree_In3_r,
                                                                                                    forkHP1_QTree_Int_snk_r,
                                                                                                    forkHP1_QTree_Int_r}));
  assign mergeHP_QTree_Int_buf_r = (& mergeHP_QTree_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_QTree_Int_buf_emitted <= 4'd0;
    else
      mergeHP_QTree_Int_buf_emitted <= (mergeHP_QTree_Int_buf_r ? 4'd0 :
                                        mergeHP_QTree_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_QTree_Int) : [(dconReadIn_QTree_Int,MemIn_QTree_Int),
                                  (dconWriteIn_QTree_Int,MemIn_QTree_Int)] > (memMergeChoice_QTree_Int,C2) (memMergeIn_QTree_Int,MemIn_QTree_Int) */
  logic [1:0] dconReadIn_QTree_Int_select_d;
  assign dconReadIn_QTree_Int_select_d = ((| dconReadIn_QTree_Int_select_q) ? dconReadIn_QTree_Int_select_q :
                                          (dconReadIn_QTree_Int_d[0] ? 2'd1 :
                                           (dconWriteIn_QTree_Int_d[0] ? 2'd2 :
                                            2'd0)));
  logic [1:0] dconReadIn_QTree_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_select_q <= 2'd0;
    else
      dconReadIn_QTree_Int_select_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                        dconReadIn_QTree_Int_select_d);
  logic [1:0] dconReadIn_QTree_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) dconReadIn_QTree_Int_emit_q <= 2'd0;
    else
      dconReadIn_QTree_Int_emit_q <= (dconReadIn_QTree_Int_done ? 2'd0 :
                                      dconReadIn_QTree_Int_emit_d);
  logic [1:0] dconReadIn_QTree_Int_emit_d;
  assign dconReadIn_QTree_Int_emit_d = (dconReadIn_QTree_Int_emit_q | ({memMergeChoice_QTree_Int_d[0],
                                                                        memMergeIn_QTree_Int_d[0]} & {memMergeChoice_QTree_Int_r,
                                                                                                      memMergeIn_QTree_Int_r}));
  logic dconReadIn_QTree_Int_done;
  assign dconReadIn_QTree_Int_done = (& dconReadIn_QTree_Int_emit_d);
  assign {dconWriteIn_QTree_Int_r,
          dconReadIn_QTree_Int_r} = (dconReadIn_QTree_Int_done ? dconReadIn_QTree_Int_select_d :
                                     2'd0);
  assign memMergeIn_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconReadIn_QTree_Int_d :
                                   ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[0])) ? dconWriteIn_QTree_Int_d :
                                    {83'd0, 1'd0}));
  assign memMergeChoice_QTree_Int_d = ((dconReadIn_QTree_Int_select_d[0] && (! dconReadIn_QTree_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((dconReadIn_QTree_Int_select_d[1] && (! dconReadIn_QTree_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_QTree_Int,
      Ty MemOut_QTree_Int) : (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) > (memOut_QTree_Int,MemOut_QTree_Int) */
  logic [65:0] memMergeIn_QTree_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_QTree_Int_dbuf_address;
  logic [65:0] memMergeIn_QTree_Int_dbuf_din;
  logic [65:0] memOut_QTree_Int_q;
  logic memOut_QTree_Int_valid;
  logic memMergeIn_QTree_Int_dbuf_we;
  logic memOut_QTree_Int_we;
  assign memMergeIn_QTree_Int_dbuf_din = memMergeIn_QTree_Int_dbuf_d[83:18];
  assign memMergeIn_QTree_Int_dbuf_address = memMergeIn_QTree_Int_dbuf_d[17:2];
  assign memMergeIn_QTree_Int_dbuf_we = (memMergeIn_QTree_Int_dbuf_d[1:1] && memMergeIn_QTree_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_QTree_Int_we <= 1'd0;
        memOut_QTree_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_QTree_Int_we <= memMergeIn_QTree_Int_dbuf_we;
        memOut_QTree_Int_valid <= memMergeIn_QTree_Int_dbuf_d[0];
        if (memMergeIn_QTree_Int_dbuf_we)
          begin
            memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address] <= memMergeIn_QTree_Int_dbuf_din;
            memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_din;
          end
        else
          memOut_QTree_Int_q <= memMergeIn_QTree_Int_dbuf_mem[memMergeIn_QTree_Int_dbuf_address];
      end
  assign memOut_QTree_Int_d = {memOut_QTree_Int_q,
                               memOut_QTree_Int_we,
                               memOut_QTree_Int_valid};
  assign memMergeIn_QTree_Int_dbuf_r = ((! memOut_QTree_Int_valid) || memOut_QTree_Int_r);
  logic [31:0] profiling_MemIn_QTree_Int_read;
  logic [31:0] profiling_MemIn_QTree_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_QTree_Int_write <= 0;
        profiling_MemIn_QTree_Int_read <= 0;
      end
    else
      if ((memMergeIn_QTree_Int_dbuf_we == 1'd1))
        profiling_MemIn_QTree_Int_write <= (profiling_MemIn_QTree_Int_write + 1);
      else
        if ((memOut_QTree_Int_valid == 1'd1))
          profiling_MemIn_QTree_Int_read <= (profiling_MemIn_QTree_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_QTree_Int) : (memMergeChoice_QTree_Int,C2) (memOut_QTree_Int_dbuf,MemOut_QTree_Int) > [(memReadOut_QTree_Int,MemOut_QTree_Int),
                                                                                                        (memWriteOut_QTree_Int,MemOut_QTree_Int)] */
  logic [1:0] memOut_QTree_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_QTree_Int_d[0] && memOut_QTree_Int_dbuf_d[0]))
      unique case (memMergeChoice_QTree_Int_d[1:1])
        1'd0: memOut_QTree_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_QTree_Int_dbuf_onehotd = 2'd2;
        default: memOut_QTree_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_QTree_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                   memOut_QTree_Int_dbuf_onehotd[0]};
  assign memWriteOut_QTree_Int_d = {memOut_QTree_Int_dbuf_d[67:1],
                                    memOut_QTree_Int_dbuf_onehotd[1]};
  assign memOut_QTree_Int_dbuf_r = (| (memOut_QTree_Int_dbuf_onehotd & {memWriteOut_QTree_Int_r,
                                                                        memReadOut_QTree_Int_r}));
  assign memMergeChoice_QTree_Int_r = memOut_QTree_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) > (memMergeIn_QTree_Int_dbuf,MemIn_QTree_Int) */
  assign memMergeIn_QTree_Int_rbuf_r = ((! memMergeIn_QTree_Int_dbuf_d[0]) || memMergeIn_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_dbuf_d <= {83'd0, 1'd0};
    else
      if (memMergeIn_QTree_Int_rbuf_r)
        memMergeIn_QTree_Int_dbuf_d <= memMergeIn_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_QTree_Int) : (memMergeIn_QTree_Int,MemIn_QTree_Int) > (memMergeIn_QTree_Int_rbuf,MemIn_QTree_Int) */
  MemIn_QTree_Int_t memMergeIn_QTree_Int_buf;
  assign memMergeIn_QTree_Int_r = (! memMergeIn_QTree_Int_buf[0]);
  assign memMergeIn_QTree_Int_rbuf_d = (memMergeIn_QTree_Int_buf[0] ? memMergeIn_QTree_Int_buf :
                                        memMergeIn_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
    else
      if ((memMergeIn_QTree_Int_rbuf_r && memMergeIn_QTree_Int_buf[0]))
        memMergeIn_QTree_Int_buf <= {83'd0, 1'd0};
      else if (((! memMergeIn_QTree_Int_rbuf_r) && (! memMergeIn_QTree_Int_buf[0])))
        memMergeIn_QTree_Int_buf <= memMergeIn_QTree_Int_d;
  
  /* dbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int_rbuf,MemOut_QTree_Int) > (memOut_QTree_Int_dbuf,MemOut_QTree_Int) */
  assign memOut_QTree_Int_rbuf_r = ((! memOut_QTree_Int_dbuf_d[0]) || memOut_QTree_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_dbuf_d <= {67'd0, 1'd0};
    else
      if (memOut_QTree_Int_rbuf_r)
        memOut_QTree_Int_dbuf_d <= memOut_QTree_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_QTree_Int) : (memOut_QTree_Int,MemOut_QTree_Int) > (memOut_QTree_Int_rbuf,MemOut_QTree_Int) */
  MemOut_QTree_Int_t memOut_QTree_Int_buf;
  assign memOut_QTree_Int_r = (! memOut_QTree_Int_buf[0]);
  assign memOut_QTree_Int_rbuf_d = (memOut_QTree_Int_buf[0] ? memOut_QTree_Int_buf :
                                    memOut_QTree_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) memOut_QTree_Int_buf <= {67'd0, 1'd0};
    else
      if ((memOut_QTree_Int_rbuf_r && memOut_QTree_Int_buf[0]))
        memOut_QTree_Int_buf <= {67'd0, 1'd0};
      else if (((! memOut_QTree_Int_rbuf_r) && (! memOut_QTree_Int_buf[0])))
        memOut_QTree_Int_buf <= memOut_QTree_Int_d;
  
  /* mergectrl (Ty C3,
           Ty Pointer_QTree_Int) : [(m1ahU_1_argbuf,Pointer_QTree_Int),
                                    (m2ai5_1_argbuf,Pointer_QTree_Int),
                                    (wstH_1_1_argbuf,Pointer_QTree_Int)] > (readMerge_choice_QTree_Int,C3) (readMerge_data_QTree_Int,Pointer_QTree_Int) */
  logic [2:0] m1ahU_1_argbuf_select_d;
  assign m1ahU_1_argbuf_select_d = ((| m1ahU_1_argbuf_select_q) ? m1ahU_1_argbuf_select_q :
                                    (m1ahU_1_argbuf_d[0] ? 3'd1 :
                                     (m2ai5_1_argbuf_d[0] ? 3'd2 :
                                      (wstH_1_1_argbuf_d[0] ? 3'd4 :
                                       3'd0))));
  logic [2:0] m1ahU_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ahU_1_argbuf_select_q <= 3'd0;
    else
      m1ahU_1_argbuf_select_q <= (m1ahU_1_argbuf_done ? 3'd0 :
                                  m1ahU_1_argbuf_select_d);
  logic [1:0] m1ahU_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ahU_1_argbuf_emit_q <= 2'd0;
    else
      m1ahU_1_argbuf_emit_q <= (m1ahU_1_argbuf_done ? 2'd0 :
                                m1ahU_1_argbuf_emit_d);
  logic [1:0] m1ahU_1_argbuf_emit_d;
  assign m1ahU_1_argbuf_emit_d = (m1ahU_1_argbuf_emit_q | ({readMerge_choice_QTree_Int_d[0],
                                                            readMerge_data_QTree_Int_d[0]} & {readMerge_choice_QTree_Int_r,
                                                                                              readMerge_data_QTree_Int_r}));
  logic m1ahU_1_argbuf_done;
  assign m1ahU_1_argbuf_done = (& m1ahU_1_argbuf_emit_d);
  assign {wstH_1_1_argbuf_r,
          m2ai5_1_argbuf_r,
          m1ahU_1_argbuf_r} = (m1ahU_1_argbuf_done ? m1ahU_1_argbuf_select_d :
                               3'd0);
  assign readMerge_data_QTree_Int_d = ((m1ahU_1_argbuf_select_d[0] && (! m1ahU_1_argbuf_emit_q[0])) ? m1ahU_1_argbuf_d :
                                       ((m1ahU_1_argbuf_select_d[1] && (! m1ahU_1_argbuf_emit_q[0])) ? m2ai5_1_argbuf_d :
                                        ((m1ahU_1_argbuf_select_d[2] && (! m1ahU_1_argbuf_emit_q[0])) ? wstH_1_1_argbuf_d :
                                         {16'd0, 1'd0})));
  assign readMerge_choice_QTree_Int_d = ((m1ahU_1_argbuf_select_d[0] && (! m1ahU_1_argbuf_emit_q[1])) ? C1_3_dc(1'd1) :
                                         ((m1ahU_1_argbuf_select_d[1] && (! m1ahU_1_argbuf_emit_q[1])) ? C2_3_dc(1'd1) :
                                          ((m1ahU_1_argbuf_select_d[2] && (! m1ahU_1_argbuf_emit_q[1])) ? C3_3_dc(1'd1) :
                                           {2'd0, 1'd0})));
  
  /* demux (Ty C3,
       Ty QTree_Int) : (readMerge_choice_QTree_Int,C3) (destructReadOut_QTree_Int,QTree_Int) > [(readPointer_QTree_Intm1ahU_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_Intm2ai5_1_argbuf,QTree_Int),
                                                                                                (readPointer_QTree_IntwstH_1_1_argbuf,QTree_Int)] */
  logic [2:0] destructReadOut_QTree_Int_onehotd;
  always_comb
    if ((readMerge_choice_QTree_Int_d[0] && destructReadOut_QTree_Int_d[0]))
      unique case (readMerge_choice_QTree_Int_d[2:1])
        2'd0: destructReadOut_QTree_Int_onehotd = 3'd1;
        2'd1: destructReadOut_QTree_Int_onehotd = 3'd2;
        2'd2: destructReadOut_QTree_Int_onehotd = 3'd4;
        default: destructReadOut_QTree_Int_onehotd = 3'd0;
      endcase
    else destructReadOut_QTree_Int_onehotd = 3'd0;
  assign readPointer_QTree_Intm1ahU_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[0]};
  assign readPointer_QTree_Intm2ai5_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                  destructReadOut_QTree_Int_onehotd[1]};
  assign readPointer_QTree_IntwstH_1_1_argbuf_d = {destructReadOut_QTree_Int_d[66:1],
                                                   destructReadOut_QTree_Int_onehotd[2]};
  assign destructReadOut_QTree_Int_r = (| (destructReadOut_QTree_Int_onehotd & {readPointer_QTree_IntwstH_1_1_argbuf_r,
                                                                                readPointer_QTree_Intm2ai5_1_argbuf_r,
                                                                                readPointer_QTree_Intm1ahU_1_argbuf_r}));
  assign readMerge_choice_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* destruct (Ty Pointer_QTree_Int,
          Dcon Pointer_QTree_Int) : (readMerge_data_QTree_Int,Pointer_QTree_Int) > [(destructReadIn_QTree_Int,Word16#)] */
  assign destructReadIn_QTree_Int_d = {readMerge_data_QTree_Int_d[16:1],
                                       readMerge_data_QTree_Int_d[0]};
  assign readMerge_data_QTree_Int_r = destructReadIn_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon ReadIn_QTree_Int) : [(destructReadIn_QTree_Int,Word16#)] > (dconReadIn_QTree_Int,MemIn_QTree_Int) */
  assign dconReadIn_QTree_Int_d = ReadIn_QTree_Int_dc((& {destructReadIn_QTree_Int_d[0]}), destructReadIn_QTree_Int_d);
  assign {destructReadIn_QTree_Int_r} = {1 {(dconReadIn_QTree_Int_r && dconReadIn_QTree_Int_d[0])}};
  
  /* destruct (Ty MemOut_QTree_Int,
          Dcon ReadOut_QTree_Int) : (memReadOut_QTree_Int,MemOut_QTree_Int) > [(destructReadOut_QTree_Int,QTree_Int)] */
  assign destructReadOut_QTree_Int_d = {memReadOut_QTree_Int_d[67:2],
                                        memReadOut_QTree_Int_d[0]};
  assign memReadOut_QTree_Int_r = destructReadOut_QTree_Int_r;
  
  /* mergectrl (Ty C10,
           Ty QTree_Int) : [(lizzieLet10_1_argbuf,QTree_Int),
                            (lizzieLet12_1_1_argbuf,QTree_Int),
                            (lizzieLet14_1_argbuf,QTree_Int),
                            (lizzieLet16_1_argbuf,QTree_Int),
                            (lizzieLet27_1_argbuf,QTree_Int),
                            (lizzieLet32_1_argbuf,QTree_Int),
                            (lizzieLet7_1_argbuf,QTree_Int),
                            (lizzieLet8_1_argbuf,QTree_Int),
                            (lizzieLet9_1_argbuf,QTree_Int),
                            (dummy_write_QTree_Int,QTree_Int)] > (writeMerge_choice_QTree_Int,C10) (writeMerge_data_QTree_Int,QTree_Int) */
  logic [9:0] lizzieLet10_1_argbuf_select_d;
  assign lizzieLet10_1_argbuf_select_d = ((| lizzieLet10_1_argbuf_select_q) ? lizzieLet10_1_argbuf_select_q :
                                          (lizzieLet10_1_argbuf_d[0] ? 10'd1 :
                                           (lizzieLet12_1_1_argbuf_d[0] ? 10'd2 :
                                            (lizzieLet14_1_argbuf_d[0] ? 10'd4 :
                                             (lizzieLet16_1_argbuf_d[0] ? 10'd8 :
                                              (lizzieLet27_1_argbuf_d[0] ? 10'd16 :
                                               (lizzieLet32_1_argbuf_d[0] ? 10'd32 :
                                                (lizzieLet7_1_argbuf_d[0] ? 10'd64 :
                                                 (lizzieLet8_1_argbuf_d[0] ? 10'd128 :
                                                  (lizzieLet9_1_argbuf_d[0] ? 10'd256 :
                                                   (dummy_write_QTree_Int_d[0] ? 10'd512 :
                                                    10'd0)))))))))));
  logic [9:0] lizzieLet10_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_select_q <= 10'd0;
    else
      lizzieLet10_1_argbuf_select_q <= (lizzieLet10_1_argbuf_done ? 10'd0 :
                                        lizzieLet10_1_argbuf_select_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet10_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet10_1_argbuf_emit_q <= (lizzieLet10_1_argbuf_done ? 2'd0 :
                                      lizzieLet10_1_argbuf_emit_d);
  logic [1:0] lizzieLet10_1_argbuf_emit_d;
  assign lizzieLet10_1_argbuf_emit_d = (lizzieLet10_1_argbuf_emit_q | ({writeMerge_choice_QTree_Int_d[0],
                                                                        writeMerge_data_QTree_Int_d[0]} & {writeMerge_choice_QTree_Int_r,
                                                                                                           writeMerge_data_QTree_Int_r}));
  logic lizzieLet10_1_argbuf_done;
  assign lizzieLet10_1_argbuf_done = (& lizzieLet10_1_argbuf_emit_d);
  assign {dummy_write_QTree_Int_r,
          lizzieLet9_1_argbuf_r,
          lizzieLet8_1_argbuf_r,
          lizzieLet7_1_argbuf_r,
          lizzieLet32_1_argbuf_r,
          lizzieLet27_1_argbuf_r,
          lizzieLet16_1_argbuf_r,
          lizzieLet14_1_argbuf_r,
          lizzieLet12_1_1_argbuf_r,
          lizzieLet10_1_argbuf_r} = (lizzieLet10_1_argbuf_done ? lizzieLet10_1_argbuf_select_d :
                                     10'd0);
  assign writeMerge_data_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet10_1_argbuf_d :
                                        ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet12_1_1_argbuf_d :
                                         ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet14_1_argbuf_d :
                                          ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet16_1_argbuf_d :
                                           ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet27_1_argbuf_d :
                                            ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet32_1_argbuf_d :
                                             ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet7_1_argbuf_d :
                                              ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet8_1_argbuf_d :
                                               ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[0])) ? lizzieLet9_1_argbuf_d :
                                                ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[0])) ? dummy_write_QTree_Int_d :
                                                 {66'd0, 1'd0}))))))))));
  assign writeMerge_choice_QTree_Int_d = ((lizzieLet10_1_argbuf_select_d[0] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C1_10_dc(1'd1) :
                                          ((lizzieLet10_1_argbuf_select_d[1] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C2_10_dc(1'd1) :
                                           ((lizzieLet10_1_argbuf_select_d[2] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C3_10_dc(1'd1) :
                                            ((lizzieLet10_1_argbuf_select_d[3] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C4_10_dc(1'd1) :
                                             ((lizzieLet10_1_argbuf_select_d[4] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C5_10_dc(1'd1) :
                                              ((lizzieLet10_1_argbuf_select_d[5] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C6_10_dc(1'd1) :
                                               ((lizzieLet10_1_argbuf_select_d[6] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C7_10_dc(1'd1) :
                                                ((lizzieLet10_1_argbuf_select_d[7] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C8_10_dc(1'd1) :
                                                 ((lizzieLet10_1_argbuf_select_d[8] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C9_10_dc(1'd1) :
                                                  ((lizzieLet10_1_argbuf_select_d[9] && (! lizzieLet10_1_argbuf_emit_q[1])) ? C10_10_dc(1'd1) :
                                                   {4'd0, 1'd0}))))))))));
  
  /* demux (Ty C10,
       Ty Pointer_QTree_Int) : (writeMerge_choice_QTree_Int,C10) (demuxWriteResult_QTree_Int,Pointer_QTree_Int) > [(writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet12_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet14_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet27_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int),
                                                                                                                   (dummy_write_QTree_Int_sink,Pointer_QTree_Int)] */
  logic [9:0] demuxWriteResult_QTree_Int_onehotd;
  always_comb
    if ((writeMerge_choice_QTree_Int_d[0] && demuxWriteResult_QTree_Int_d[0]))
      unique case (writeMerge_choice_QTree_Int_d[4:1])
        4'd0: demuxWriteResult_QTree_Int_onehotd = 10'd1;
        4'd1: demuxWriteResult_QTree_Int_onehotd = 10'd2;
        4'd2: demuxWriteResult_QTree_Int_onehotd = 10'd4;
        4'd3: demuxWriteResult_QTree_Int_onehotd = 10'd8;
        4'd4: demuxWriteResult_QTree_Int_onehotd = 10'd16;
        4'd5: demuxWriteResult_QTree_Int_onehotd = 10'd32;
        4'd6: demuxWriteResult_QTree_Int_onehotd = 10'd64;
        4'd7: demuxWriteResult_QTree_Int_onehotd = 10'd128;
        4'd8: demuxWriteResult_QTree_Int_onehotd = 10'd256;
        4'd9: demuxWriteResult_QTree_Int_onehotd = 10'd512;
        default: demuxWriteResult_QTree_Int_onehotd = 10'd0;
      endcase
    else demuxWriteResult_QTree_Int_onehotd = 10'd0;
  assign writeQTree_IntlizzieLet10_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[0]};
  assign writeQTree_IntlizzieLet12_1_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                   demuxWriteResult_QTree_Int_onehotd[1]};
  assign writeQTree_IntlizzieLet14_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[2]};
  assign writeQTree_IntlizzieLet16_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[3]};
  assign writeQTree_IntlizzieLet27_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[4]};
  assign writeQTree_IntlizzieLet32_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                 demuxWriteResult_QTree_Int_onehotd[5]};
  assign writeQTree_IntlizzieLet7_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[6]};
  assign writeQTree_IntlizzieLet8_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[7]};
  assign writeQTree_IntlizzieLet9_1_argbuf_d = {demuxWriteResult_QTree_Int_d[16:1],
                                                demuxWriteResult_QTree_Int_onehotd[8]};
  assign dummy_write_QTree_Int_sink_d = {demuxWriteResult_QTree_Int_d[16:1],
                                         demuxWriteResult_QTree_Int_onehotd[9]};
  assign demuxWriteResult_QTree_Int_r = (| (demuxWriteResult_QTree_Int_onehotd & {dummy_write_QTree_Int_sink_r,
                                                                                  writeQTree_IntlizzieLet9_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet8_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet7_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet32_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet27_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet16_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet14_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet12_1_1_argbuf_r,
                                                                                  writeQTree_IntlizzieLet10_1_argbuf_r}));
  assign writeMerge_choice_QTree_Int_r = demuxWriteResult_QTree_Int_r;
  
  /* dcon (Ty MemIn_QTree_Int,
      Dcon WriteIn_QTree_Int) : [(forkHP1_QTree_In3,Word16#),
                                 (writeMerge_data_QTree_Int,QTree_Int)] > (dconWriteIn_QTree_Int,MemIn_QTree_Int) */
  assign dconWriteIn_QTree_Int_d = WriteIn_QTree_Int_dc((& {forkHP1_QTree_In3_d[0],
                                                            writeMerge_data_QTree_Int_d[0]}), forkHP1_QTree_In3_d, writeMerge_data_QTree_Int_d);
  assign {forkHP1_QTree_In3_r,
          writeMerge_data_QTree_Int_r} = {2 {(dconWriteIn_QTree_Int_r && dconWriteIn_QTree_Int_d[0])}};
  
  /* dcon (Ty Pointer_QTree_Int,
      Dcon Pointer_QTree_Int) : [(forkHP1_QTree_In4,Word16#)] > (dconPtr_QTree_Int,Pointer_QTree_Int) */
  assign dconPtr_QTree_Int_d = Pointer_QTree_Int_dc((& {forkHP1_QTree_In4_d[0]}), forkHP1_QTree_In4_d);
  assign {forkHP1_QTree_In4_r} = {1 {(dconPtr_QTree_Int_r && dconPtr_QTree_Int_d[0])}};
  
  /* demux (Ty MemOut_QTree_Int,
       Ty Pointer_QTree_Int) : (memWriteOut_QTree_Int,MemOut_QTree_Int) (dconPtr_QTree_Int,Pointer_QTree_Int) > [(_44,Pointer_QTree_Int),
                                                                                                                 (demuxWriteResult_QTree_Int,Pointer_QTree_Int)] */
  logic [1:0] dconPtr_QTree_Int_onehotd;
  always_comb
    if ((memWriteOut_QTree_Int_d[0] && dconPtr_QTree_Int_d[0]))
      unique case (memWriteOut_QTree_Int_d[1:1])
        1'd0: dconPtr_QTree_Int_onehotd = 2'd1;
        1'd1: dconPtr_QTree_Int_onehotd = 2'd2;
        default: dconPtr_QTree_Int_onehotd = 2'd0;
      endcase
    else dconPtr_QTree_Int_onehotd = 2'd0;
  assign _44_d = {dconPtr_QTree_Int_d[16:1],
                  dconPtr_QTree_Int_onehotd[0]};
  assign demuxWriteResult_QTree_Int_d = {dconPtr_QTree_Int_d[16:1],
                                         dconPtr_QTree_Int_onehotd[1]};
  assign dconPtr_QTree_Int_r = (| (dconPtr_QTree_Int_onehotd & {demuxWriteResult_QTree_Int_r,
                                                                _44_r}));
  assign memWriteOut_QTree_Int_r = dconPtr_QTree_Int_r;
  
  /* const (Ty Word16#,
       Lit 0) : (go__9,Go) > (initHP_CTf'_f'_Int_Int_Int_Int,Word16#) */
  assign \initHP_CTf'_f'_Int_Int_Int_Int_d  = {16'd0, go__9_d[0]};
  assign go__9_r = \initHP_CTf'_f'_Int_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf'_f'_Int_Int_Int_Int1,Go) > (incrHP_CTf'_f'_Int_Int_Int_Int,Word16#) */
  assign \incrHP_CTf'_f'_Int_Int_Int_Int_d  = {16'd1,
                                               \incrHP_CTf'_f'_Int_Int_Int_Int1_d [0]};
  assign \incrHP_CTf'_f'_Int_Int_Int_Int1_r  = \incrHP_CTf'_f'_Int_Int_Int_Int_r ;
  
  /* merge (Ty Go) : [(go__10,Go),
                 (incrHP_CTf'_f'_Int_Int_Int_Int2,Go)] > (incrHP_mergeCTf'_f'_Int_Int_Int_Int,Go) */
  logic [1:0] \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected ;
  logic [1:0] \incrHP_mergeCTf'_f'_Int_Int_Int_Int_select ;
  always_comb
    begin
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected  = 2'd0;
      if ((| \incrHP_mergeCTf'_f'_Int_Int_Int_Int_select ))
        \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected  = \incrHP_mergeCTf'_f'_Int_Int_Int_Int_select ;
      else
        if (go__10_d[0])
          \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected [0] = 1'd1;
        else if (\incrHP_CTf'_f'_Int_Int_Int_Int2_d [0])
          \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_select  <= 2'd0;
    else
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_select  <= (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_r  ? 2'd0 :
                                                       \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected );
  always_comb
    if (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected [0])
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_d  = go__10_d;
    else if (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected [1])
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_d  = \incrHP_CTf'_f'_Int_Int_Int_Int2_d ;
    else \incrHP_mergeCTf'_f'_Int_Int_Int_Int_d  = 1'd0;
  assign {\incrHP_CTf'_f'_Int_Int_Int_Int2_r ,
          go__10_r} = (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_r  ? \incrHP_mergeCTf'_f'_Int_Int_Int_Int_selected  :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf,Go) > [(incrHP_CTf'_f'_Int_Int_Int_Int1,Go),
                                                               (incrHP_CTf'_f'_Int_Int_Int_Int2,Go)] */
  logic [1:0] \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted ;
  logic [1:0] \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_done ;
  assign \incrHP_CTf'_f'_Int_Int_Int_Int1_d  = (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted [0]));
  assign \incrHP_CTf'_f'_Int_Int_Int_Int2_d  = (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_d [0] && (! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted [1]));
  assign \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_done  = (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted  | ({\incrHP_CTf'_f'_Int_Int_Int_Int2_d [0],
                                                                                                                 \incrHP_CTf'_f'_Int_Int_Int_Int1_d [0]} & {\incrHP_CTf'_f'_Int_Int_Int_Int2_r ,
                                                                                                                                                            \incrHP_CTf'_f'_Int_Int_Int_Int1_r }));
  assign \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_r  = (& \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted  <= 2'd0;
    else
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_emitted  <= (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_r  ? 2'd0 :
                                                            \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_done );
  
  /* op_add (Ty Word16#) : (incrHP_CTf'_f'_Int_Int_Int_Int,Word16#) (forkHP1_CTf'_f'_Int_Int_Int_Int,Word16#) > (addHP_CTf'_f'_Int_Int_Int_Int,Word16#) */
  assign \addHP_CTf'_f'_Int_Int_Int_Int_d  = {(\incrHP_CTf'_f'_Int_Int_Int_Int_d [16:1] + \forkHP1_CTf'_f'_Int_Int_Int_Int_d [16:1]),
                                              (\incrHP_CTf'_f'_Int_Int_Int_Int_d [0] && \forkHP1_CTf'_f'_Int_Int_Int_Int_d [0])};
  assign {\incrHP_CTf'_f'_Int_Int_Int_Int_r ,
          \forkHP1_CTf'_f'_Int_Int_Int_Int_r } = {2 {(\addHP_CTf'_f'_Int_Int_Int_Int_r  && \addHP_CTf'_f'_Int_Int_Int_Int_d [0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf'_f'_Int_Int_Int_Int,Word16#),
                      (addHP_CTf'_f'_Int_Int_Int_Int,Word16#)] > (mergeHP_CTf'_f'_Int_Int_Int_Int,Word16#) */
  logic [1:0] \mergeHP_CTf'_f'_Int_Int_Int_Int_selected ;
  logic [1:0] \mergeHP_CTf'_f'_Int_Int_Int_Int_select ;
  always_comb
    begin
      \mergeHP_CTf'_f'_Int_Int_Int_Int_selected  = 2'd0;
      if ((| \mergeHP_CTf'_f'_Int_Int_Int_Int_select ))
        \mergeHP_CTf'_f'_Int_Int_Int_Int_selected  = \mergeHP_CTf'_f'_Int_Int_Int_Int_select ;
      else
        if (\initHP_CTf'_f'_Int_Int_Int_Int_d [0])
          \mergeHP_CTf'_f'_Int_Int_Int_Int_selected [0] = 1'd1;
        else if (\addHP_CTf'_f'_Int_Int_Int_Int_d [0])
          \mergeHP_CTf'_f'_Int_Int_Int_Int_selected [1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_Int_Int_Int_select  <= 2'd0;
    else
      \mergeHP_CTf'_f'_Int_Int_Int_Int_select  <= (\mergeHP_CTf'_f'_Int_Int_Int_Int_r  ? 2'd0 :
                                                   \mergeHP_CTf'_f'_Int_Int_Int_Int_selected );
  always_comb
    if (\mergeHP_CTf'_f'_Int_Int_Int_Int_selected [0])
      \mergeHP_CTf'_f'_Int_Int_Int_Int_d  = \initHP_CTf'_f'_Int_Int_Int_Int_d ;
    else if (\mergeHP_CTf'_f'_Int_Int_Int_Int_selected [1])
      \mergeHP_CTf'_f'_Int_Int_Int_Int_d  = \addHP_CTf'_f'_Int_Int_Int_Int_d ;
    else \mergeHP_CTf'_f'_Int_Int_Int_Int_d  = {16'd0, 1'd0};
  assign {\addHP_CTf'_f'_Int_Int_Int_Int_r ,
          \initHP_CTf'_f'_Int_Int_Int_Int_r } = (\mergeHP_CTf'_f'_Int_Int_Int_Int_r  ? \mergeHP_CTf'_f'_Int_Int_Int_Int_selected  :
                                                 2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf'_f'_Int_Int_Int_Int,Go) > (incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf,Go) */
  Go_t \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d ;
  logic \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_r ;
  assign \incrHP_mergeCTf'_f'_Int_Int_Int_Int_r  = ((! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d [0]) || \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d  <= 1'd0;
    else
      if (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_r )
        \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d  <= \incrHP_mergeCTf'_f'_Int_Int_Int_Int_d ;
  Go_t \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf ;
  assign \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_r  = (! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf [0]);
  assign \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_d  = (\incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf [0] ? \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf  :
                                                        \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf  <= 1'd0;
    else
      if ((\incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_r  && \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf [0]))
        \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf  <= 1'd0;
      else if (((! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_buf_r ) && (! \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf [0])))
        \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_buf  <= \incrHP_mergeCTf'_f'_Int_Int_Int_Int_bufchan_d ;
  
  /* buf (Ty Word16#) : (mergeHP_CTf'_f'_Int_Int_Int_Int,Word16#) > (mergeHP_CTf'_f'_Int_Int_Int_Int_buf,Word16#) */
  \Word16#_t  \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d ;
  logic \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_r ;
  assign \mergeHP_CTf'_f'_Int_Int_Int_Int_r  = ((! \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d [0]) || \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\mergeHP_CTf'_f'_Int_Int_Int_Int_r )
        \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d  <= \mergeHP_CTf'_f'_Int_Int_Int_Int_d ;
  \Word16#_t  \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf ;
  assign \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_r  = (! \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf [0]);
  assign \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d  = (\mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf [0] ? \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf  :
                                                    \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_r  && \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf [0]))
        \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_r ) && (! \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf [0])))
        \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_buf  <= \mergeHP_CTf'_f'_Int_Int_Int_Int_bufchan_d ;
  
  /* fork (Ty Word16#) : (mergeHP_CTf'_f'_Int_Int_Int_Int_buf,Word16#) > [(forkHP1_CTf'_f'_Int_Int_Int_Int,Word16#),
                                                                     (forkHP1_CTf'_f'_Int_Int_Int_In2,Word16#),
                                                                     (forkHP1_CTf'_f'_Int_Int_Int_In3,Word16#)] */
  logic [2:0] \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted ;
  logic [2:0] \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_done ;
  assign \forkHP1_CTf'_f'_Int_Int_Int_Int_d  = {\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [16:1],
                                                (\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted [0]))};
  assign \forkHP1_CTf'_f'_Int_Int_Int_In2_d  = {\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [16:1],
                                                (\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted [1]))};
  assign \forkHP1_CTf'_f'_Int_Int_Int_In3_d  = {\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [16:1],
                                                (\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_d [0] && (! \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted [2]))};
  assign \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_done  = (\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted  | ({\forkHP1_CTf'_f'_Int_Int_Int_In3_d [0],
                                                                                                         \forkHP1_CTf'_f'_Int_Int_Int_In2_d [0],
                                                                                                         \forkHP1_CTf'_f'_Int_Int_Int_Int_d [0]} & {\forkHP1_CTf'_f'_Int_Int_Int_In3_r ,
                                                                                                                                                    \forkHP1_CTf'_f'_Int_Int_Int_In2_r ,
                                                                                                                                                    \forkHP1_CTf'_f'_Int_Int_Int_Int_r }));
  assign \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_r  = (& \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted  <= 3'd0;
    else
      \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_emitted  <= (\mergeHP_CTf'_f'_Int_Int_Int_Int_buf_r  ? 3'd0 :
                                                        \mergeHP_CTf'_f'_Int_Int_Int_Int_buf_done );
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf'_f'_Int_Int_Int_Int) : [(dconReadIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int),
                                                (dconWriteIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int)] > (memMergeChoice_CTf'_f'_Int_Int_Int_Int,C2) (memMergeIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int) */
  logic [1:0] \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d ;
  assign \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d  = ((| \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_q ) ? \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_q  :
                                                          (\dconReadIn_CTf'_f'_Int_Int_Int_Int_d [0] ? 2'd1 :
                                                           (\dconWriteIn_CTf'_f'_Int_Int_Int_Int_d [0] ? 2'd2 :
                                                            2'd0)));
  logic [1:0] \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_q  <= 2'd0;
    else
      \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_q  <= (\dconReadIn_CTf'_f'_Int_Int_Int_Int_done  ? 2'd0 :
                                                        \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d );
  logic [1:0] \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q  <= 2'd0;
    else
      \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q  <= (\dconReadIn_CTf'_f'_Int_Int_Int_Int_done  ? 2'd0 :
                                                      \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_d );
  logic [1:0] \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_d ;
  assign \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_d  = (\dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q  | ({\memMergeChoice_CTf'_f'_Int_Int_Int_Int_d [0],
                                                                                                        \memMergeIn_CTf'_f'_Int_Int_Int_Int_d [0]} & {\memMergeChoice_CTf'_f'_Int_Int_Int_Int_r ,
                                                                                                                                                      \memMergeIn_CTf'_f'_Int_Int_Int_Int_r }));
  logic \dconReadIn_CTf'_f'_Int_Int_Int_Int_done ;
  assign \dconReadIn_CTf'_f'_Int_Int_Int_Int_done  = (& \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_d );
  assign {\dconWriteIn_CTf'_f'_Int_Int_Int_Int_r ,
          \dconReadIn_CTf'_f'_Int_Int_Int_Int_r } = (\dconReadIn_CTf'_f'_Int_Int_Int_Int_done  ? \dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d  :
                                                     2'd0);
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_d  = ((\dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d [0] && (! \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q [0])) ? \dconReadIn_CTf'_f'_Int_Int_Int_Int_d  :
                                                   ((\dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d [1] && (! \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q [0])) ? \dconWriteIn_CTf'_f'_Int_Int_Int_Int_d  :
                                                    {116'd0, 1'd0}));
  assign \memMergeChoice_CTf'_f'_Int_Int_Int_Int_d  = ((\dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d [0] && (! \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q [1])) ? C1_2_dc(1'd1) :
                                                       ((\dconReadIn_CTf'_f'_Int_Int_Int_Int_select_d [1] && (! \dconReadIn_CTf'_f'_Int_Int_Int_Int_emit_q [1])) ? C2_2_dc(1'd1) :
                                                        {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf'_f'_Int_Int_Int_Int,
      Ty MemOut_CTf'_f'_Int_Int_Int_Int) : (memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf,MemIn_CTf'_f'_Int_Int_Int_Int) > (memOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int) */
  logic [98:0] \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_mem [65535:0];
  logic [15:0] \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_address ;
  logic [98:0] \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_din ;
  logic [98:0] \memOut_CTf'_f'_Int_Int_Int_Int_q ;
  logic \memOut_CTf'_f'_Int_Int_Int_Int_valid ;
  logic \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_we ;
  logic \memOut_CTf'_f'_Int_Int_Int_Int_we ;
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_din  = \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [116:18];
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_address  = \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [17:2];
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_we  = (\memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [1:1] && \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \memOut_CTf'_f'_Int_Int_Int_Int_we  <= 1'd0;
        \memOut_CTf'_f'_Int_Int_Int_Int_valid  <= 1'd0;
      end
    else
      begin
        \memOut_CTf'_f'_Int_Int_Int_Int_we  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_we ;
        \memOut_CTf'_f'_Int_Int_Int_Int_valid  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [0];
        if (\memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_we )
          begin
            \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_mem [\memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_address ] <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_din ;
            \memOut_CTf'_f'_Int_Int_Int_Int_q  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_din ;
          end
        else
          \memOut_CTf'_f'_Int_Int_Int_Int_q  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_mem [\memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_address ];
      end
  assign \memOut_CTf'_f'_Int_Int_Int_Int_d  = {\memOut_CTf'_f'_Int_Int_Int_Int_q ,
                                               \memOut_CTf'_f'_Int_Int_Int_Int_we ,
                                               \memOut_CTf'_f'_Int_Int_Int_Int_valid };
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_r  = ((! \memOut_CTf'_f'_Int_Int_Int_Int_valid ) || \memOut_CTf'_f'_Int_Int_Int_Int_r );
  logic [31:0] \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_read ;
  logic [31:0] \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_write ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_write  <= 0;
        \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_read  <= 0;
      end
    else
      if ((\memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_we  == 1'd1))
        \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_write  <= (\profiling_MemIn_CTf'_f'_Int_Int_Int_Int_write  + 1);
      else
        if ((\memOut_CTf'_f'_Int_Int_Int_Int_valid  == 1'd1))
          \profiling_MemIn_CTf'_f'_Int_Int_Int_Int_read  <= (\profiling_MemIn_CTf'_f'_Int_Int_Int_Int_read  + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf'_f'_Int_Int_Int_Int) : (memMergeChoice_CTf'_f'_Int_Int_Int_Int,C2) (memOut_CTf'_f'_Int_Int_Int_Int_dbuf,MemOut_CTf'_f'_Int_Int_Int_Int) > [(memReadOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                (memWriteOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int)] */
  logic [1:0] \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd ;
  always_comb
    if ((\memMergeChoice_CTf'_f'_Int_Int_Int_Int_d [0] && \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d [0]))
      unique case (\memMergeChoice_CTf'_f'_Int_Int_Int_Int_d [1:1])
        1'd0: \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd  = 2'd1;
        1'd1: \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd  = 2'd2;
        default: \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd  = 2'd0;
      endcase
    else \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd  = 2'd0;
  assign \memReadOut_CTf'_f'_Int_Int_Int_Int_d  = {\memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d [100:1],
                                                   \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd [0]};
  assign \memWriteOut_CTf'_f'_Int_Int_Int_Int_d  = {\memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d [100:1],
                                                    \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd [1]};
  assign \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_r  = (| (\memOut_CTf'_f'_Int_Int_Int_Int_dbuf_onehotd  & {\memWriteOut_CTf'_f'_Int_Int_Int_Int_r ,
                                                                                                        \memReadOut_CTf'_f'_Int_Int_Int_Int_r }));
  assign \memMergeChoice_CTf'_f'_Int_Int_Int_Int_r  = \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_r ;
  
  /* dbuf (Ty MemIn_CTf'_f'_Int_Int_Int_Int) : (memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf,MemIn_CTf'_f'_Int_Int_Int_Int) > (memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf,MemIn_CTf'_f'_Int_Int_Int_Int) */
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_r  = ((! \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d [0]) || \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d  <= {116'd0, 1'd0};
    else
      if (\memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_r )
        \memMergeIn_CTf'_f'_Int_Int_Int_Int_dbuf_d  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemIn_CTf'_f'_Int_Int_Int_Int) : (memMergeIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int) > (memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf,MemIn_CTf'_f'_Int_Int_Int_Int) */
  \MemIn_CTf'_f'_Int_Int_Int_Int_t  \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf ;
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_r  = (! \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf [0]);
  assign \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_d  = (\memMergeIn_CTf'_f'_Int_Int_Int_Int_buf [0] ? \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf  :
                                                        \memMergeIn_CTf'_f'_Int_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf  <= {116'd0, 1'd0};
    else
      if ((\memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_r  && \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf [0]))
        \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf  <= {116'd0, 1'd0};
      else if (((! \memMergeIn_CTf'_f'_Int_Int_Int_Int_rbuf_r ) && (! \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf [0])))
        \memMergeIn_CTf'_f'_Int_Int_Int_Int_buf  <= \memMergeIn_CTf'_f'_Int_Int_Int_Int_d ;
  
  /* dbuf (Ty MemOut_CTf'_f'_Int_Int_Int_Int) : (memOut_CTf'_f'_Int_Int_Int_Int_rbuf,MemOut_CTf'_f'_Int_Int_Int_Int) > (memOut_CTf'_f'_Int_Int_Int_Int_dbuf,MemOut_CTf'_f'_Int_Int_Int_Int) */
  assign \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_r  = ((! \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d [0]) || \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d  <= {100'd0, 1'd0};
    else
      if (\memOut_CTf'_f'_Int_Int_Int_Int_rbuf_r )
        \memOut_CTf'_f'_Int_Int_Int_Int_dbuf_d  <= \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_d ;
  
  /* rbuf (Ty MemOut_CTf'_f'_Int_Int_Int_Int) : (memOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int) > (memOut_CTf'_f'_Int_Int_Int_Int_rbuf,MemOut_CTf'_f'_Int_Int_Int_Int) */
  \MemOut_CTf'_f'_Int_Int_Int_Int_t  \memOut_CTf'_f'_Int_Int_Int_Int_buf ;
  assign \memOut_CTf'_f'_Int_Int_Int_Int_r  = (! \memOut_CTf'_f'_Int_Int_Int_Int_buf [0]);
  assign \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_d  = (\memOut_CTf'_f'_Int_Int_Int_Int_buf [0] ? \memOut_CTf'_f'_Int_Int_Int_Int_buf  :
                                                    \memOut_CTf'_f'_Int_Int_Int_Int_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \memOut_CTf'_f'_Int_Int_Int_Int_buf  <= {100'd0, 1'd0};
    else
      if ((\memOut_CTf'_f'_Int_Int_Int_Int_rbuf_r  && \memOut_CTf'_f'_Int_Int_Int_Int_buf [0]))
        \memOut_CTf'_f'_Int_Int_Int_Int_buf  <= {100'd0, 1'd0};
      else if (((! \memOut_CTf'_f'_Int_Int_Int_Int_rbuf_r ) && (! \memOut_CTf'_f'_Int_Int_Int_Int_buf [0])))
        \memOut_CTf'_f'_Int_Int_Int_Int_buf  <= \memOut_CTf'_f'_Int_Int_Int_Int_d ;
  
  /* destruct (Ty Pointer_CTf'_f'_Int_Int_Int_Int,
          Dcon Pointer_CTf'_f'_Int_Int_Int_Int) : (scfarg_0_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > [(destructReadIn_CTf'_f'_Int_Int_Int_Int,Word16#)] */
  assign \destructReadIn_CTf'_f'_Int_Int_Int_Int_d  = {scfarg_0_1_1_argbuf_d[16:1],
                                                       scfarg_0_1_1_argbuf_d[0]};
  assign scfarg_0_1_1_argbuf_r = \destructReadIn_CTf'_f'_Int_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTf'_f'_Int_Int_Int_Int,
      Dcon ReadIn_CTf'_f'_Int_Int_Int_Int) : [(destructReadIn_CTf'_f'_Int_Int_Int_Int,Word16#)] > (dconReadIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int) */
  assign \dconReadIn_CTf'_f'_Int_Int_Int_Int_d  = \ReadIn_CTf'_f'_Int_Int_Int_Int_dc ((& {\destructReadIn_CTf'_f'_Int_Int_Int_Int_d [0]}), \destructReadIn_CTf'_f'_Int_Int_Int_Int_d );
  assign {\destructReadIn_CTf'_f'_Int_Int_Int_Int_r } = {1 {(\dconReadIn_CTf'_f'_Int_Int_Int_Int_r  && \dconReadIn_CTf'_f'_Int_Int_Int_Int_d [0])}};
  
  /* destruct (Ty MemOut_CTf'_f'_Int_Int_Int_Int,
          Dcon ReadOut_CTf'_f'_Int_Int_Int_Int) : (memReadOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int) > [(readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf,CTf'_f'_Int_Int_Int_Int)] */
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_d  = {\memReadOut_CTf'_f'_Int_Int_Int_Int_d [100:2],
                                                                       \memReadOut_CTf'_f'_Int_Int_Int_Int_d [0]};
  assign \memReadOut_CTf'_f'_Int_Int_Int_Int_r  = \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_r ;
  
  /* mergectrl (Ty C5,
           Ty CTf'_f'_Int_Int_Int_Int) : [(lizzieLet11_2_1_argbuf,CTf'_f'_Int_Int_Int_Int),
                                          (lizzieLet17_1_argbuf,CTf'_f'_Int_Int_Int_Int),
                                          (lizzieLet24_1_argbuf,CTf'_f'_Int_Int_Int_Int),
                                          (lizzieLet25_1_argbuf,CTf'_f'_Int_Int_Int_Int),
                                          (lizzieLet26_1_argbuf,CTf'_f'_Int_Int_Int_Int)] > (writeMerge_choice_CTf'_f'_Int_Int_Int_Int,C5) (writeMerge_data_CTf'_f'_Int_Int_Int_Int,CTf'_f'_Int_Int_Int_Int) */
  logic [4:0] lizzieLet11_2_1_argbuf_select_d;
  assign lizzieLet11_2_1_argbuf_select_d = ((| lizzieLet11_2_1_argbuf_select_q) ? lizzieLet11_2_1_argbuf_select_q :
                                            (lizzieLet11_2_1_argbuf_d[0] ? 5'd1 :
                                             (lizzieLet17_1_argbuf_d[0] ? 5'd2 :
                                              (lizzieLet24_1_argbuf_d[0] ? 5'd4 :
                                               (lizzieLet25_1_argbuf_d[0] ? 5'd8 :
                                                (lizzieLet26_1_argbuf_d[0] ? 5'd16 :
                                                 5'd0))))));
  logic [4:0] lizzieLet11_2_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_2_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet11_2_1_argbuf_select_q <= (lizzieLet11_2_1_argbuf_done ? 5'd0 :
                                          lizzieLet11_2_1_argbuf_select_d);
  logic [1:0] lizzieLet11_2_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet11_2_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet11_2_1_argbuf_emit_q <= (lizzieLet11_2_1_argbuf_done ? 2'd0 :
                                        lizzieLet11_2_1_argbuf_emit_d);
  logic [1:0] lizzieLet11_2_1_argbuf_emit_d;
  assign lizzieLet11_2_1_argbuf_emit_d = (lizzieLet11_2_1_argbuf_emit_q | ({\writeMerge_choice_CTf'_f'_Int_Int_Int_Int_d [0],
                                                                            \writeMerge_data_CTf'_f'_Int_Int_Int_Int_d [0]} & {\writeMerge_choice_CTf'_f'_Int_Int_Int_Int_r ,
                                                                                                                               \writeMerge_data_CTf'_f'_Int_Int_Int_Int_r }));
  logic lizzieLet11_2_1_argbuf_done;
  assign lizzieLet11_2_1_argbuf_done = (& lizzieLet11_2_1_argbuf_emit_d);
  assign {lizzieLet26_1_argbuf_r,
          lizzieLet25_1_argbuf_r,
          lizzieLet24_1_argbuf_r,
          lizzieLet17_1_argbuf_r,
          lizzieLet11_2_1_argbuf_r} = (lizzieLet11_2_1_argbuf_done ? lizzieLet11_2_1_argbuf_select_d :
                                       5'd0);
  assign \writeMerge_data_CTf'_f'_Int_Int_Int_Int_d  = ((lizzieLet11_2_1_argbuf_select_d[0] && (! lizzieLet11_2_1_argbuf_emit_q[0])) ? lizzieLet11_2_1_argbuf_d :
                                                        ((lizzieLet11_2_1_argbuf_select_d[1] && (! lizzieLet11_2_1_argbuf_emit_q[0])) ? lizzieLet17_1_argbuf_d :
                                                         ((lizzieLet11_2_1_argbuf_select_d[2] && (! lizzieLet11_2_1_argbuf_emit_q[0])) ? lizzieLet24_1_argbuf_d :
                                                          ((lizzieLet11_2_1_argbuf_select_d[3] && (! lizzieLet11_2_1_argbuf_emit_q[0])) ? lizzieLet25_1_argbuf_d :
                                                           ((lizzieLet11_2_1_argbuf_select_d[4] && (! lizzieLet11_2_1_argbuf_emit_q[0])) ? lizzieLet26_1_argbuf_d :
                                                            {99'd0, 1'd0})))));
  assign \writeMerge_choice_CTf'_f'_Int_Int_Int_Int_d  = ((lizzieLet11_2_1_argbuf_select_d[0] && (! lizzieLet11_2_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                          ((lizzieLet11_2_1_argbuf_select_d[1] && (! lizzieLet11_2_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                           ((lizzieLet11_2_1_argbuf_select_d[2] && (! lizzieLet11_2_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                            ((lizzieLet11_2_1_argbuf_select_d[3] && (! lizzieLet11_2_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                             ((lizzieLet11_2_1_argbuf_select_d[4] && (! lizzieLet11_2_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                              {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeMerge_choice_CTf'_f'_Int_Int_Int_Int,C5) (demuxWriteResult_CTf'_f'_Int_Int_Int_Int,Pointer_CTf'_f'_Int_Int_Int_Int) > [(writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                          (writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                          (writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                          (writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                          (writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [4:0] \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd ;
  always_comb
    if ((\writeMerge_choice_CTf'_f'_Int_Int_Int_Int_d [0] && \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [0]))
      unique case (\writeMerge_choice_CTf'_f'_Int_Int_Int_Int_d [3:1])
        3'd0: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd1;
        3'd1: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd2;
        3'd2: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd4;
        3'd3: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd8;
        3'd4: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd16;
        default: \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd0;
      endcase
    else \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  = 5'd0;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                                   \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd [0]};
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                                 \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd [1]};
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                                 \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd [2]};
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                                 \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd [3]};
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_d  = {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                                 \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd [4]};
  assign \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_r  = (| (\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_onehotd  & {\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_r ,
                                                                                                                  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_r ,
                                                                                                                  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_r ,
                                                                                                                  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_r ,
                                                                                                                  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_r }));
  assign \writeMerge_choice_CTf'_f'_Int_Int_Int_Int_r  = \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_r ;
  
  /* dcon (Ty MemIn_CTf'_f'_Int_Int_Int_Int,
      Dcon WriteIn_CTf'_f'_Int_Int_Int_Int) : [(forkHP1_CTf'_f'_Int_Int_Int_In2,Word16#),
                                               (writeMerge_data_CTf'_f'_Int_Int_Int_Int,CTf'_f'_Int_Int_Int_Int)] > (dconWriteIn_CTf'_f'_Int_Int_Int_Int,MemIn_CTf'_f'_Int_Int_Int_Int) */
  assign \dconWriteIn_CTf'_f'_Int_Int_Int_Int_d  = \WriteIn_CTf'_f'_Int_Int_Int_Int_dc ((& {\forkHP1_CTf'_f'_Int_Int_Int_In2_d [0],
                                                                                            \writeMerge_data_CTf'_f'_Int_Int_Int_Int_d [0]}), \forkHP1_CTf'_f'_Int_Int_Int_In2_d , \writeMerge_data_CTf'_f'_Int_Int_Int_Int_d );
  assign {\forkHP1_CTf'_f'_Int_Int_Int_In2_r ,
          \writeMerge_data_CTf'_f'_Int_Int_Int_Int_r } = {2 {(\dconWriteIn_CTf'_f'_Int_Int_Int_Int_r  && \dconWriteIn_CTf'_f'_Int_Int_Int_Int_d [0])}};
  
  /* dcon (Ty Pointer_CTf'_f'_Int_Int_Int_Int,
      Dcon Pointer_CTf'_f'_Int_Int_Int_Int) : [(forkHP1_CTf'_f'_Int_Int_Int_In3,Word16#)] > (dconPtr_CTf'_f'_Int_Int_Int_Int,Pointer_CTf'_f'_Int_Int_Int_Int) */
  assign \dconPtr_CTf'_f'_Int_Int_Int_Int_d  = \Pointer_CTf'_f'_Int_Int_Int_Int_dc ((& {\forkHP1_CTf'_f'_Int_Int_Int_In3_d [0]}), \forkHP1_CTf'_f'_Int_Int_Int_In3_d );
  assign {\forkHP1_CTf'_f'_Int_Int_Int_In3_r } = {1 {(\dconPtr_CTf'_f'_Int_Int_Int_Int_r  && \dconPtr_CTf'_f'_Int_Int_Int_Int_d [0])}};
  
  /* demux (Ty MemOut_CTf'_f'_Int_Int_Int_Int,
       Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (memWriteOut_CTf'_f'_Int_Int_Int_Int,MemOut_CTf'_f'_Int_Int_Int_Int) (dconPtr_CTf'_f'_Int_Int_Int_Int,Pointer_CTf'_f'_Int_Int_Int_Int) > [(_43,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                                                                                       (demuxWriteResult_CTf'_f'_Int_Int_Int_Int,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [1:0] \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd ;
  always_comb
    if ((\memWriteOut_CTf'_f'_Int_Int_Int_Int_d [0] && \dconPtr_CTf'_f'_Int_Int_Int_Int_d [0]))
      unique case (\memWriteOut_CTf'_f'_Int_Int_Int_Int_d [1:1])
        1'd0: \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd  = 2'd1;
        1'd1: \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd  = 2'd2;
        default: \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd  = 2'd0;
      endcase
    else \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd  = 2'd0;
  assign _43_d = {\dconPtr_CTf'_f'_Int_Int_Int_Int_d [16:1],
                  \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd [0]};
  assign \demuxWriteResult_CTf'_f'_Int_Int_Int_Int_d  = {\dconPtr_CTf'_f'_Int_Int_Int_Int_d [16:1],
                                                         \dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd [1]};
  assign \dconPtr_CTf'_f'_Int_Int_Int_Int_r  = (| (\dconPtr_CTf'_f'_Int_Int_Int_Int_onehotd  & {\demuxWriteResult_CTf'_f'_Int_Int_Int_Int_r ,
                                                                                                _43_r}));
  assign \memWriteOut_CTf'_f'_Int_Int_Int_Int_r  = \dconPtr_CTf'_f'_Int_Int_Int_Int_r ;
  
  /* const (Ty Word16#,
       Lit 0) : (go__11,Go) > (initHP_CTf_f_Int_Int_Int_Int,Word16#) */
  assign initHP_CTf_f_Int_Int_Int_Int_d = {16'd0, go__11_d[0]};
  assign go__11_r = initHP_CTf_f_Int_Int_Int_Int_r;
  
  /* const (Ty Word16#,
       Lit 1) : (incrHP_CTf_f_Int_Int_Int_Int1,Go) > (incrHP_CTf_f_Int_Int_Int_Int,Word16#) */
  assign incrHP_CTf_f_Int_Int_Int_Int_d = {16'd1,
                                           incrHP_CTf_f_Int_Int_Int_Int1_d[0]};
  assign incrHP_CTf_f_Int_Int_Int_Int1_r = incrHP_CTf_f_Int_Int_Int_Int_r;
  
  /* merge (Ty Go) : [(go__12,Go),
                 (incrHP_CTf_f_Int_Int_Int_Int2,Go)] > (incrHP_mergeCTf_f_Int_Int_Int_Int,Go) */
  logic [1:0] incrHP_mergeCTf_f_Int_Int_Int_Int_selected;
  logic [1:0] incrHP_mergeCTf_f_Int_Int_Int_Int_select;
  always_comb
    begin
      incrHP_mergeCTf_f_Int_Int_Int_Int_selected = 2'd0;
      if ((| incrHP_mergeCTf_f_Int_Int_Int_Int_select))
        incrHP_mergeCTf_f_Int_Int_Int_Int_selected = incrHP_mergeCTf_f_Int_Int_Int_Int_select;
      else
        if (go__12_d[0])
          incrHP_mergeCTf_f_Int_Int_Int_Int_selected[0] = 1'd1;
        else if (incrHP_CTf_f_Int_Int_Int_Int2_d[0])
          incrHP_mergeCTf_f_Int_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTf_f_Int_Int_Int_Int_select <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_Int_Int_Int_select <= (incrHP_mergeCTf_f_Int_Int_Int_Int_r ? 2'd0 :
                                                   incrHP_mergeCTf_f_Int_Int_Int_Int_selected);
  always_comb
    if (incrHP_mergeCTf_f_Int_Int_Int_Int_selected[0])
      incrHP_mergeCTf_f_Int_Int_Int_Int_d = go__12_d;
    else if (incrHP_mergeCTf_f_Int_Int_Int_Int_selected[1])
      incrHP_mergeCTf_f_Int_Int_Int_Int_d = incrHP_CTf_f_Int_Int_Int_Int2_d;
    else incrHP_mergeCTf_f_Int_Int_Int_Int_d = 1'd0;
  assign {incrHP_CTf_f_Int_Int_Int_Int2_r,
          go__12_r} = (incrHP_mergeCTf_f_Int_Int_Int_Int_r ? incrHP_mergeCTf_f_Int_Int_Int_Int_selected :
                       2'd0);
  
  /* fork (Ty Go) : (incrHP_mergeCTf_f_Int_Int_Int_Int_buf,Go) > [(incrHP_CTf_f_Int_Int_Int_Int1,Go),
                                                             (incrHP_CTf_f_Int_Int_Int_Int2,Go)] */
  logic [1:0] incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted;
  logic [1:0] incrHP_mergeCTf_f_Int_Int_Int_Int_buf_done;
  assign incrHP_CTf_f_Int_Int_Int_Int1_d = (incrHP_mergeCTf_f_Int_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted[0]));
  assign incrHP_CTf_f_Int_Int_Int_Int2_d = (incrHP_mergeCTf_f_Int_Int_Int_Int_buf_d[0] && (! incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted[1]));
  assign incrHP_mergeCTf_f_Int_Int_Int_Int_buf_done = (incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted | ({incrHP_CTf_f_Int_Int_Int_Int2_d[0],
                                                                                                         incrHP_CTf_f_Int_Int_Int_Int1_d[0]} & {incrHP_CTf_f_Int_Int_Int_Int2_r,
                                                                                                                                                incrHP_CTf_f_Int_Int_Int_Int1_r}));
  assign incrHP_mergeCTf_f_Int_Int_Int_Int_buf_r = (& incrHP_mergeCTf_f_Int_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted <= 2'd0;
    else
      incrHP_mergeCTf_f_Int_Int_Int_Int_buf_emitted <= (incrHP_mergeCTf_f_Int_Int_Int_Int_buf_r ? 2'd0 :
                                                        incrHP_mergeCTf_f_Int_Int_Int_Int_buf_done);
  
  /* op_add (Ty Word16#) : (incrHP_CTf_f_Int_Int_Int_Int,Word16#) (forkHP1_CTf_f_Int_Int_Int_Int,Word16#) > (addHP_CTf_f_Int_Int_Int_Int,Word16#) */
  assign addHP_CTf_f_Int_Int_Int_Int_d = {(incrHP_CTf_f_Int_Int_Int_Int_d[16:1] + forkHP1_CTf_f_Int_Int_Int_Int_d[16:1]),
                                          (incrHP_CTf_f_Int_Int_Int_Int_d[0] && forkHP1_CTf_f_Int_Int_Int_Int_d[0])};
  assign {incrHP_CTf_f_Int_Int_Int_Int_r,
          forkHP1_CTf_f_Int_Int_Int_Int_r} = {2 {(addHP_CTf_f_Int_Int_Int_Int_r && addHP_CTf_f_Int_Int_Int_Int_d[0])}};
  
  /* merge (Ty Word16#) : [(initHP_CTf_f_Int_Int_Int_Int,Word16#),
                      (addHP_CTf_f_Int_Int_Int_Int,Word16#)] > (mergeHP_CTf_f_Int_Int_Int_Int,Word16#) */
  logic [1:0] mergeHP_CTf_f_Int_Int_Int_Int_selected;
  logic [1:0] mergeHP_CTf_f_Int_Int_Int_Int_select;
  always_comb
    begin
      mergeHP_CTf_f_Int_Int_Int_Int_selected = 2'd0;
      if ((| mergeHP_CTf_f_Int_Int_Int_Int_select))
        mergeHP_CTf_f_Int_Int_Int_Int_selected = mergeHP_CTf_f_Int_Int_Int_Int_select;
      else
        if (initHP_CTf_f_Int_Int_Int_Int_d[0])
          mergeHP_CTf_f_Int_Int_Int_Int_selected[0] = 1'd1;
        else if (addHP_CTf_f_Int_Int_Int_Int_d[0])
          mergeHP_CTf_f_Int_Int_Int_Int_selected[1] = 1'd1;
    end
  always_ff @(posedge clk)
    if ((reset == 1'd1)) mergeHP_CTf_f_Int_Int_Int_Int_select <= 2'd0;
    else
      mergeHP_CTf_f_Int_Int_Int_Int_select <= (mergeHP_CTf_f_Int_Int_Int_Int_r ? 2'd0 :
                                               mergeHP_CTf_f_Int_Int_Int_Int_selected);
  always_comb
    if (mergeHP_CTf_f_Int_Int_Int_Int_selected[0])
      mergeHP_CTf_f_Int_Int_Int_Int_d = initHP_CTf_f_Int_Int_Int_Int_d;
    else if (mergeHP_CTf_f_Int_Int_Int_Int_selected[1])
      mergeHP_CTf_f_Int_Int_Int_Int_d = addHP_CTf_f_Int_Int_Int_Int_d;
    else mergeHP_CTf_f_Int_Int_Int_Int_d = {16'd0, 1'd0};
  assign {addHP_CTf_f_Int_Int_Int_Int_r,
          initHP_CTf_f_Int_Int_Int_Int_r} = (mergeHP_CTf_f_Int_Int_Int_Int_r ? mergeHP_CTf_f_Int_Int_Int_Int_selected :
                                             2'd0);
  
  /* buf (Ty Go) : (incrHP_mergeCTf_f_Int_Int_Int_Int,Go) > (incrHP_mergeCTf_f_Int_Int_Int_Int_buf,Go) */
  Go_t incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d;
  logic incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_r;
  assign incrHP_mergeCTf_f_Int_Int_Int_Int_r = ((! incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d[0]) || incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d <= 1'd0;
    else
      if (incrHP_mergeCTf_f_Int_Int_Int_Int_r)
        incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d <= incrHP_mergeCTf_f_Int_Int_Int_Int_d;
  Go_t incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf;
  assign incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_r = (! incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf[0]);
  assign incrHP_mergeCTf_f_Int_Int_Int_Int_buf_d = (incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf[0] ? incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf :
                                                    incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf <= 1'd0;
    else
      if ((incrHP_mergeCTf_f_Int_Int_Int_Int_buf_r && incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf[0]))
        incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf <= 1'd0;
      else if (((! incrHP_mergeCTf_f_Int_Int_Int_Int_buf_r) && (! incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf[0])))
        incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_buf <= incrHP_mergeCTf_f_Int_Int_Int_Int_bufchan_d;
  
  /* buf (Ty Word16#) : (mergeHP_CTf_f_Int_Int_Int_Int,Word16#) > (mergeHP_CTf_f_Int_Int_Int_Int_buf,Word16#) */
  \Word16#_t  mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d;
  logic mergeHP_CTf_f_Int_Int_Int_Int_bufchan_r;
  assign mergeHP_CTf_f_Int_Int_Int_Int_r = ((! mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d[0]) || mergeHP_CTf_f_Int_Int_Int_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (mergeHP_CTf_f_Int_Int_Int_Int_r)
        mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d <= mergeHP_CTf_f_Int_Int_Int_Int_d;
  \Word16#_t  mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf;
  assign mergeHP_CTf_f_Int_Int_Int_Int_bufchan_r = (! mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf[0]);
  assign mergeHP_CTf_f_Int_Int_Int_Int_buf_d = (mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf[0] ? mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf :
                                                mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((mergeHP_CTf_f_Int_Int_Int_Int_buf_r && mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf[0]))
        mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! mergeHP_CTf_f_Int_Int_Int_Int_buf_r) && (! mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf[0])))
        mergeHP_CTf_f_Int_Int_Int_Int_bufchan_buf <= mergeHP_CTf_f_Int_Int_Int_Int_bufchan_d;
  
  /* fork (Ty Word16#) : (mergeHP_CTf_f_Int_Int_Int_Int_buf,Word16#) > [(forkHP1_CTf_f_Int_Int_Int_Int,Word16#),
                                                                   (forkHP1_CTf_f_Int_Int_Int_In2,Word16#),
                                                                   (forkHP1_CTf_f_Int_Int_Int_In3,Word16#)] */
  logic [2:0] mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted;
  logic [2:0] mergeHP_CTf_f_Int_Int_Int_Int_buf_done;
  assign forkHP1_CTf_f_Int_Int_Int_Int_d = {mergeHP_CTf_f_Int_Int_Int_Int_buf_d[16:1],
                                            (mergeHP_CTf_f_Int_Int_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted[0]))};
  assign forkHP1_CTf_f_Int_Int_Int_In2_d = {mergeHP_CTf_f_Int_Int_Int_Int_buf_d[16:1],
                                            (mergeHP_CTf_f_Int_Int_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted[1]))};
  assign forkHP1_CTf_f_Int_Int_Int_In3_d = {mergeHP_CTf_f_Int_Int_Int_Int_buf_d[16:1],
                                            (mergeHP_CTf_f_Int_Int_Int_Int_buf_d[0] && (! mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted[2]))};
  assign mergeHP_CTf_f_Int_Int_Int_Int_buf_done = (mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted | ({forkHP1_CTf_f_Int_Int_Int_In3_d[0],
                                                                                                 forkHP1_CTf_f_Int_Int_Int_In2_d[0],
                                                                                                 forkHP1_CTf_f_Int_Int_Int_Int_d[0]} & {forkHP1_CTf_f_Int_Int_Int_In3_r,
                                                                                                                                        forkHP1_CTf_f_Int_Int_Int_In2_r,
                                                                                                                                        forkHP1_CTf_f_Int_Int_Int_Int_r}));
  assign mergeHP_CTf_f_Int_Int_Int_Int_buf_r = (& mergeHP_CTf_f_Int_Int_Int_Int_buf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted <= 3'd0;
    else
      mergeHP_CTf_f_Int_Int_Int_Int_buf_emitted <= (mergeHP_CTf_f_Int_Int_Int_Int_buf_r ? 3'd0 :
                                                    mergeHP_CTf_f_Int_Int_Int_Int_buf_done);
  
  /* mergectrl (Ty C2,
           Ty MemIn_CTf_f_Int_Int_Int_Int) : [(dconReadIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int),
                                              (dconWriteIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int)] > (memMergeChoice_CTf_f_Int_Int_Int_Int,C2) (memMergeIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int) */
  logic [1:0] dconReadIn_CTf_f_Int_Int_Int_Int_select_d;
  assign dconReadIn_CTf_f_Int_Int_Int_Int_select_d = ((| dconReadIn_CTf_f_Int_Int_Int_Int_select_q) ? dconReadIn_CTf_f_Int_Int_Int_Int_select_q :
                                                      (dconReadIn_CTf_f_Int_Int_Int_Int_d[0] ? 2'd1 :
                                                       (dconWriteIn_CTf_f_Int_Int_Int_Int_d[0] ? 2'd2 :
                                                        2'd0)));
  logic [1:0] dconReadIn_CTf_f_Int_Int_Int_Int_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTf_f_Int_Int_Int_Int_select_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_Int_Int_Int_select_q <= (dconReadIn_CTf_f_Int_Int_Int_Int_done ? 2'd0 :
                                                    dconReadIn_CTf_f_Int_Int_Int_Int_select_d);
  logic [1:0] dconReadIn_CTf_f_Int_Int_Int_Int_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      dconReadIn_CTf_f_Int_Int_Int_Int_emit_q <= 2'd0;
    else
      dconReadIn_CTf_f_Int_Int_Int_Int_emit_q <= (dconReadIn_CTf_f_Int_Int_Int_Int_done ? 2'd0 :
                                                  dconReadIn_CTf_f_Int_Int_Int_Int_emit_d);
  logic [1:0] dconReadIn_CTf_f_Int_Int_Int_Int_emit_d;
  assign dconReadIn_CTf_f_Int_Int_Int_Int_emit_d = (dconReadIn_CTf_f_Int_Int_Int_Int_emit_q | ({memMergeChoice_CTf_f_Int_Int_Int_Int_d[0],
                                                                                                memMergeIn_CTf_f_Int_Int_Int_Int_d[0]} & {memMergeChoice_CTf_f_Int_Int_Int_Int_r,
                                                                                                                                          memMergeIn_CTf_f_Int_Int_Int_Int_r}));
  logic dconReadIn_CTf_f_Int_Int_Int_Int_done;
  assign dconReadIn_CTf_f_Int_Int_Int_Int_done = (& dconReadIn_CTf_f_Int_Int_Int_Int_emit_d);
  assign {dconWriteIn_CTf_f_Int_Int_Int_Int_r,
          dconReadIn_CTf_f_Int_Int_Int_Int_r} = (dconReadIn_CTf_f_Int_Int_Int_Int_done ? dconReadIn_CTf_f_Int_Int_Int_Int_select_d :
                                                 2'd0);
  assign memMergeIn_CTf_f_Int_Int_Int_Int_d = ((dconReadIn_CTf_f_Int_Int_Int_Int_select_d[0] && (! dconReadIn_CTf_f_Int_Int_Int_Int_emit_q[0])) ? dconReadIn_CTf_f_Int_Int_Int_Int_d :
                                               ((dconReadIn_CTf_f_Int_Int_Int_Int_select_d[1] && (! dconReadIn_CTf_f_Int_Int_Int_Int_emit_q[0])) ? dconWriteIn_CTf_f_Int_Int_Int_Int_d :
                                                {100'd0, 1'd0}));
  assign memMergeChoice_CTf_f_Int_Int_Int_Int_d = ((dconReadIn_CTf_f_Int_Int_Int_Int_select_d[0] && (! dconReadIn_CTf_f_Int_Int_Int_Int_emit_q[1])) ? C1_2_dc(1'd1) :
                                                   ((dconReadIn_CTf_f_Int_Int_Int_Int_select_d[1] && (! dconReadIn_CTf_f_Int_Int_Int_Int_emit_q[1])) ? C2_2_dc(1'd1) :
                                                    {1'd0, 1'd0}));
  
  /* bram (Ty MemIn_CTf_f_Int_Int_Int_Int,
      Ty MemOut_CTf_f_Int_Int_Int_Int) : (memMergeIn_CTf_f_Int_Int_Int_Int_dbuf,MemIn_CTf_f_Int_Int_Int_Int) > (memOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int) */
  logic [82:0] memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_mem[65535:0];
  logic [15:0] memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_address;
  logic [82:0] memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_din;
  logic [82:0] memOut_CTf_f_Int_Int_Int_Int_q;
  logic memOut_CTf_f_Int_Int_Int_Int_valid;
  logic memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_we;
  logic memOut_CTf_f_Int_Int_Int_Int_we;
  assign memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_din = memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[100:18];
  assign memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_address = memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[17:2];
  assign memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_we = (memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[1:1] && memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[0]);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        memOut_CTf_f_Int_Int_Int_Int_we <= 1'd0;
        memOut_CTf_f_Int_Int_Int_Int_valid <= 1'd0;
      end
    else
      begin
        memOut_CTf_f_Int_Int_Int_Int_we <= memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_we;
        memOut_CTf_f_Int_Int_Int_Int_valid <= memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[0];
        if (memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_we)
          begin
            memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_mem[memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_address] <= memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_din;
            memOut_CTf_f_Int_Int_Int_Int_q <= memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_din;
          end
        else
          memOut_CTf_f_Int_Int_Int_Int_q <= memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_mem[memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_address];
      end
  assign memOut_CTf_f_Int_Int_Int_Int_d = {memOut_CTf_f_Int_Int_Int_Int_q,
                                           memOut_CTf_f_Int_Int_Int_Int_we,
                                           memOut_CTf_f_Int_Int_Int_Int_valid};
  assign memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_r = ((! memOut_CTf_f_Int_Int_Int_Int_valid) || memOut_CTf_f_Int_Int_Int_Int_r);
  logic [31:0] profiling_MemIn_CTf_f_Int_Int_Int_Int_read;
  logic [31:0] profiling_MemIn_CTf_f_Int_Int_Int_Int_write;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      begin
        profiling_MemIn_CTf_f_Int_Int_Int_Int_write <= 0;
        profiling_MemIn_CTf_f_Int_Int_Int_Int_read <= 0;
      end
    else
      if ((memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_we == 1'd1))
        profiling_MemIn_CTf_f_Int_Int_Int_Int_write <= (profiling_MemIn_CTf_f_Int_Int_Int_Int_write + 1);
      else
        if ((memOut_CTf_f_Int_Int_Int_Int_valid == 1'd1))
          profiling_MemIn_CTf_f_Int_Int_Int_Int_read <= (profiling_MemIn_CTf_f_Int_Int_Int_Int_read + 1);
  
  /* demux (Ty C2,
       Ty MemOut_CTf_f_Int_Int_Int_Int) : (memMergeChoice_CTf_f_Int_Int_Int_Int,C2) (memOut_CTf_f_Int_Int_Int_Int_dbuf,MemOut_CTf_f_Int_Int_Int_Int) > [(memReadOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int),
                                                                                                                                                        (memWriteOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int)] */
  logic [1:0] memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd;
  always_comb
    if ((memMergeChoice_CTf_f_Int_Int_Int_Int_d[0] && memOut_CTf_f_Int_Int_Int_Int_dbuf_d[0]))
      unique case (memMergeChoice_CTf_f_Int_Int_Int_Int_d[1:1])
        1'd0: memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd = 2'd1;
        1'd1: memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd = 2'd2;
        default: memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd = 2'd0;
      endcase
    else memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd = 2'd0;
  assign memReadOut_CTf_f_Int_Int_Int_Int_d = {memOut_CTf_f_Int_Int_Int_Int_dbuf_d[84:1],
                                               memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd[0]};
  assign memWriteOut_CTf_f_Int_Int_Int_Int_d = {memOut_CTf_f_Int_Int_Int_Int_dbuf_d[84:1],
                                                memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd[1]};
  assign memOut_CTf_f_Int_Int_Int_Int_dbuf_r = (| (memOut_CTf_f_Int_Int_Int_Int_dbuf_onehotd & {memWriteOut_CTf_f_Int_Int_Int_Int_r,
                                                                                                memReadOut_CTf_f_Int_Int_Int_Int_r}));
  assign memMergeChoice_CTf_f_Int_Int_Int_Int_r = memOut_CTf_f_Int_Int_Int_Int_dbuf_r;
  
  /* dbuf (Ty MemIn_CTf_f_Int_Int_Int_Int) : (memMergeIn_CTf_f_Int_Int_Int_Int_rbuf,MemIn_CTf_f_Int_Int_Int_Int) > (memMergeIn_CTf_f_Int_Int_Int_Int_dbuf,MemIn_CTf_f_Int_Int_Int_Int) */
  assign memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_r = ((! memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d[0]) || memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d <= {100'd0, 1'd0};
    else
      if (memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_r)
        memMergeIn_CTf_f_Int_Int_Int_Int_dbuf_d <= memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemIn_CTf_f_Int_Int_Int_Int) : (memMergeIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int) > (memMergeIn_CTf_f_Int_Int_Int_Int_rbuf,MemIn_CTf_f_Int_Int_Int_Int) */
  MemIn_CTf_f_Int_Int_Int_Int_t memMergeIn_CTf_f_Int_Int_Int_Int_buf;
  assign memMergeIn_CTf_f_Int_Int_Int_Int_r = (! memMergeIn_CTf_f_Int_Int_Int_Int_buf[0]);
  assign memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_d = (memMergeIn_CTf_f_Int_Int_Int_Int_buf[0] ? memMergeIn_CTf_f_Int_Int_Int_Int_buf :
                                                    memMergeIn_CTf_f_Int_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memMergeIn_CTf_f_Int_Int_Int_Int_buf <= {100'd0, 1'd0};
    else
      if ((memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_r && memMergeIn_CTf_f_Int_Int_Int_Int_buf[0]))
        memMergeIn_CTf_f_Int_Int_Int_Int_buf <= {100'd0, 1'd0};
      else if (((! memMergeIn_CTf_f_Int_Int_Int_Int_rbuf_r) && (! memMergeIn_CTf_f_Int_Int_Int_Int_buf[0])))
        memMergeIn_CTf_f_Int_Int_Int_Int_buf <= memMergeIn_CTf_f_Int_Int_Int_Int_d;
  
  /* dbuf (Ty MemOut_CTf_f_Int_Int_Int_Int) : (memOut_CTf_f_Int_Int_Int_Int_rbuf,MemOut_CTf_f_Int_Int_Int_Int) > (memOut_CTf_f_Int_Int_Int_Int_dbuf,MemOut_CTf_f_Int_Int_Int_Int) */
  assign memOut_CTf_f_Int_Int_Int_Int_rbuf_r = ((! memOut_CTf_f_Int_Int_Int_Int_dbuf_d[0]) || memOut_CTf_f_Int_Int_Int_Int_dbuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTf_f_Int_Int_Int_Int_dbuf_d <= {84'd0, 1'd0};
    else
      if (memOut_CTf_f_Int_Int_Int_Int_rbuf_r)
        memOut_CTf_f_Int_Int_Int_Int_dbuf_d <= memOut_CTf_f_Int_Int_Int_Int_rbuf_d;
  
  /* rbuf (Ty MemOut_CTf_f_Int_Int_Int_Int) : (memOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int) > (memOut_CTf_f_Int_Int_Int_Int_rbuf,MemOut_CTf_f_Int_Int_Int_Int) */
  MemOut_CTf_f_Int_Int_Int_Int_t memOut_CTf_f_Int_Int_Int_Int_buf;
  assign memOut_CTf_f_Int_Int_Int_Int_r = (! memOut_CTf_f_Int_Int_Int_Int_buf[0]);
  assign memOut_CTf_f_Int_Int_Int_Int_rbuf_d = (memOut_CTf_f_Int_Int_Int_Int_buf[0] ? memOut_CTf_f_Int_Int_Int_Int_buf :
                                                memOut_CTf_f_Int_Int_Int_Int_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      memOut_CTf_f_Int_Int_Int_Int_buf <= {84'd0, 1'd0};
    else
      if ((memOut_CTf_f_Int_Int_Int_Int_rbuf_r && memOut_CTf_f_Int_Int_Int_Int_buf[0]))
        memOut_CTf_f_Int_Int_Int_Int_buf <= {84'd0, 1'd0};
      else if (((! memOut_CTf_f_Int_Int_Int_Int_rbuf_r) && (! memOut_CTf_f_Int_Int_Int_Int_buf[0])))
        memOut_CTf_f_Int_Int_Int_Int_buf <= memOut_CTf_f_Int_Int_Int_Int_d;
  
  /* destruct (Ty Pointer_CTf_f_Int_Int_Int_Int,
          Dcon Pointer_CTf_f_Int_Int_Int_Int) : (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > [(destructReadIn_CTf_f_Int_Int_Int_Int,Word16#)] */
  assign destructReadIn_CTf_f_Int_Int_Int_Int_d = {scfarg_0_2_1_argbuf_d[16:1],
                                                   scfarg_0_2_1_argbuf_d[0]};
  assign scfarg_0_2_1_argbuf_r = destructReadIn_CTf_f_Int_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int_Int_Int_Int,
      Dcon ReadIn_CTf_f_Int_Int_Int_Int) : [(destructReadIn_CTf_f_Int_Int_Int_Int,Word16#)] > (dconReadIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int) */
  assign dconReadIn_CTf_f_Int_Int_Int_Int_d = ReadIn_CTf_f_Int_Int_Int_Int_dc((& {destructReadIn_CTf_f_Int_Int_Int_Int_d[0]}), destructReadIn_CTf_f_Int_Int_Int_Int_d);
  assign {destructReadIn_CTf_f_Int_Int_Int_Int_r} = {1 {(dconReadIn_CTf_f_Int_Int_Int_Int_r && dconReadIn_CTf_f_Int_Int_Int_Int_d[0])}};
  
  /* destruct (Ty MemOut_CTf_f_Int_Int_Int_Int,
          Dcon ReadOut_CTf_f_Int_Int_Int_Int) : (memReadOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int) > [(readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf,CTf_f_Int_Int_Int_Int)] */
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_d = {memReadOut_CTf_f_Int_Int_Int_Int_d[84:2],
                                                                   memReadOut_CTf_f_Int_Int_Int_Int_d[0]};
  assign memReadOut_CTf_f_Int_Int_Int_Int_r = readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_r;
  
  /* mergectrl (Ty C5,
           Ty CTf_f_Int_Int_Int_Int) : [(lizzieLet15_1_argbuf,CTf_f_Int_Int_Int_Int),
                                        (lizzieLet18_1_argbuf,CTf_f_Int_Int_Int_Int),
                                        (lizzieLet29_1_argbuf,CTf_f_Int_Int_Int_Int),
                                        (lizzieLet30_1_argbuf,CTf_f_Int_Int_Int_Int),
                                        (lizzieLet31_1_argbuf,CTf_f_Int_Int_Int_Int)] > (writeMerge_choice_CTf_f_Int_Int_Int_Int,C5) (writeMerge_data_CTf_f_Int_Int_Int_Int,CTf_f_Int_Int_Int_Int) */
  logic [4:0] lizzieLet15_1_argbuf_select_d;
  assign lizzieLet15_1_argbuf_select_d = ((| lizzieLet15_1_argbuf_select_q) ? lizzieLet15_1_argbuf_select_q :
                                          (lizzieLet15_1_argbuf_d[0] ? 5'd1 :
                                           (lizzieLet18_1_argbuf_d[0] ? 5'd2 :
                                            (lizzieLet29_1_argbuf_d[0] ? 5'd4 :
                                             (lizzieLet30_1_argbuf_d[0] ? 5'd8 :
                                              (lizzieLet31_1_argbuf_d[0] ? 5'd16 :
                                               5'd0))))));
  logic [4:0] lizzieLet15_1_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_argbuf_select_q <= 5'd0;
    else
      lizzieLet15_1_argbuf_select_q <= (lizzieLet15_1_argbuf_done ? 5'd0 :
                                        lizzieLet15_1_argbuf_select_d);
  logic [1:0] lizzieLet15_1_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet15_1_argbuf_emit_q <= 2'd0;
    else
      lizzieLet15_1_argbuf_emit_q <= (lizzieLet15_1_argbuf_done ? 2'd0 :
                                      lizzieLet15_1_argbuf_emit_d);
  logic [1:0] lizzieLet15_1_argbuf_emit_d;
  assign lizzieLet15_1_argbuf_emit_d = (lizzieLet15_1_argbuf_emit_q | ({writeMerge_choice_CTf_f_Int_Int_Int_Int_d[0],
                                                                        writeMerge_data_CTf_f_Int_Int_Int_Int_d[0]} & {writeMerge_choice_CTf_f_Int_Int_Int_Int_r,
                                                                                                                       writeMerge_data_CTf_f_Int_Int_Int_Int_r}));
  logic lizzieLet15_1_argbuf_done;
  assign lizzieLet15_1_argbuf_done = (& lizzieLet15_1_argbuf_emit_d);
  assign {lizzieLet31_1_argbuf_r,
          lizzieLet30_1_argbuf_r,
          lizzieLet29_1_argbuf_r,
          lizzieLet18_1_argbuf_r,
          lizzieLet15_1_argbuf_r} = (lizzieLet15_1_argbuf_done ? lizzieLet15_1_argbuf_select_d :
                                     5'd0);
  assign writeMerge_data_CTf_f_Int_Int_Int_Int_d = ((lizzieLet15_1_argbuf_select_d[0] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet15_1_argbuf_d :
                                                    ((lizzieLet15_1_argbuf_select_d[1] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet18_1_argbuf_d :
                                                     ((lizzieLet15_1_argbuf_select_d[2] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet29_1_argbuf_d :
                                                      ((lizzieLet15_1_argbuf_select_d[3] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet30_1_argbuf_d :
                                                       ((lizzieLet15_1_argbuf_select_d[4] && (! lizzieLet15_1_argbuf_emit_q[0])) ? lizzieLet31_1_argbuf_d :
                                                        {83'd0, 1'd0})))));
  assign writeMerge_choice_CTf_f_Int_Int_Int_Int_d = ((lizzieLet15_1_argbuf_select_d[0] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C1_5_dc(1'd1) :
                                                      ((lizzieLet15_1_argbuf_select_d[1] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C2_5_dc(1'd1) :
                                                       ((lizzieLet15_1_argbuf_select_d[2] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C3_5_dc(1'd1) :
                                                        ((lizzieLet15_1_argbuf_select_d[3] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C4_5_dc(1'd1) :
                                                         ((lizzieLet15_1_argbuf_select_d[4] && (! lizzieLet15_1_argbuf_emit_q[1])) ? C5_5_dc(1'd1) :
                                                          {3'd0, 1'd0})))));
  
  /* demux (Ty C5,
       Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeMerge_choice_CTf_f_Int_Int_Int_Int,C5) (demuxWriteResult_CTf_f_Int_Int_Int_Int,Pointer_CTf_f_Int_Int_Int_Int) > [(writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                                                                  (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                                                                  (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                                                                  (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                                                                  (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int)] */
  logic [4:0] demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd;
  always_comb
    if ((writeMerge_choice_CTf_f_Int_Int_Int_Int_d[0] && demuxWriteResult_CTf_f_Int_Int_Int_Int_d[0]))
      unique case (writeMerge_choice_CTf_f_Int_Int_Int_Int_d[3:1])
        3'd0: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd1;
        3'd1: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd2;
        3'd2: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd4;
        3'd3: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd8;
        3'd4: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd16;
        default: demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd0;
      endcase
    else demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd = 5'd0;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_Int_Int_d[16:1],
                                                             demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd[0]};
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_Int_Int_d[16:1],
                                                             demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd[1]};
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_Int_Int_d[16:1],
                                                             demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd[2]};
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_Int_Int_d[16:1],
                                                             demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd[3]};
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_d = {demuxWriteResult_CTf_f_Int_Int_Int_Int_d[16:1],
                                                             demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd[4]};
  assign demuxWriteResult_CTf_f_Int_Int_Int_Int_r = (| (demuxWriteResult_CTf_f_Int_Int_Int_Int_onehotd & {writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_r,
                                                                                                          writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_r,
                                                                                                          writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_r,
                                                                                                          writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_r,
                                                                                                          writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_r}));
  assign writeMerge_choice_CTf_f_Int_Int_Int_Int_r = demuxWriteResult_CTf_f_Int_Int_Int_Int_r;
  
  /* dcon (Ty MemIn_CTf_f_Int_Int_Int_Int,
      Dcon WriteIn_CTf_f_Int_Int_Int_Int) : [(forkHP1_CTf_f_Int_Int_Int_In2,Word16#),
                                             (writeMerge_data_CTf_f_Int_Int_Int_Int,CTf_f_Int_Int_Int_Int)] > (dconWriteIn_CTf_f_Int_Int_Int_Int,MemIn_CTf_f_Int_Int_Int_Int) */
  assign dconWriteIn_CTf_f_Int_Int_Int_Int_d = WriteIn_CTf_f_Int_Int_Int_Int_dc((& {forkHP1_CTf_f_Int_Int_Int_In2_d[0],
                                                                                    writeMerge_data_CTf_f_Int_Int_Int_Int_d[0]}), forkHP1_CTf_f_Int_Int_Int_In2_d, writeMerge_data_CTf_f_Int_Int_Int_Int_d);
  assign {forkHP1_CTf_f_Int_Int_Int_In2_r,
          writeMerge_data_CTf_f_Int_Int_Int_Int_r} = {2 {(dconWriteIn_CTf_f_Int_Int_Int_Int_r && dconWriteIn_CTf_f_Int_Int_Int_Int_d[0])}};
  
  /* dcon (Ty Pointer_CTf_f_Int_Int_Int_Int,
      Dcon Pointer_CTf_f_Int_Int_Int_Int) : [(forkHP1_CTf_f_Int_Int_Int_In3,Word16#)] > (dconPtr_CTf_f_Int_Int_Int_Int,Pointer_CTf_f_Int_Int_Int_Int) */
  assign dconPtr_CTf_f_Int_Int_Int_Int_d = Pointer_CTf_f_Int_Int_Int_Int_dc((& {forkHP1_CTf_f_Int_Int_Int_In3_d[0]}), forkHP1_CTf_f_Int_Int_Int_In3_d);
  assign {forkHP1_CTf_f_Int_Int_Int_In3_r} = {1 {(dconPtr_CTf_f_Int_Int_Int_Int_r && dconPtr_CTf_f_Int_Int_Int_Int_d[0])}};
  
  /* demux (Ty MemOut_CTf_f_Int_Int_Int_Int,
       Ty Pointer_CTf_f_Int_Int_Int_Int) : (memWriteOut_CTf_f_Int_Int_Int_Int,MemOut_CTf_f_Int_Int_Int_Int) (dconPtr_CTf_f_Int_Int_Int_Int,Pointer_CTf_f_Int_Int_Int_Int) > [(_42,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                                                                             (demuxWriteResult_CTf_f_Int_Int_Int_Int,Pointer_CTf_f_Int_Int_Int_Int)] */
  logic [1:0] dconPtr_CTf_f_Int_Int_Int_Int_onehotd;
  always_comb
    if ((memWriteOut_CTf_f_Int_Int_Int_Int_d[0] && dconPtr_CTf_f_Int_Int_Int_Int_d[0]))
      unique case (memWriteOut_CTf_f_Int_Int_Int_Int_d[1:1])
        1'd0: dconPtr_CTf_f_Int_Int_Int_Int_onehotd = 2'd1;
        1'd1: dconPtr_CTf_f_Int_Int_Int_Int_onehotd = 2'd2;
        default: dconPtr_CTf_f_Int_Int_Int_Int_onehotd = 2'd0;
      endcase
    else dconPtr_CTf_f_Int_Int_Int_Int_onehotd = 2'd0;
  assign _42_d = {dconPtr_CTf_f_Int_Int_Int_Int_d[16:1],
                  dconPtr_CTf_f_Int_Int_Int_Int_onehotd[0]};
  assign demuxWriteResult_CTf_f_Int_Int_Int_Int_d = {dconPtr_CTf_f_Int_Int_Int_Int_d[16:1],
                                                     dconPtr_CTf_f_Int_Int_Int_Int_onehotd[1]};
  assign dconPtr_CTf_f_Int_Int_Int_Int_r = (| (dconPtr_CTf_f_Int_Int_Int_Int_onehotd & {demuxWriteResult_CTf_f_Int_Int_Int_Int_r,
                                                                                        _42_r}));
  assign memWriteOut_CTf_f_Int_Int_Int_Int_r = dconPtr_CTf_f_Int_Int_Int_Int_r;
  
  /* source (Ty Go) : > (sourceGo,Go) */
  
  /* source (Ty Pointer_QTree_Int) : > (m1ahS_0,Pointer_QTree_Int) */
  
  /* source (Ty Pointer_QTree_Int) : > (m2ahT_1,Pointer_QTree_Int) */
  
  /* destruct (Ty TupGo___Pointer_QTree_Int,
          Dcon TupGo___Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) > [($wnnz_IntTupGo___Pointer_QTree_Intgo_7,Go),
                                                                                                                ($wnnz_IntTupGo___Pointer_QTree_IntwstH,Pointer_QTree_Int)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Int_1_done ;
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_d  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [0]));
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwstH_d  = {\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [16:1],
                                                       (\$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted [1]))};
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_done  = (\$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  | ({\$wnnz_IntTupGo___Pointer_QTree_IntwstH_d [0],
                                                                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_d [0]} & {\$wnnz_IntTupGo___Pointer_QTree_IntwstH_r ,
                                                                                                                                                             \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_r }));
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Int_1_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  ? 2'd0 :
                                                         \$wnnz_IntTupGo___Pointer_QTree_Int_1_done );
  
  /* fork (Ty Go) : ($wnnz_IntTupGo___Pointer_QTree_Intgo_7,Go) > [(go_7_1,Go),
                                                              (go_7_2,Go)] */
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted ;
  logic [1:0] \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_done ;
  assign go_7_1_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_7_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted [0]));
  assign go_7_2_d = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_7_d [0] && (! \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted [1]));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_done  = (\$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted  | ({go_7_2_d[0],
                                                                                                               go_7_1_d[0]} & {go_7_2_r,
                                                                                                                               go_7_1_r}));
  assign \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_r  = (& \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted  <= 2'd0;
    else
      \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_emitted  <= (\$wnnz_IntTupGo___Pointer_QTree_Intgo_7_r  ? 2'd0 :
                                                           \$wnnz_IntTupGo___Pointer_QTree_Intgo_7_done );
  
  /* buf (Ty Pointer_QTree_Int) : ($wnnz_IntTupGo___Pointer_QTree_IntwstH,Pointer_QTree_Int) > (wstH_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d ;
  logic \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_r ;
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwstH_r  = ((! \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d [0]) || \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d  <= {16'd0,
                                                             1'd0};
    else
      if (\$wnnz_IntTupGo___Pointer_QTree_IntwstH_r )
        \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d  <= \$wnnz_IntTupGo___Pointer_QTree_IntwstH_d ;
  Pointer_QTree_Int_t \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf ;
  assign \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_r  = (! \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf [0]);
  assign wstH_1_argbuf_d = (\$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf [0] ? \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf  :
                            \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf  <= {16'd0,
                                                               1'd0};
    else
      if ((wstH_1_argbuf_r && \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf [0]))
        \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf  <= {16'd0,
                                                                 1'd0};
      else if (((! wstH_1_argbuf_r) && (! \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf [0])))
        \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_buf  <= \$wnnz_IntTupGo___Pointer_QTree_IntwstH_bufchan_d ;
  
  /* dcon (Ty Int,Dcon I#) : [($wnnz_Int_resbuf,Int#)] > (es_7_1I#,Int) */
  assign \es_7_1I#_d  = \I#_dc ((& {\$wnnz_Int_resbuf_d [0]}), \$wnnz_Int_resbuf_d );
  assign {\$wnnz_Int_resbuf_r } = {1 {(\es_7_1I#_r  && \es_7_1I#_d [0])}};
  
  /* mergectrl (Ty C2,
           Ty TupGo___MyDTInt_Bool___Int) : [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int),
                                             (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int)] > (applyfnInt_Bool_5_choice,C2) (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) */
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d = ((| applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q :
                                                                   (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0] ? 2'd1 :
                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0] ? 2'd2 :
                                                                     2'd0)));
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                                 applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? 2'd0 :
                                                               applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  logic [1:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q | ({applyfnInt_Bool_5_choice_d[0],
                                                                                                                          applyfnInt_Bool_5_data_d[0]} & {applyfnInt_Bool_5_choice_r,
                                                                                                                                                          applyfnInt_Bool_5_data_r}));
  logic applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_d);
  assign {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r,
          applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r} = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_done ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d :
                                                              2'd0);
  assign applyfnInt_Bool_5_data_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d :
                                     ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[0])) ? applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d :
                                      {32'd0, 1'd0}));
  assign applyfnInt_Bool_5_choice_d = ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C1_2_dc(1'd1) :
                                       ((applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_select_d[1] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_emit_q[1])) ? C2_2_dc(1'd1) :
                                        {1'd0, 1'd0}));
  
  /* fork (Ty MyDTInt_Bool) : (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool) > [(arg0_1,MyDTInt_Bool),
                                                                                           (arg0_2,MyDTInt_Bool),
                                                                                           (arg0_3,MyDTInt_Bool)] */
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted;
  logic [2:0] applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done;
  assign arg0_1_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[0]));
  assign arg0_2_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[1]));
  assign arg0_3_d = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0] && (! applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted[2]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done = (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted | ({arg0_3_d[0],
                                                                                                                             arg0_2_d[0],
                                                                                                                             arg0_1_d[0]} & {arg0_3_r,
                                                                                                                                             arg0_2_r,
                                                                                                                                             arg0_1_r}));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r = (& applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= 3'd0;
    else
      applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_emitted <= (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r ? 3'd0 :
                                                                  applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_done);
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_1,MyBool) > (applyfnInt_Bool_5_resbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_1_bufchan_d;
  logic applyfnInt_Bool_5_1_bufchan_r;
  assign applyfnInt_Bool_5_1_r = ((! applyfnInt_Bool_5_1_bufchan_d[0]) || applyfnInt_Bool_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_1_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_1_r)
        applyfnInt_Bool_5_1_bufchan_d <= applyfnInt_Bool_5_1_d;
  MyBool_t applyfnInt_Bool_5_1_bufchan_buf;
  assign applyfnInt_Bool_5_1_bufchan_r = (! applyfnInt_Bool_5_1_bufchan_buf[0]);
  assign applyfnInt_Bool_5_resbuf_d = (applyfnInt_Bool_5_1_bufchan_buf[0] ? applyfnInt_Bool_5_1_bufchan_buf :
                                       applyfnInt_Bool_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_resbuf_r && applyfnInt_Bool_5_1_bufchan_buf[0]))
        applyfnInt_Bool_5_1_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_resbuf_r) && (! applyfnInt_Bool_5_1_bufchan_buf[0])))
        applyfnInt_Bool_5_1_bufchan_buf <= applyfnInt_Bool_5_1_bufchan_d;
  
  /* buf (Ty MyBool) : (applyfnInt_Bool_5_2,MyBool) > (applyfnInt_Bool_5_2_argbuf,MyBool) */
  MyBool_t applyfnInt_Bool_5_2_bufchan_d;
  logic applyfnInt_Bool_5_2_bufchan_r;
  assign applyfnInt_Bool_5_2_r = ((! applyfnInt_Bool_5_2_bufchan_d[0]) || applyfnInt_Bool_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_bufchan_d <= {1'd0, 1'd0};
    else
      if (applyfnInt_Bool_5_2_r)
        applyfnInt_Bool_5_2_bufchan_d <= applyfnInt_Bool_5_2_d;
  MyBool_t applyfnInt_Bool_5_2_bufchan_buf;
  assign applyfnInt_Bool_5_2_bufchan_r = (! applyfnInt_Bool_5_2_bufchan_buf[0]);
  assign applyfnInt_Bool_5_2_argbuf_d = (applyfnInt_Bool_5_2_bufchan_buf[0] ? applyfnInt_Bool_5_2_bufchan_buf :
                                         applyfnInt_Bool_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((applyfnInt_Bool_5_2_argbuf_r && applyfnInt_Bool_5_2_bufchan_buf[0]))
        applyfnInt_Bool_5_2_bufchan_buf <= {1'd0, 1'd0};
      else if (((! applyfnInt_Bool_5_2_argbuf_r) && (! applyfnInt_Bool_5_2_bufchan_buf[0])))
        applyfnInt_Bool_5_2_bufchan_buf <= applyfnInt_Bool_5_2_bufchan_d;
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_2_argbuf,MyBool) > [(es_7_1_1,MyBool),
                                                          (es_7_1_2,MyBool),
                                                          (es_7_1_3,MyBool),
                                                          (es_7_1_4,MyBool),
                                                          (es_7_1_5,MyBool),
                                                          (es_7_1_6,MyBool)] */
  logic [5:0] applyfnInt_Bool_5_2_argbuf_emitted;
  logic [5:0] applyfnInt_Bool_5_2_argbuf_done;
  assign es_7_1_1_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[0]))};
  assign es_7_1_2_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[1]))};
  assign es_7_1_3_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[2]))};
  assign es_7_1_4_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[3]))};
  assign es_7_1_5_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[4]))};
  assign es_7_1_6_d = {applyfnInt_Bool_5_2_argbuf_d[1:1],
                       (applyfnInt_Bool_5_2_argbuf_d[0] && (! applyfnInt_Bool_5_2_argbuf_emitted[5]))};
  assign applyfnInt_Bool_5_2_argbuf_done = (applyfnInt_Bool_5_2_argbuf_emitted | ({es_7_1_6_d[0],
                                                                                   es_7_1_5_d[0],
                                                                                   es_7_1_4_d[0],
                                                                                   es_7_1_3_d[0],
                                                                                   es_7_1_2_d[0],
                                                                                   es_7_1_1_d[0]} & {es_7_1_6_r,
                                                                                                     es_7_1_5_r,
                                                                                                     es_7_1_4_r,
                                                                                                     es_7_1_3_r,
                                                                                                     es_7_1_2_r,
                                                                                                     es_7_1_1_r}));
  assign applyfnInt_Bool_5_2_argbuf_r = (& applyfnInt_Bool_5_2_argbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_2_argbuf_emitted <= 6'd0;
    else
      applyfnInt_Bool_5_2_argbuf_emitted <= (applyfnInt_Bool_5_2_argbuf_r ? 6'd0 :
                                             applyfnInt_Bool_5_2_argbuf_done);
  
  /* demux (Ty C2,
       Ty MyBool) : (applyfnInt_Bool_5_choice,C2) (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) > [(applyfnInt_Bool_5_1,MyBool),
                                                                                                                                 (applyfnInt_Bool_5_2,MyBool)] */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd;
  always_comb
    if ((applyfnInt_Bool_5_choice_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[0]))
      unique case (applyfnInt_Bool_5_choice_d[1:1])
        1'd0:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd1;
        1'd1:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd2;
        default:
          lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
      endcase
    else
      lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd = 2'd0;
  assign applyfnInt_Bool_5_1_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[0]};
  assign applyfnInt_Bool_5_2_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d[1:1],
                                  lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd[1]};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r = (| (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_onehotd & {applyfnInt_Bool_5_2_r,
                                                                                                                                                                  applyfnInt_Bool_5_1_r}));
  assign applyfnInt_Bool_5_choice_r = lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r;
  
  /* destruct (Ty TupGo___MyDTInt_Bool___Int,
          Dcon TupGo___MyDTInt_Bool___Int) : (applyfnInt_Bool_5_data,TupGo___MyDTInt_Bool___Int) > [(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8,Go),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0,MyDTInt_Bool),
                                                                                                    (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int)] */
  logic [2:0] applyfnInt_Bool_5_data_emitted;
  logic [2:0] applyfnInt_Bool_5_data_done;
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[0]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d = (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[1]));
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d = {applyfnInt_Bool_5_data_d[32:1],
                                                              (applyfnInt_Bool_5_data_d[0] && (! applyfnInt_Bool_5_data_emitted[2]))};
  assign applyfnInt_Bool_5_data_done = (applyfnInt_Bool_5_data_emitted | ({applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_d[0],
                                                                           applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]} & {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg0_r,
                                                                                                                                    applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r}));
  assign applyfnInt_Bool_5_data_r = (& applyfnInt_Bool_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_data_emitted <= 3'd0;
    else
      applyfnInt_Bool_5_data_emitted <= (applyfnInt_Bool_5_data_r ? 3'd0 :
                                         applyfnInt_Bool_5_data_done);
  
  /* fork (Ty MyBool) : (applyfnInt_Bool_5_resbuf,MyBool) > [(es_2_1,MyBool),
                                                        (es_2_2,MyBool),
                                                        (es_2_3,MyBool),
                                                        (es_2_4,MyBool),
                                                        (es_2_5,MyBool),
                                                        (es_2_6,MyBool),
                                                        (es_2_7,MyBool)] */
  logic [6:0] applyfnInt_Bool_5_resbuf_emitted;
  logic [6:0] applyfnInt_Bool_5_resbuf_done;
  assign es_2_1_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[0]))};
  assign es_2_2_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[1]))};
  assign es_2_3_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[2]))};
  assign es_2_4_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[3]))};
  assign es_2_5_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[4]))};
  assign es_2_6_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[5]))};
  assign es_2_7_d = {applyfnInt_Bool_5_resbuf_d[1:1],
                     (applyfnInt_Bool_5_resbuf_d[0] && (! applyfnInt_Bool_5_resbuf_emitted[6]))};
  assign applyfnInt_Bool_5_resbuf_done = (applyfnInt_Bool_5_resbuf_emitted | ({es_2_7_d[0],
                                                                               es_2_6_d[0],
                                                                               es_2_5_d[0],
                                                                               es_2_4_d[0],
                                                                               es_2_3_d[0],
                                                                               es_2_2_d[0],
                                                                               es_2_1_d[0]} & {es_2_7_r,
                                                                                               es_2_6_r,
                                                                                               es_2_5_r,
                                                                                               es_2_4_r,
                                                                                               es_2_3_r,
                                                                                               es_2_2_r,
                                                                                               es_2_1_r}));
  assign applyfnInt_Bool_5_resbuf_r = (& applyfnInt_Bool_5_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Bool_5_resbuf_emitted <= 7'd0;
    else
      applyfnInt_Bool_5_resbuf_emitted <= (applyfnInt_Bool_5_resbuf_r ? 7'd0 :
                                           applyfnInt_Bool_5_resbuf_done);
  
  /* mergectrl (Ty C2,
           Ty TupGo___MyDTInt_Int___Int) : [(applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int),
                                            (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2,TupGo___MyDTInt_Int___Int)] > (applyfnInt_Int_5_choice,C2) (applyfnInt_Int_5_data,TupGo___MyDTInt_Int___Int) */
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d = ((| applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q :
                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0] ? 2'd1 :
                                                                  (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d[0] ? 2'd2 :
                                                                   2'd0)));
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q <= 2'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_q <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? 2'd0 :
                                                               applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? 2'd0 :
                                                             applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q | ({applyfnInt_Int_5_choice_d[0],
                                                                                                                      applyfnInt_Int_5_data_d[0]} & {applyfnInt_Int_5_choice_r,
                                                                                                                                                     applyfnInt_Int_5_data_r}));
  logic applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_d);
  assign {applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r,
          applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r} = (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_done ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d :
                                                            2'd0);
  assign applyfnInt_Int_5_data_d = ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d :
                                    ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[1] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[0])) ? applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d :
                                     {32'd0, 1'd0}));
  assign applyfnInt_Int_5_choice_d = ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C1_2_dc(1'd1) :
                                      ((applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_select_d[1] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_emit_q[1])) ? C2_2_dc(1'd1) :
                                       {1'd0, 1'd0}));
  
  /* fork (Ty MyDTInt_Int) : (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int) > [(arg0_2_1,MyDTInt_Int),
                                                                                         (arg0_2_2,MyDTInt_Int),
                                                                                         (arg0_2_3,MyDTInt_Int)] */
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted;
  logic [2:0] applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done;
  assign arg0_2_1_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[0]));
  assign arg0_2_2_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[1]));
  assign arg0_2_3_d = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0] && (! applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted[2]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done = (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted | ({arg0_2_3_d[0],
                                                                                                                             arg0_2_2_d[0],
                                                                                                                             arg0_2_1_d[0]} & {arg0_2_3_r,
                                                                                                                                               arg0_2_2_r,
                                                                                                                                               arg0_2_1_r}));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r = (& applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= 3'd0;
    else
      applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_emitted <= (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r ? 3'd0 :
                                                                  applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_5_1,Int) > (applyfnInt_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_5_1_bufchan_d;
  logic applyfnInt_Int_5_1_bufchan_r;
  assign applyfnInt_Int_5_1_r = ((! applyfnInt_Int_5_1_bufchan_d[0]) || applyfnInt_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_1_r)
        applyfnInt_Int_5_1_bufchan_d <= applyfnInt_Int_5_1_d;
  Int_t applyfnInt_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_5_1_bufchan_r = (! applyfnInt_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_5_resbuf_d = (applyfnInt_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_5_1_bufchan_buf :
                                      applyfnInt_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_resbuf_r && applyfnInt_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_resbuf_r) && (! applyfnInt_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_5_1_bufchan_buf <= applyfnInt_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_5_2,Int) > (applyfnInt_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_5_2_bufchan_d;
  logic applyfnInt_Int_5_2_bufchan_r;
  assign applyfnInt_Int_5_2_r = ((! applyfnInt_Int_5_2_bufchan_d[0]) || applyfnInt_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_2_r)
        applyfnInt_Int_5_2_bufchan_d <= applyfnInt_Int_5_2_d;
  Int_t applyfnInt_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_5_2_bufchan_r = (! applyfnInt_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_5_2_argbuf_d = (applyfnInt_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_5_2_bufchan_buf :
                                        applyfnInt_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_5_2_argbuf_r && applyfnInt_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_5_2_argbuf_r) && (! applyfnInt_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_5_2_bufchan_buf <= applyfnInt_Int_5_2_bufchan_d;
  
  /* dcon (Ty QTree_Int,
      Dcon QVal_Int) : [(applyfnInt_Int_5_2_argbuf,Int)] > (es_8_1QVal_Int,QTree_Int) */
  assign es_8_1QVal_Int_d = QVal_Int_dc((& {applyfnInt_Int_5_2_argbuf_d[0]}), applyfnInt_Int_5_2_argbuf_d);
  assign {applyfnInt_Int_5_2_argbuf_r} = {1 {(es_8_1QVal_Int_r && es_8_1QVal_Int_d[0])}};
  
  /* demux (Ty C2,
       Ty Int) : (applyfnInt_Int_5_choice,C2) (es_0_1_1I#_mux_mux,Int) > [(applyfnInt_Int_5_1,Int),
                                                                          (applyfnInt_Int_5_2,Int)] */
  logic [1:0] \es_0_1_1I#_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_5_choice_d[0] && \es_0_1_1I#_mux_mux_d [0]))
      unique case (applyfnInt_Int_5_choice_d[1:1])
        1'd0: \es_0_1_1I#_mux_mux_onehotd  = 2'd1;
        1'd1: \es_0_1_1I#_mux_mux_onehotd  = 2'd2;
        default: \es_0_1_1I#_mux_mux_onehotd  = 2'd0;
      endcase
    else \es_0_1_1I#_mux_mux_onehotd  = 2'd0;
  assign applyfnInt_Int_5_1_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [0]};
  assign applyfnInt_Int_5_2_d = {\es_0_1_1I#_mux_mux_d [32:1],
                                 \es_0_1_1I#_mux_mux_onehotd [1]};
  assign \es_0_1_1I#_mux_mux_r  = (| (\es_0_1_1I#_mux_mux_onehotd  & {applyfnInt_Int_5_2_r,
                                                                      applyfnInt_Int_5_1_r}));
  assign applyfnInt_Int_5_choice_r = \es_0_1_1I#_mux_mux_r ;
  
  /* destruct (Ty TupGo___MyDTInt_Int___Int,
          Dcon TupGo___MyDTInt_Int___Int) : (applyfnInt_Int_5_data,TupGo___MyDTInt_Int___Int) > [(applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9,Go),
                                                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2,MyDTInt_Int),
                                                                                                 (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int)] */
  logic [2:0] applyfnInt_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_5_data_done;
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d = (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[0]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d = (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[1]));
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d = {applyfnInt_Int_5_data_d[32:1],
                                                              (applyfnInt_Int_5_data_d[0] && (! applyfnInt_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_5_data_done = (applyfnInt_Int_5_data_emitted | ({applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0],
                                                                         applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_d[0],
                                                                         applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]} & {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r,
                                                                                                                                applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg0_2_r,
                                                                                                                                applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r}));
  assign applyfnInt_Int_5_data_r = (& applyfnInt_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_5_data_emitted <= (applyfnInt_Int_5_data_r ? 3'd0 :
                                        applyfnInt_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_5_resbuf,Int) > (es_4_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_5_resbuf_r = ((! applyfnInt_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_5_resbuf_r)
        applyfnInt_Int_5_resbuf_bufchan_d <= applyfnInt_Int_5_resbuf_d;
  Int_t applyfnInt_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_5_resbuf_bufchan_buf[0]);
  assign es_4_1_1_argbuf_d = (applyfnInt_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_5_resbuf_bufchan_buf :
                              applyfnInt_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_4_1_1_argbuf_r && applyfnInt_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_4_1_1_argbuf_r) && (! applyfnInt_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_5_resbuf_bufchan_d;
  
  /* mergectrl (Ty C3,
           Ty TupMyDTInt_Int_Int___Int___Int) : [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int),
                                                 (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int)] > (applyfnInt_Int_Int_5_choice,C3) (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d = ((| applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q :
                                                                          (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0] ? 3'd1 :
                                                                           (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0] ? 3'd2 :
                                                                            (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0] ? 3'd4 :
                                                                             3'd0))));
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 3'd0 :
                                                                        applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= 2'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? 2'd0 :
                                                                      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  logic [1:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q | ({applyfnInt_Int_Int_5_choice_d[0],
                                                                                                                                        applyfnInt_Int_Int_5_data_d[0]} & {applyfnInt_Int_Int_5_choice_r,
                                                                                                                                                                           applyfnInt_Int_Int_5_data_r}));
  logic applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_d);
  assign {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r,
          applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r} = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_done ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d :
                                                                     3'd0);
  assign applyfnInt_Int_Int_5_data_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d :
                                        ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d :
                                         ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[0])) ? applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d :
                                          {64'd0, 1'd0})));
  assign applyfnInt_Int_Int_5_choice_d = ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C1_3_dc(1'd1) :
                                          ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[1] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C2_3_dc(1'd1) :
                                           ((applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_select_d[2] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_emit_q[1])) ? C3_3_dc(1'd1) :
                                            {2'd0, 1'd0})));
  
  /* fork (Ty MyDTInt_Int_Int) : (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int) > [(arg0_4_1,MyDTInt_Int_Int),
                                                                                                          (arg0_4_2,MyDTInt_Int_Int),
                                                                                                          (arg0_4_3,MyDTInt_Int_Int)] */
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted;
  logic [2:0] applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done;
  assign arg0_4_1_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[0]));
  assign arg0_4_2_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[1]));
  assign arg0_4_3_d = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0] && (! applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted[2]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done = (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted | ({arg0_4_3_d[0],
                                                                                                                                               arg0_4_2_d[0],
                                                                                                                                               arg0_4_1_d[0]} & {arg0_4_3_r,
                                                                                                                                                                 arg0_4_2_r,
                                                                                                                                                                 arg0_4_1_r}));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r = (& applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_emitted <= (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r ? 3'd0 :
                                                                           applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_1,Int) > (applyfnInt_Int_Int_5_resbuf,Int) */
  Int_t applyfnInt_Int_Int_5_1_bufchan_d;
  logic applyfnInt_Int_Int_5_1_bufchan_r;
  assign applyfnInt_Int_Int_5_1_r = ((! applyfnInt_Int_Int_5_1_bufchan_d[0]) || applyfnInt_Int_Int_5_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_1_r)
        applyfnInt_Int_Int_5_1_bufchan_d <= applyfnInt_Int_Int_5_1_d;
  Int_t applyfnInt_Int_Int_5_1_bufchan_buf;
  assign applyfnInt_Int_Int_5_1_bufchan_r = (! applyfnInt_Int_Int_5_1_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_resbuf_d = (applyfnInt_Int_Int_5_1_bufchan_buf[0] ? applyfnInt_Int_Int_5_1_bufchan_buf :
                                          applyfnInt_Int_Int_5_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_resbuf_r && applyfnInt_Int_Int_5_1_bufchan_buf[0]))
        applyfnInt_Int_Int_5_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_resbuf_r) && (! applyfnInt_Int_Int_5_1_bufchan_buf[0])))
        applyfnInt_Int_Int_5_1_bufchan_buf <= applyfnInt_Int_Int_5_1_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2,Int) > (applyfnInt_Int_Int_5_2_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_bufchan_d;
  logic applyfnInt_Int_Int_5_2_bufchan_r;
  assign applyfnInt_Int_Int_5_2_r = ((! applyfnInt_Int_Int_5_2_bufchan_d[0]) || applyfnInt_Int_Int_5_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_r)
        applyfnInt_Int_Int_5_2_bufchan_d <= applyfnInt_Int_Int_5_2_d;
  Int_t applyfnInt_Int_Int_5_2_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_bufchan_r = (! applyfnInt_Int_Int_5_2_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_2_argbuf_d = (applyfnInt_Int_Int_5_2_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_bufchan_buf :
                                            applyfnInt_Int_Int_5_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_2_argbuf_r && applyfnInt_Int_Int_5_2_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_2_argbuf_r) && (! applyfnInt_Int_Int_5_2_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_bufchan_buf <= applyfnInt_Int_Int_5_2_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_2_argbuf,Int) > (es_6_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_2_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_2_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_2_argbuf_r = ((! applyfnInt_Int_Int_5_2_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_2_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_2_argbuf_r)
        applyfnInt_Int_Int_5_2_argbuf_bufchan_d <= applyfnInt_Int_Int_5_2_argbuf_d;
  Int_t applyfnInt_Int_Int_5_2_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_2_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0]);
  assign es_6_1_1_argbuf_d = (applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_2_argbuf_bufchan_buf :
                              applyfnInt_Int_Int_5_2_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_6_1_1_argbuf_r && applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_6_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_2_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_2_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_2_argbuf_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3,Int) > (applyfnInt_Int_Int_5_3_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_bufchan_d;
  logic applyfnInt_Int_Int_5_3_bufchan_r;
  assign applyfnInt_Int_Int_5_3_r = ((! applyfnInt_Int_Int_5_3_bufchan_d[0]) || applyfnInt_Int_Int_5_3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_r)
        applyfnInt_Int_Int_5_3_bufchan_d <= applyfnInt_Int_Int_5_3_d;
  Int_t applyfnInt_Int_Int_5_3_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_bufchan_r = (! applyfnInt_Int_Int_5_3_bufchan_buf[0]);
  assign applyfnInt_Int_Int_5_3_argbuf_d = (applyfnInt_Int_Int_5_3_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_bufchan_buf :
                                            applyfnInt_Int_Int_5_3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((applyfnInt_Int_Int_5_3_argbuf_r && applyfnInt_Int_Int_5_3_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_bufchan_buf <= {32'd0, 1'd0};
      else if (((! applyfnInt_Int_Int_5_3_argbuf_r) && (! applyfnInt_Int_Int_5_3_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_bufchan_buf <= applyfnInt_Int_Int_5_3_bufchan_d;
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_3_argbuf,Int) > (es_10_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_3_argbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_3_argbuf_r = ((! applyfnInt_Int_Int_5_3_argbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_3_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_3_argbuf_r)
        applyfnInt_Int_Int_5_3_argbuf_bufchan_d <= applyfnInt_Int_Int_5_3_argbuf_d;
  Int_t applyfnInt_Int_Int_5_3_argbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_3_argbuf_bufchan_r = (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]);
  assign es_10_1_argbuf_d = (applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_3_argbuf_bufchan_buf :
                             applyfnInt_Int_Int_5_3_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_10_1_argbuf_r && applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_10_1_argbuf_r) && (! applyfnInt_Int_Int_5_3_argbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_3_argbuf_bufchan_buf <= applyfnInt_Int_Int_5_3_argbuf_bufchan_d;
  
  /* demux (Ty C3,
       Ty Int) : (applyfnInt_Int_Int_5_choice,C3) (es_0_2_1I#_mux_mux_mux,Int) > [(applyfnInt_Int_Int_5_1,Int),
                                                                                  (applyfnInt_Int_Int_5_2,Int),
                                                                                  (applyfnInt_Int_Int_5_3,Int)] */
  logic [2:0] \es_0_2_1I#_mux_mux_mux_onehotd ;
  always_comb
    if ((applyfnInt_Int_Int_5_choice_d[0] && \es_0_2_1I#_mux_mux_mux_d [0]))
      unique case (applyfnInt_Int_Int_5_choice_d[2:1])
        2'd0: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd1;
        2'd1: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd2;
        2'd2: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd4;
        default: \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd0;
      endcase
    else \es_0_2_1I#_mux_mux_mux_onehotd  = 3'd0;
  assign applyfnInt_Int_Int_5_1_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [0]};
  assign applyfnInt_Int_Int_5_2_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [1]};
  assign applyfnInt_Int_Int_5_3_d = {\es_0_2_1I#_mux_mux_mux_d [32:1],
                                     \es_0_2_1I#_mux_mux_mux_onehotd [2]};
  assign \es_0_2_1I#_mux_mux_mux_r  = (| (\es_0_2_1I#_mux_mux_mux_onehotd  & {applyfnInt_Int_Int_5_3_r,
                                                                              applyfnInt_Int_Int_5_2_r,
                                                                              applyfnInt_Int_Int_5_1_r}));
  assign applyfnInt_Int_Int_5_choice_r = \es_0_2_1I#_mux_mux_mux_r ;
  
  /* destruct (Ty TupMyDTInt_Int_Int___Int___Int,
          Dcon TupMyDTInt_Int_Int___Int___Int) : (applyfnInt_Int_Int_5_data,TupMyDTInt_Int_Int___Int___Int) > [(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4,MyDTInt_Int_Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int),
                                                                                                               (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int)] */
  logic [2:0] applyfnInt_Int_Int_5_data_emitted;
  logic [2:0] applyfnInt_Int_Int_5_data_done;
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d = (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[0]));
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d = {applyfnInt_Int_Int_5_data_d[32:1],
                                                                     (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[1]))};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d = {applyfnInt_Int_Int_5_data_d[64:33],
                                                                       (applyfnInt_Int_Int_5_data_d[0] && (! applyfnInt_Int_Int_5_data_emitted[2]))};
  assign applyfnInt_Int_Int_5_data_done = (applyfnInt_Int_Int_5_data_emitted | ({applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0],
                                                                                 applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_d[0]} & {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r,
                                                                                                                                                   applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg0_4_r}));
  assign applyfnInt_Int_Int_5_data_r = (& applyfnInt_Int_Int_5_data_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) applyfnInt_Int_Int_5_data_emitted <= 3'd0;
    else
      applyfnInt_Int_Int_5_data_emitted <= (applyfnInt_Int_Int_5_data_r ? 3'd0 :
                                            applyfnInt_Int_Int_5_data_done);
  
  /* buf (Ty Int) : (applyfnInt_Int_Int_5_resbuf,Int) > (es_1_1_argbuf,Int) */
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_d;
  logic applyfnInt_Int_Int_5_resbuf_bufchan_r;
  assign applyfnInt_Int_Int_5_resbuf_r = ((! applyfnInt_Int_Int_5_resbuf_bufchan_d[0]) || applyfnInt_Int_Int_5_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_d <= {32'd0, 1'd0};
    else
      if (applyfnInt_Int_Int_5_resbuf_r)
        applyfnInt_Int_Int_5_resbuf_bufchan_d <= applyfnInt_Int_Int_5_resbuf_d;
  Int_t applyfnInt_Int_Int_5_resbuf_bufchan_buf;
  assign applyfnInt_Int_Int_5_resbuf_bufchan_r = (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]);
  assign es_1_1_argbuf_d = (applyfnInt_Int_Int_5_resbuf_bufchan_buf[0] ? applyfnInt_Int_Int_5_resbuf_bufchan_buf :
                            applyfnInt_Int_Int_5_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_1_1_argbuf_r && applyfnInt_Int_Int_5_resbuf_bufchan_buf[0]))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_1_1_argbuf_r) && (! applyfnInt_Int_Int_5_resbuf_bufchan_buf[0])))
        applyfnInt_Int_Int_5_resbuf_bufchan_buf <= applyfnInt_Int_Int_5_resbuf_bufchan_d;
  
  /* demux (Ty MyDTInt_Bool,
       Ty Int) : (arg0_1,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1,Int) > [(arg0_1Dcon_eqZero,Int)] */
  assign arg0_1Dcon_eqZero_d = {applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[32:1],
                                (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0])};
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_r = (arg0_1Dcon_eqZero_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  assign arg0_1_r = (arg0_1Dcon_eqZero_r && (arg0_1_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intarg1_d[0]));
  
  /* fork (Ty Int) : (arg0_1Dcon_eqZero,Int) > [(arg0_1Dcon_eqZero_1,Int),
                                           (arg0_1Dcon_eqZero_2,Int),
                                           (arg0_1Dcon_eqZero_3,Int),
                                           (arg0_1Dcon_eqZero_4,Int)] */
  logic [3:0] arg0_1Dcon_eqZero_emitted;
  logic [3:0] arg0_1Dcon_eqZero_done;
  assign arg0_1Dcon_eqZero_1_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[0]))};
  assign arg0_1Dcon_eqZero_2_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[1]))};
  assign arg0_1Dcon_eqZero_3_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[2]))};
  assign arg0_1Dcon_eqZero_4_d = {arg0_1Dcon_eqZero_d[32:1],
                                  (arg0_1Dcon_eqZero_d[0] && (! arg0_1Dcon_eqZero_emitted[3]))};
  assign arg0_1Dcon_eqZero_done = (arg0_1Dcon_eqZero_emitted | ({arg0_1Dcon_eqZero_4_d[0],
                                                                 arg0_1Dcon_eqZero_3_d[0],
                                                                 arg0_1Dcon_eqZero_2_d[0],
                                                                 arg0_1Dcon_eqZero_1_d[0]} & {arg0_1Dcon_eqZero_4_r,
                                                                                              arg0_1Dcon_eqZero_3_r,
                                                                                              arg0_1Dcon_eqZero_2_r,
                                                                                              arg0_1Dcon_eqZero_1_r}));
  assign arg0_1Dcon_eqZero_r = (& arg0_1Dcon_eqZero_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_1Dcon_eqZero_emitted <= 4'd0;
    else
      arg0_1Dcon_eqZero_emitted <= (arg0_1Dcon_eqZero_r ? 4'd0 :
                                    arg0_1Dcon_eqZero_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_1Dcon_eqZero_1I#,Int) > [(x1aph_destruct,Int#)] */
  assign x1aph_destruct_d = {\arg0_1Dcon_eqZero_1I#_d [32:1],
                             \arg0_1Dcon_eqZero_1I#_d [0]};
  assign \arg0_1Dcon_eqZero_1I#_r  = x1aph_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_1Dcon_eqZero_2,Int) (arg0_1Dcon_eqZero_1,Int) > [(arg0_1Dcon_eqZero_1I#,Int)] */
  assign \arg0_1Dcon_eqZero_1I#_d  = {arg0_1Dcon_eqZero_1_d[32:1],
                                      (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0])};
  assign arg0_1Dcon_eqZero_1_r = (\arg0_1Dcon_eqZero_1I#_r  && (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0]));
  assign arg0_1Dcon_eqZero_2_r = (\arg0_1Dcon_eqZero_1I#_r  && (arg0_1Dcon_eqZero_2_d[0] && arg0_1Dcon_eqZero_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_1Dcon_eqZero_3,Int) (arg0_2Dcon_eqZero,Go) > [(arg0_1Dcon_eqZero_3I#,Go)] */
  assign \arg0_1Dcon_eqZero_3I#_d  = (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]);
  assign arg0_2Dcon_eqZero_r = (\arg0_1Dcon_eqZero_3I#_r  && (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]));
  assign arg0_1Dcon_eqZero_3_r = (\arg0_1Dcon_eqZero_3I#_r  && (arg0_1Dcon_eqZero_3_d[0] && arg0_2Dcon_eqZero_d[0]));
  
  /* fork (Ty Go) : (arg0_1Dcon_eqZero_3I#,Go) > [(arg0_1Dcon_eqZero_3I#_1,Go),
                                             (arg0_1Dcon_eqZero_3I#_2,Go),
                                             (arg0_1Dcon_eqZero_3I#_3,Go)] */
  logic [2:0] \arg0_1Dcon_eqZero_3I#_emitted ;
  logic [2:0] \arg0_1Dcon_eqZero_3I#_done ;
  assign \arg0_1Dcon_eqZero_3I#_1_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [0]));
  assign \arg0_1Dcon_eqZero_3I#_2_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [1]));
  assign \arg0_1Dcon_eqZero_3I#_3_d  = (\arg0_1Dcon_eqZero_3I#_d [0] && (! \arg0_1Dcon_eqZero_3I#_emitted [2]));
  assign \arg0_1Dcon_eqZero_3I#_done  = (\arg0_1Dcon_eqZero_3I#_emitted  | ({\arg0_1Dcon_eqZero_3I#_3_d [0],
                                                                             \arg0_1Dcon_eqZero_3I#_2_d [0],
                                                                             \arg0_1Dcon_eqZero_3I#_1_d [0]} & {\arg0_1Dcon_eqZero_3I#_3_r ,
                                                                                                                \arg0_1Dcon_eqZero_3I#_2_r ,
                                                                                                                \arg0_1Dcon_eqZero_3I#_1_r }));
  assign \arg0_1Dcon_eqZero_3I#_r  = (& \arg0_1Dcon_eqZero_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_emitted  <= 3'd0;
    else
      \arg0_1Dcon_eqZero_3I#_emitted  <= (\arg0_1Dcon_eqZero_3I#_r  ? 3'd0 :
                                          \arg0_1Dcon_eqZero_3I#_done );
  
  /* buf (Ty Go) : (arg0_1Dcon_eqZero_3I#_1,Go) > (arg0_1Dcon_eqZero_3I#_1_argbuf,Go) */
  Go_t \arg0_1Dcon_eqZero_3I#_1_bufchan_d ;
  logic \arg0_1Dcon_eqZero_3I#_1_bufchan_r ;
  assign \arg0_1Dcon_eqZero_3I#_1_r  = ((! \arg0_1Dcon_eqZero_3I#_1_bufchan_d [0]) || \arg0_1Dcon_eqZero_3I#_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_1_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_eqZero_3I#_1_r )
        \arg0_1Dcon_eqZero_3I#_1_bufchan_d  <= \arg0_1Dcon_eqZero_3I#_1_d ;
  Go_t \arg0_1Dcon_eqZero_3I#_1_bufchan_buf ;
  assign \arg0_1Dcon_eqZero_3I#_1_bufchan_r  = (! \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0]);
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_d  = (\arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0] ? \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  :
                                               \arg0_1Dcon_eqZero_3I#_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_eqZero_3I#_1_argbuf_r  && \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0]))
        \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_eqZero_3I#_1_argbuf_r ) && (! \arg0_1Dcon_eqZero_3I#_1_bufchan_buf [0])))
        \arg0_1Dcon_eqZero_3I#_1_bufchan_buf  <= \arg0_1Dcon_eqZero_3I#_1_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 0) : (arg0_1Dcon_eqZero_3I#_1_argbuf,Go) > (arg0_1Dcon_eqZero_3I#_1_argbuf_0,Int#) */
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_0_d  = {32'd0,
                                                 \arg0_1Dcon_eqZero_3I#_1_argbuf_d [0]};
  assign \arg0_1Dcon_eqZero_3I#_1_argbuf_r  = \arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ;
  
  /* op_eq (Ty Int#) : (arg0_1Dcon_eqZero_3I#_1_argbuf_0,Int#) (x1aph_destruct,Int#) > (lizzieLet1_1wild1X19_1_Eq,Bool) */
  assign lizzieLet1_1wild1X19_1_Eq_d = {(\arg0_1Dcon_eqZero_3I#_1_argbuf_0_d [32:1] == x1aph_destruct_d[32:1]),
                                        (\arg0_1Dcon_eqZero_3I#_1_argbuf_0_d [0] && x1aph_destruct_d[0])};
  assign {\arg0_1Dcon_eqZero_3I#_1_argbuf_0_r ,
          x1aph_destruct_r} = {2 {(lizzieLet1_1wild1X19_1_Eq_r && lizzieLet1_1wild1X19_1_Eq_d[0])}};
  
  /* buf (Ty Go) : (arg0_1Dcon_eqZero_3I#_2,Go) > (arg0_1Dcon_eqZero_3I#_2_argbuf,Go) */
  Go_t \arg0_1Dcon_eqZero_3I#_2_bufchan_d ;
  logic \arg0_1Dcon_eqZero_3I#_2_bufchan_r ;
  assign \arg0_1Dcon_eqZero_3I#_2_r  = ((! \arg0_1Dcon_eqZero_3I#_2_bufchan_d [0]) || \arg0_1Dcon_eqZero_3I#_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_2_bufchan_d  <= 1'd0;
    else
      if (\arg0_1Dcon_eqZero_3I#_2_r )
        \arg0_1Dcon_eqZero_3I#_2_bufchan_d  <= \arg0_1Dcon_eqZero_3I#_2_d ;
  Go_t \arg0_1Dcon_eqZero_3I#_2_bufchan_buf ;
  assign \arg0_1Dcon_eqZero_3I#_2_bufchan_r  = (! \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0]);
  assign \arg0_1Dcon_eqZero_3I#_2_argbuf_d  = (\arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0] ? \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  :
                                               \arg0_1Dcon_eqZero_3I#_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_1Dcon_eqZero_3I#_2_argbuf_r  && \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0]))
        \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= 1'd0;
      else if (((! \arg0_1Dcon_eqZero_3I#_2_argbuf_r ) && (! \arg0_1Dcon_eqZero_3I#_2_bufchan_buf [0])))
        \arg0_1Dcon_eqZero_3I#_2_bufchan_buf  <= \arg0_1Dcon_eqZero_3I#_2_bufchan_d ;
  
  /* dcon (Ty TupGo___Bool,
      Dcon TupGo___Bool) : [(arg0_1Dcon_eqZero_3I#_2_argbuf,Go),
                            (lizzieLet2_1_argbuf,Bool)] > (boolConvert_1TupGo___Bool_1,TupGo___Bool) */
  assign boolConvert_1TupGo___Bool_1_d = TupGo___Bool_dc((& {\arg0_1Dcon_eqZero_3I#_2_argbuf_d [0],
                                                             lizzieLet2_1_argbuf_d[0]}), \arg0_1Dcon_eqZero_3I#_2_argbuf_d , lizzieLet2_1_argbuf_d);
  assign {\arg0_1Dcon_eqZero_3I#_2_argbuf_r ,
          lizzieLet2_1_argbuf_r} = {2 {(boolConvert_1TupGo___Bool_1_r && boolConvert_1TupGo___Bool_1_d[0])}};
  
  /* mux (Ty Int,
     Ty MyBool) : (arg0_1Dcon_eqZero_4,Int) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[1:1],
                                                                             (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  assign arg0_1Dcon_eqZero_4_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r && (arg0_1Dcon_eqZero_4_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0]));
  
  /* demux (Ty MyDTInt_Bool,
       Ty Go) : (arg0_2,MyDTInt_Bool) (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8,Go) > [(arg0_2Dcon_eqZero,Go)] */
  assign arg0_2Dcon_eqZero_d = (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]);
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_r = (arg0_2Dcon_eqZero_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]));
  assign arg0_2_r = (arg0_2Dcon_eqZero_r && (arg0_2_d[0] && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Intgo_8_d[0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Int) : (arg0_2_1,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1,Int) > [(arg0_2_1Dcon_main1,Int)] */
  assign arg0_2_1Dcon_main1_d = {applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[32:1],
                                 (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0])};
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  assign arg0_2_1_r = (arg0_2_1Dcon_main1_r && (arg0_2_1_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intarg1_1_d[0]));
  
  /* fork (Ty Int) : (arg0_2_1Dcon_main1,Int) > [(arg0_2_1Dcon_main1_1,Int),
                                            (arg0_2_1Dcon_main1_2,Int),
                                            (arg0_2_1Dcon_main1_3,Int),
                                            (arg0_2_1Dcon_main1_4,Int)] */
  logic [3:0] arg0_2_1Dcon_main1_emitted;
  logic [3:0] arg0_2_1Dcon_main1_done;
  assign arg0_2_1Dcon_main1_1_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[0]))};
  assign arg0_2_1Dcon_main1_2_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[1]))};
  assign arg0_2_1Dcon_main1_3_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[2]))};
  assign arg0_2_1Dcon_main1_4_d = {arg0_2_1Dcon_main1_d[32:1],
                                   (arg0_2_1Dcon_main1_d[0] && (! arg0_2_1Dcon_main1_emitted[3]))};
  assign arg0_2_1Dcon_main1_done = (arg0_2_1Dcon_main1_emitted | ({arg0_2_1Dcon_main1_4_d[0],
                                                                   arg0_2_1Dcon_main1_3_d[0],
                                                                   arg0_2_1Dcon_main1_2_d[0],
                                                                   arg0_2_1Dcon_main1_1_d[0]} & {arg0_2_1Dcon_main1_4_r,
                                                                                                 arg0_2_1Dcon_main1_3_r,
                                                                                                 arg0_2_1Dcon_main1_2_r,
                                                                                                 arg0_2_1Dcon_main1_1_r}));
  assign arg0_2_1Dcon_main1_r = (& arg0_2_1Dcon_main1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) arg0_2_1Dcon_main1_emitted <= 4'd0;
    else
      arg0_2_1Dcon_main1_emitted <= (arg0_2_1Dcon_main1_r ? 4'd0 :
                                     arg0_2_1Dcon_main1_done);
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_2_1Dcon_main1_1I#,Int) > [(xap7_destruct,Int#)] */
  assign xap7_destruct_d = {\arg0_2_1Dcon_main1_1I#_d [32:1],
                            \arg0_2_1Dcon_main1_1I#_d [0]};
  assign \arg0_2_1Dcon_main1_1I#_r  = xap7_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_2_1Dcon_main1_2,Int) (arg0_2_1Dcon_main1_1,Int) > [(arg0_2_1Dcon_main1_1I#,Int)] */
  assign \arg0_2_1Dcon_main1_1I#_d  = {arg0_2_1Dcon_main1_1_d[32:1],
                                       (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0])};
  assign arg0_2_1Dcon_main1_1_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  assign arg0_2_1Dcon_main1_2_r = (\arg0_2_1Dcon_main1_1I#_r  && (arg0_2_1Dcon_main1_2_d[0] && arg0_2_1Dcon_main1_1_d[0]));
  
  /* demux (Ty Int,
       Ty Go) : (arg0_2_1Dcon_main1_3,Int) (arg0_2_2Dcon_main1,Go) > [(arg0_2_1Dcon_main1_3I#,Go)] */
  assign \arg0_2_1Dcon_main1_3I#_d  = (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]);
  assign arg0_2_2Dcon_main1_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  assign arg0_2_1Dcon_main1_3_r = (\arg0_2_1Dcon_main1_3I#_r  && (arg0_2_1Dcon_main1_3_d[0] && arg0_2_2Dcon_main1_d[0]));
  
  /* buf (Ty Go) : (arg0_2_1Dcon_main1_3I#,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) */
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  logic \arg0_2_1Dcon_main1_3I#_bufchan_r ;
  assign \arg0_2_1Dcon_main1_3I#_r  = ((! \arg0_2_1Dcon_main1_3I#_bufchan_d [0]) || \arg0_2_1Dcon_main1_3I#_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_d  <= 1'd0;
    else
      if (\arg0_2_1Dcon_main1_3I#_r )
        \arg0_2_1Dcon_main1_3I#_bufchan_d  <= \arg0_2_1Dcon_main1_3I#_d ;
  Go_t \arg0_2_1Dcon_main1_3I#_bufchan_buf ;
  assign \arg0_2_1Dcon_main1_3I#_bufchan_r  = (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]);
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_d  = (\arg0_2_1Dcon_main1_3I#_bufchan_buf [0] ? \arg0_2_1Dcon_main1_3I#_bufchan_buf  :
                                                \arg0_2_1Dcon_main1_3I#_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
    else
      if ((\arg0_2_1Dcon_main1_3I#_1_argbuf_r  && \arg0_2_1Dcon_main1_3I#_bufchan_buf [0]))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= 1'd0;
      else if (((! \arg0_2_1Dcon_main1_3I#_1_argbuf_r ) && (! \arg0_2_1Dcon_main1_3I#_bufchan_buf [0])))
        \arg0_2_1Dcon_main1_3I#_bufchan_buf  <= \arg0_2_1Dcon_main1_3I#_bufchan_d ;
  
  /* const (Ty Int#,
       Lit 2) : (arg0_2_1Dcon_main1_3I#_1_argbuf,Go) > (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) */
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d  = {32'd2,
                                                  \arg0_2_1Dcon_main1_3I#_1_argbuf_d [0]};
  assign \arg0_2_1Dcon_main1_3I#_1_argbuf_r  = \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r ;
  
  /* mux (Ty Int,
     Ty Int) : (arg0_2_1Dcon_main1_4,Int) [(es_0_1_1I#,Int)] > (es_0_1_1I#_mux,Int) */
  assign \es_0_1_1I#_mux_d  = {\es_0_1_1I#_d [32:1],
                               (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0])};
  assign \es_0_1_1I#_r  = (\es_0_1_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0]));
  assign arg0_2_1Dcon_main1_4_r = (\es_0_1_1I#_mux_r  && (arg0_2_1Dcon_main1_4_d[0] && \es_0_1_1I#_d [0]));
  
  /* demux (Ty MyDTInt_Int,
       Ty Go) : (arg0_2_2,MyDTInt_Int) (applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9,Go) > [(arg0_2_2Dcon_main1,Go)] */
  assign arg0_2_2Dcon_main1_d = (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]);
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]));
  assign arg0_2_2_r = (arg0_2_2Dcon_main1_r && (arg0_2_2_d[0] && applyfnInt_Int_5TupGo___MyDTInt_Int___Intgo_9_d[0]));
  
  /* mux (Ty MyDTInt_Int,
     Ty Int) : (arg0_2_3,MyDTInt_Int) [(es_0_1_1I#_mux,Int)] > (es_0_1_1I#_mux_mux,Int) */
  assign \es_0_1_1I#_mux_mux_d  = {\es_0_1_1I#_mux_d [32:1],
                                   (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0])};
  assign \es_0_1_1I#_mux_r  = (\es_0_1_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0]));
  assign arg0_2_3_r = (\es_0_1_1I#_mux_mux_r  && (arg0_2_3_d[0] && \es_0_1_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Bool,
     Ty MyBool) : (arg0_3,MyDTInt_Bool) [(lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[1:1],
                                                                                 (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0])};
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  assign arg0_3_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_mux_r && (arg0_3_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_1,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2,Int) > [(arg0_4_1Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_4_1Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[32:1],
                                              (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_r = (\arg0_4_1Dcon_$fNumInt_$ctimes_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  assign arg0_4_1_r = (\arg0_4_1Dcon_$fNumInt_$ctimes_r  && (arg0_4_1_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg1_2_d[0]));
  
  /* demux (Ty MyDTInt_Int_Int,
       Ty Int) : (arg0_4_2,MyDTInt_Int_Int) (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2,Int) > [(arg0_4_2Dcon_$fNumInt_$c*,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_d  = {applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[32:1],
                                              (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0])};
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  assign arg0_4_2_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_r  && (arg0_4_2_d[0] && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Intarg2_d[0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_1,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_2,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_3,Int),
                                                   (arg0_4_2Dcon_$fNumInt_$c*_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_done ;
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_2_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_4_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_d [32:1],
                                                (\arg0_4_2Dcon_$fNumInt_$ctimes_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_done  = (\arg0_4_2Dcon_$fNumInt_$ctimes_emitted  | ({\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0],
                                                                                             \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$ctimes_4_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_3_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_2_r ,
                                                                                                                                        \arg0_4_2Dcon_$fNumInt_$ctimes_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_r  = (& \arg0_4_2Dcon_$fNumInt_$ctimes_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$ctimes_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$ctimes_emitted  <= (\arg0_4_2Dcon_$fNumInt_$ctimes_r  ? 4'd0 :
                                                  \arg0_4_2Dcon_$fNumInt_$ctimes_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c*_1I#,Int) > [(xa1m0_destruct,Int#)] */
  assign xa1m0_destruct_d = {\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  = xa1m0_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_2,Int) (arg0_4_2Dcon_$fNumInt_$c*_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_1_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_1_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_2_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3,Int) (arg0_4_1Dcon_$fNumInt_$c*,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d  = {\arg0_4_1Dcon_$fNumInt_$ctimes_d [32:1],
                                                  (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0])};
  assign \arg0_4_1Dcon_$fNumInt_$ctimes_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3_d [0] && \arg0_4_1Dcon_$fNumInt_$ctimes_d [0]));
  
  /* fork (Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_1,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_2,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_3,Int),
                                                       (arg0_4_2Dcon_$fNumInt_$c*_3I#_4,Int)] */
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted ;
  logic [3:0] \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done ;
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [0]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [1]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [2]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [32:1],
                                                    (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_d [0] && (! \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted [3]))};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  | ({\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0],
                                                                                                     \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]} & {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r ,
                                                                                                                                                    \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r }));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  = (& \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= 4'd0;
    else
      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_emitted  <= (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_r  ? 4'd0 :
                                                      \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_done );
  
  /* destruct (Ty Int,
          Dcon I#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_1I#,Int) > [(ya1m1_destruct,Int#)] */
  assign ya1m1_destruct_d = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [32:1],
                             \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d [0]};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  = ya1m1_destruct_r;
  
  /* demux (Ty Int,
       Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_2,Int) (arg0_4_2Dcon_$fNumInt_$c*_3I#_1,Int) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_1I#,Int)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_d  = {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [32:1],
                                                      (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0])};
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_2_d [0] && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_1_d [0]));
  
  /* demux (Ty Int,
       Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_3,Int) (xa1m0_destruct,Int#) > [(arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#,Int#)] */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d  = {xa1m0_destruct_d[32:1],
                                                      (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0])};
  assign xa1m0_destruct_r = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_r  = (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3_d [0] && xa1m0_destruct_d[0]));
  
  /* op_mul (Ty Int#) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#,Int#) (ya1m1_destruct,Int#) > (arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#) */
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d  = {(\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [32:1] * ya1m1_destruct_d[32:1]),
                                                                     (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_d [0] && ya1m1_destruct_d[0])};
  assign {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_r ,
          ya1m1_destruct_r} = {2 {(\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r  && \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(arg0_4_2Dcon_$fNumInt_$c*_3I#_3I#_1ya1m1_1_Mul32,Int#)] > (es_0_2_1I#,Int) */
  assign \es_0_2_1I#_d  = \I#_dc ((& {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d [0]}), \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_d );
  assign {\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_3I#_1ya1m1_1_Mul32_r } = {1 {(\es_0_2_1I#_r  && \es_0_2_1I#_d [0])}};
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_3I#_4,Int) [(es_0_2_1I#,Int)] > (es_0_2_1I#_mux,Int) */
  assign \es_0_2_1I#_mux_d  = {\es_0_2_1I#_d [32:1],
                               (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_2_1I#_d [0])};
  assign \es_0_2_1I#_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_r  = (\es_0_2_1I#_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_3I#_4_d [0] && \es_0_2_1I#_d [0]));
  
  /* mux (Ty Int,
     Ty Int) : (arg0_4_2Dcon_$fNumInt_$c*_4,Int) [(es_0_2_1I#_mux,Int)] > (es_0_2_1I#_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_d  = {\es_0_2_1I#_mux_d [32:1],
                                   (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_2_1I#_mux_d [0])};
  assign \es_0_2_1I#_mux_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_2_1I#_mux_d [0]));
  assign \arg0_4_2Dcon_$fNumInt_$ctimes_4_r  = (\es_0_2_1I#_mux_mux_r  && (\arg0_4_2Dcon_$fNumInt_$ctimes_4_d [0] && \es_0_2_1I#_mux_d [0]));
  
  /* mux (Ty MyDTInt_Int_Int,
     Ty Int) : (arg0_4_3,MyDTInt_Int_Int) [(es_0_2_1I#_mux_mux,Int)] > (es_0_2_1I#_mux_mux_mux,Int) */
  assign \es_0_2_1I#_mux_mux_mux_d  = {\es_0_2_1I#_mux_mux_d [32:1],
                                       (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0])};
  assign \es_0_2_1I#_mux_mux_r  = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  assign arg0_4_3_r = (\es_0_2_1I#_mux_mux_mux_r  && (arg0_4_3_d[0] && \es_0_2_1I#_mux_mux_d [0]));
  
  /* destruct (Ty TupGo___Bool,
          Dcon TupGo___Bool) : (boolConvert_1TupGo___Bool_1,TupGo___Bool) > [(boolConvert_1TupGo___Boolgo_1,Go),
                                                                             (boolConvert_1TupGo___Boolbool,Bool)] */
  logic [1:0] boolConvert_1TupGo___Bool_1_emitted;
  logic [1:0] boolConvert_1TupGo___Bool_1_done;
  assign boolConvert_1TupGo___Boolgo_1_d = (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[0]));
  assign boolConvert_1TupGo___Boolbool_d = {boolConvert_1TupGo___Bool_1_d[1:1],
                                            (boolConvert_1TupGo___Bool_1_d[0] && (! boolConvert_1TupGo___Bool_1_emitted[1]))};
  assign boolConvert_1TupGo___Bool_1_done = (boolConvert_1TupGo___Bool_1_emitted | ({boolConvert_1TupGo___Boolbool_d[0],
                                                                                     boolConvert_1TupGo___Boolgo_1_d[0]} & {boolConvert_1TupGo___Boolbool_r,
                                                                                                                            boolConvert_1TupGo___Boolgo_1_r}));
  assign boolConvert_1TupGo___Bool_1_r = (& boolConvert_1TupGo___Bool_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Bool_1_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Bool_1_emitted <= (boolConvert_1TupGo___Bool_1_r ? 2'd0 :
                                              boolConvert_1TupGo___Bool_1_done);
  
  /* fork (Ty Bool) : (boolConvert_1TupGo___Boolbool,Bool) > [(bool_1,Bool),
                                                         (bool_2,Bool)] */
  logic [1:0] boolConvert_1TupGo___Boolbool_emitted;
  logic [1:0] boolConvert_1TupGo___Boolbool_done;
  assign bool_1_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[0]))};
  assign bool_2_d = {boolConvert_1TupGo___Boolbool_d[1:1],
                     (boolConvert_1TupGo___Boolbool_d[0] && (! boolConvert_1TupGo___Boolbool_emitted[1]))};
  assign boolConvert_1TupGo___Boolbool_done = (boolConvert_1TupGo___Boolbool_emitted | ({bool_2_d[0],
                                                                                         bool_1_d[0]} & {bool_2_r,
                                                                                                         bool_1_r}));
  assign boolConvert_1TupGo___Boolbool_r = (& boolConvert_1TupGo___Boolbool_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1TupGo___Boolbool_emitted <= 2'd0;
    else
      boolConvert_1TupGo___Boolbool_emitted <= (boolConvert_1TupGo___Boolbool_r ? 2'd0 :
                                                boolConvert_1TupGo___Boolbool_done);
  
  /* fork (Ty MyBool) : (boolConvert_1_resbuf,MyBool) > [(lizzieLet3_1,MyBool),
                                                    (lizzieLet3_2,MyBool)] */
  logic [1:0] boolConvert_1_resbuf_emitted;
  logic [1:0] boolConvert_1_resbuf_done;
  assign lizzieLet3_1_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[0]))};
  assign lizzieLet3_2_d = {boolConvert_1_resbuf_d[1:1],
                           (boolConvert_1_resbuf_d[0] && (! boolConvert_1_resbuf_emitted[1]))};
  assign boolConvert_1_resbuf_done = (boolConvert_1_resbuf_emitted | ({lizzieLet3_2_d[0],
                                                                       lizzieLet3_1_d[0]} & {lizzieLet3_2_r,
                                                                                             lizzieLet3_1_r}));
  assign boolConvert_1_resbuf_r = (& boolConvert_1_resbuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) boolConvert_1_resbuf_emitted <= 2'd0;
    else
      boolConvert_1_resbuf_emitted <= (boolConvert_1_resbuf_r ? 2'd0 :
                                       boolConvert_1_resbuf_done);
  
  /* demux (Ty Bool,
       Ty Go) : (bool_1,Bool) (boolConvert_1TupGo___Boolgo_1,Go) > [(bool_1False,Go),
                                                                    (bool_1True,Go)] */
  logic [1:0] boolConvert_1TupGo___Boolgo_1_onehotd;
  always_comb
    if ((bool_1_d[0] && boolConvert_1TupGo___Boolgo_1_d[0]))
      unique case (bool_1_d[1:1])
        1'd0: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd1;
        1'd1: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd2;
        default: boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
      endcase
    else boolConvert_1TupGo___Boolgo_1_onehotd = 2'd0;
  assign bool_1False_d = boolConvert_1TupGo___Boolgo_1_onehotd[0];
  assign bool_1True_d = boolConvert_1TupGo___Boolgo_1_onehotd[1];
  assign boolConvert_1TupGo___Boolgo_1_r = (| (boolConvert_1TupGo___Boolgo_1_onehotd & {bool_1True_r,
                                                                                        bool_1False_r}));
  assign bool_1_r = boolConvert_1TupGo___Boolgo_1_r;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(bool_1False,Go)] > (bool_1False_1MyFalse,MyBool) */
  assign bool_1False_1MyFalse_d = MyFalse_dc((& {bool_1False_d[0]}), bool_1False_d);
  assign {bool_1False_r} = {1 {(bool_1False_1MyFalse_r && bool_1False_1MyFalse_d[0])}};
  
  /* buf (Ty MyBool) : (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) > (boolConvert_1_resbuf,MyBool) */
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  logic bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_r = ((! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d[0]) || bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= {1'd0,
                                                               1'd0};
    else
      if (bool_1False_1MyFalsebool_1True_1MyTrue_mux_r)
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_d;
  MyBool_t bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf;
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_r = (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]);
  assign boolConvert_1_resbuf_d = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0] ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf :
                                   bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                 1'd0};
    else
      if ((boolConvert_1_resbuf_r && bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0]))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= {1'd0,
                                                                   1'd0};
      else if (((! boolConvert_1_resbuf_r) && (! bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf[0])))
        bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_buf <= bool_1False_1MyFalsebool_1True_1MyTrue_mux_bufchan_d;
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(bool_1True,Go)] > (bool_1True_1MyTrue,MyBool) */
  assign bool_1True_1MyTrue_d = MyTrue_dc((& {bool_1True_d[0]}), bool_1True_d);
  assign {bool_1True_r} = {1 {(bool_1True_1MyTrue_r && bool_1True_1MyTrue_d[0])}};
  
  /* mux (Ty Bool,
     Ty MyBool) : (bool_2,Bool) [(bool_1False_1MyFalse,MyBool),
                                 (bool_1True_1MyTrue,MyBool)] > (bool_1False_1MyFalsebool_1True_1MyTrue_mux,MyBool) */
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux;
  logic [1:0] bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot;
  always_comb
    unique case (bool_2_d[1:1])
      1'd0:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd1,
                                                            bool_1False_1MyFalse_d};
      1'd1:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd2,
                                                            bool_1True_1MyTrue_d};
      default:
        {bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot,
         bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux} = {2'd0,
                                                            {1'd0, 1'd0}};
    endcase
  assign bool_1False_1MyFalsebool_1True_1MyTrue_mux_d = {bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[1:1],
                                                         (bool_1False_1MyFalsebool_1True_1MyTrue_mux_mux[0] && bool_2_d[0])};
  assign bool_2_r = (bool_1False_1MyFalsebool_1True_1MyTrue_mux_d[0] && bool_1False_1MyFalsebool_1True_1MyTrue_mux_r);
  assign {bool_1True_1MyTrue_r,
          bool_1False_1MyFalse_r} = (bool_2_r ? bool_1False_1MyFalsebool_1True_1MyTrue_mux_onehot :
                                     2'd0);
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) > [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10,Go),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1,Pointer_QTree_Int),
                                                                                                                                                                                       (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] */
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted;
  logic [2:0] call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done;
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[0]));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[16:1],
                                                                                  (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[1]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[32:17],
                                                                                (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0] && (! call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted[2]))};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done = (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted | ({call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d[0],
                                                                                                                                                             call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d[0]} & {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r,
                                                                                                                                                                                                                                         call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_r,
                                                                                                                                                                                                                                         call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_r}));
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r = (& call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= 3'd0;
    else
      call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_emitted <= (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r ? 3'd0 :
                                                                                  call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_done);
  
  /* rbuf (Ty Go) : (call_$wnnz_Int_goConst,Go) > (call_$wnnz_Int_initBufi,Go) */
  Go_t call_$wnnz_Int_goConst_buf;
  assign call_$wnnz_Int_goConst_r = (! call_$wnnz_Int_goConst_buf[0]);
  assign call_$wnnz_Int_initBufi_d = (call_$wnnz_Int_goConst_buf[0] ? call_$wnnz_Int_goConst_buf :
                                      call_$wnnz_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goConst_buf <= 1'd0;
    else
      if ((call_$wnnz_Int_initBufi_r && call_$wnnz_Int_goConst_buf[0]))
        call_$wnnz_Int_goConst_buf <= 1'd0;
      else if (((! call_$wnnz_Int_initBufi_r) && (! call_$wnnz_Int_goConst_buf[0])))
        call_$wnnz_Int_goConst_buf <= call_$wnnz_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_$wnnz_Int_goMux1,Go),
                           (lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf,Go),
                           (lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf,Go),
                           (lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf,Go),
                           (lizzieLet4_3QNode_Int_1_argbuf,Go)] > (go_10_goMux_choice,C5) (go_10_goMux_data,Go) */
  logic [4:0] call_$wnnz_Int_goMux1_select_d;
  assign call_$wnnz_Int_goMux1_select_d = ((| call_$wnnz_Int_goMux1_select_q) ? call_$wnnz_Int_goMux1_select_q :
                                           (call_$wnnz_Int_goMux1_d[0] ? 5'd1 :
                                            (lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_d[0] ? 5'd2 :
                                             (lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_d[0] ? 5'd4 :
                                              (lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_d[0] ? 5'd8 :
                                               (lizzieLet4_3QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                5'd0))))));
  logic [4:0] call_$wnnz_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_select_q <= 5'd0;
    else
      call_$wnnz_Int_goMux1_select_q <= (call_$wnnz_Int_goMux1_done ? 5'd0 :
                                         call_$wnnz_Int_goMux1_select_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_goMux1_emit_q <= 2'd0;
    else
      call_$wnnz_Int_goMux1_emit_q <= (call_$wnnz_Int_goMux1_done ? 2'd0 :
                                       call_$wnnz_Int_goMux1_emit_d);
  logic [1:0] call_$wnnz_Int_goMux1_emit_d;
  assign call_$wnnz_Int_goMux1_emit_d = (call_$wnnz_Int_goMux1_emit_q | ({go_10_goMux_choice_d[0],
                                                                          go_10_goMux_data_d[0]} & {go_10_goMux_choice_r,
                                                                                                    go_10_goMux_data_r}));
  logic call_$wnnz_Int_goMux1_done;
  assign call_$wnnz_Int_goMux1_done = (& call_$wnnz_Int_goMux1_emit_d);
  assign {lizzieLet4_3QNode_Int_1_argbuf_r,
          lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_r,
          lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_r,
          lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_r,
          call_$wnnz_Int_goMux1_r} = (call_$wnnz_Int_goMux1_done ? call_$wnnz_Int_goMux1_select_d :
                                      5'd0);
  assign go_10_goMux_data_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? call_$wnnz_Int_goMux1_d :
                               ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_d :
                                ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_d :
                                 ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_d :
                                  ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[0])) ? lizzieLet4_3QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_10_goMux_choice_d = ((call_$wnnz_Int_goMux1_select_d[0] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_$wnnz_Int_goMux1_select_d[1] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_$wnnz_Int_goMux1_select_d[2] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_$wnnz_Int_goMux1_select_d[3] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_$wnnz_Int_goMux1_select_d[4] && (! call_$wnnz_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_$wnnz_Int_initBuf,Go) > [(call_$wnnz_Int_unlockFork1,Go),
                                              (call_$wnnz_Int_unlockFork2,Go),
                                              (call_$wnnz_Int_unlockFork3,Go)] */
  logic [2:0] call_$wnnz_Int_initBuf_emitted;
  logic [2:0] call_$wnnz_Int_initBuf_done;
  assign call_$wnnz_Int_unlockFork1_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[0]));
  assign call_$wnnz_Int_unlockFork2_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[1]));
  assign call_$wnnz_Int_unlockFork3_d = (call_$wnnz_Int_initBuf_d[0] && (! call_$wnnz_Int_initBuf_emitted[2]));
  assign call_$wnnz_Int_initBuf_done = (call_$wnnz_Int_initBuf_emitted | ({call_$wnnz_Int_unlockFork3_d[0],
                                                                           call_$wnnz_Int_unlockFork2_d[0],
                                                                           call_$wnnz_Int_unlockFork1_d[0]} & {call_$wnnz_Int_unlockFork3_r,
                                                                                                               call_$wnnz_Int_unlockFork2_r,
                                                                                                               call_$wnnz_Int_unlockFork1_r}));
  assign call_$wnnz_Int_initBuf_r = (& call_$wnnz_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_emitted <= 3'd0;
    else
      call_$wnnz_Int_initBuf_emitted <= (call_$wnnz_Int_initBuf_r ? 3'd0 :
                                         call_$wnnz_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_$wnnz_Int_initBufi,Go) > (call_$wnnz_Int_initBuf,Go) */
  assign call_$wnnz_Int_initBufi_r = ((! call_$wnnz_Int_initBuf_d[0]) || call_$wnnz_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_$wnnz_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_$wnnz_Int_initBufi_r)
        call_$wnnz_Int_initBuf_d <= call_$wnnz_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_$wnnz_Int_unlockFork1,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10,Go)] > (call_$wnnz_Int_goMux1,Go) */
  assign call_$wnnz_Int_goMux1_d = (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d[0]);
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d[0]));
  assign call_$wnnz_Int_unlockFork1_r = (call_$wnnz_Int_goMux1_r && (call_$wnnz_Int_unlockFork1_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intgo_10_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_$wnnz_Int_unlockFork2,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1,Pointer_QTree_Int)] > (call_$wnnz_Int_goMux2,Pointer_QTree_Int) */
  assign call_$wnnz_Int_goMux2_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d[16:1],
                                    (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d[0]));
  assign call_$wnnz_Int_unlockFork2_r = (call_$wnnz_Int_goMux2_r && (call_$wnnz_Int_unlockFork2_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_IntwstH_1_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CT$wnnz_Int) : (call_$wnnz_Int_unlockFork3,Go) [(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0,Pointer_CT$wnnz_Int)] > (call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int) */
  assign call_$wnnz_Int_goMux3_d = {call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[16:1],
                                    (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0])};
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  assign call_$wnnz_Int_unlockFork3_r = (call_$wnnz_Int_goMux3_r && (call_$wnnz_Int_unlockFork3_d[0] && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Intsc_0_d[0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int) : (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int) > [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8,Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                   (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [7:0] \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted ;
  logic [7:0] \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_done ;
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [0]));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [16:1],
                                                                                                                                                                               (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [1]))};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [2]));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [3]));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [48:17],
                                                                                                                                                                              (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [4]))};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [5]));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [6]));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [64:49],
                                                                                                                                                                                (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0] && (! \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted [7]))};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_done  = (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted  | ({\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d [0],
                                                                                                                                                                                                                                                                                                                                                         \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d [0]} & {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_r ,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_r }));
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_r  = (& \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted  <= 8'd0;
    else
      \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_emitted  <= (\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_r  ? 8'd0 :
                                                                                                                                                                                \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_done );
  
  /* rbuf (Ty Go) : (call_f'_f'_Int_Int_Int_Int_goConst,Go) > (call_f'_f'_Int_Int_Int_Int_initBufi,Go) */
  Go_t \call_f'_f'_Int_Int_Int_Int_goConst_buf ;
  assign \call_f'_f'_Int_Int_Int_Int_goConst_r  = (! \call_f'_f'_Int_Int_Int_Int_goConst_buf [0]);
  assign \call_f'_f'_Int_Int_Int_Int_initBufi_d  = (\call_f'_f'_Int_Int_Int_Int_goConst_buf [0] ? \call_f'_f'_Int_Int_Int_Int_goConst_buf  :
                                                    \call_f'_f'_Int_Int_Int_Int_goConst_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_Int_goConst_buf  <= 1'd0;
    else
      if ((\call_f'_f'_Int_Int_Int_Int_initBufi_r  && \call_f'_f'_Int_Int_Int_Int_goConst_buf [0]))
        \call_f'_f'_Int_Int_Int_Int_goConst_buf  <= 1'd0;
      else if (((! \call_f'_f'_Int_Int_Int_Int_initBufi_r ) && (! \call_f'_f'_Int_Int_Int_Int_goConst_buf [0])))
        \call_f'_f'_Int_Int_Int_Int_goConst_buf  <= \call_f'_f'_Int_Int_Int_Int_goConst_d ;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f'_f'_Int_Int_Int_Int_goMux1,Go),
                           (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf,Go),
                           (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf,Go),
                           (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf,Go),
                           (lizzieLet6_4QNode_Int_1_argbuf,Go)] > (go_11_goMux_choice,C5) (go_11_goMux_data,Go) */
  logic [4:0] \call_f'_f'_Int_Int_Int_Int_goMux1_select_d ;
  assign \call_f'_f'_Int_Int_Int_Int_goMux1_select_d  = ((| \call_f'_f'_Int_Int_Int_Int_goMux1_select_q ) ? \call_f'_f'_Int_Int_Int_Int_goMux1_select_q  :
                                                         (\call_f'_f'_Int_Int_Int_Int_goMux1_d [0] ? 5'd1 :
                                                          (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_d [0] ? 5'd2 :
                                                           (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_d [0] ? 5'd4 :
                                                            (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_d [0] ? 5'd8 :
                                                             (lizzieLet6_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                              5'd0))))));
  logic [4:0] \call_f'_f'_Int_Int_Int_Int_goMux1_select_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_Int_goMux1_select_q  <= 5'd0;
    else
      \call_f'_f'_Int_Int_Int_Int_goMux1_select_q  <= (\call_f'_f'_Int_Int_Int_Int_goMux1_done  ? 5'd0 :
                                                       \call_f'_f'_Int_Int_Int_Int_goMux1_select_d );
  logic [1:0] \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q ;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q  <= 2'd0;
    else
      \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q  <= (\call_f'_f'_Int_Int_Int_Int_goMux1_done  ? 2'd0 :
                                                     \call_f'_f'_Int_Int_Int_Int_goMux1_emit_d );
  logic [1:0] \call_f'_f'_Int_Int_Int_Int_goMux1_emit_d ;
  assign \call_f'_f'_Int_Int_Int_Int_goMux1_emit_d  = (\call_f'_f'_Int_Int_Int_Int_goMux1_emit_q  | ({go_11_goMux_choice_d[0],
                                                                                                      go_11_goMux_data_d[0]} & {go_11_goMux_choice_r,
                                                                                                                                go_11_goMux_data_r}));
  logic \call_f'_f'_Int_Int_Int_Int_goMux1_done ;
  assign \call_f'_f'_Int_Int_Int_Int_goMux1_done  = (& \call_f'_f'_Int_Int_Int_Int_goMux1_emit_d );
  assign {lizzieLet6_4QNode_Int_1_argbuf_r,
          \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_r ,
          \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_r ,
          \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_r ,
          \call_f'_f'_Int_Int_Int_Int_goMux1_r } = (\call_f'_f'_Int_Int_Int_Int_goMux1_done  ? \call_f'_f'_Int_Int_Int_Int_goMux1_select_d  :
                                                    5'd0);
  assign go_11_goMux_data_d = ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [0] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [0])) ? \call_f'_f'_Int_Int_Int_Int_goMux1_d  :
                               ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [1] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_d  :
                                ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [2] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_d  :
                                 ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [3] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [0])) ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_d  :
                                  ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [4] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [0])) ? lizzieLet6_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_11_goMux_choice_d = ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [0] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [1])) ? C1_5_dc(1'd1) :
                                 ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [1] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [1])) ? C2_5_dc(1'd1) :
                                  ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [2] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [1])) ? C3_5_dc(1'd1) :
                                   ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [3] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [1])) ? C4_5_dc(1'd1) :
                                    ((\call_f'_f'_Int_Int_Int_Int_goMux1_select_d [4] && (! \call_f'_f'_Int_Int_Int_Int_goMux1_emit_q [1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f'_f'_Int_Int_Int_Int_initBuf,Go) > [(call_f'_f'_Int_Int_Int_Int_unlockFork1,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork2,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork3,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork4,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork5,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork6,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork7,Go),
                                                          (call_f'_f'_Int_Int_Int_Int_unlockFork8,Go)] */
  logic [7:0] \call_f'_f'_Int_Int_Int_Int_initBuf_emitted ;
  logic [7:0] \call_f'_f'_Int_Int_Int_Int_initBuf_done ;
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork1_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork2_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [1]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork3_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [2]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork4_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [3]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork5_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [4]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork6_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [5]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork7_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [6]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork8_d  = (\call_f'_f'_Int_Int_Int_Int_initBuf_d [0] && (! \call_f'_f'_Int_Int_Int_Int_initBuf_emitted [7]));
  assign \call_f'_f'_Int_Int_Int_Int_initBuf_done  = (\call_f'_f'_Int_Int_Int_Int_initBuf_emitted  | ({\call_f'_f'_Int_Int_Int_Int_unlockFork8_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork7_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork6_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork5_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork4_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork3_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork2_d [0],
                                                                                                       \call_f'_f'_Int_Int_Int_Int_unlockFork1_d [0]} & {\call_f'_f'_Int_Int_Int_Int_unlockFork8_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork7_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork6_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork5_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork4_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork3_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork2_r ,
                                                                                                                                                         \call_f'_f'_Int_Int_Int_Int_unlockFork1_r }));
  assign \call_f'_f'_Int_Int_Int_Int_initBuf_r  = (& \call_f'_f'_Int_Int_Int_Int_initBuf_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_Int_initBuf_emitted  <= 8'd0;
    else
      \call_f'_f'_Int_Int_Int_Int_initBuf_emitted  <= (\call_f'_f'_Int_Int_Int_Int_initBuf_r  ? 8'd0 :
                                                       \call_f'_f'_Int_Int_Int_Int_initBuf_done );
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f'_f'_Int_Int_Int_Int_initBufi,Go) > (call_f'_f'_Int_Int_Int_Int_initBuf,Go) */
  assign \call_f'_f'_Int_Int_Int_Int_initBufi_r  = ((! \call_f'_f'_Int_Int_Int_Int_initBuf_d [0]) || \call_f'_f'_Int_Int_Int_Int_initBuf_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \call_f'_f'_Int_Int_Int_Int_initBuf_d  <= Go_dc(1'd1);
    else
      if (\call_f'_f'_Int_Int_Int_Int_initBufi_r )
        \call_f'_f'_Int_Int_Int_Int_initBuf_d  <= \call_f'_f'_Int_Int_Int_Int_initBufi_d ;
  
  /* mux (Ty Go,
     Ty Go) : (call_f'_f'_Int_Int_Int_Int_unlockFork1,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11,Go)] > (call_f'_f'_Int_Int_Int_Int_goMux1,Go) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux1_d  = (\call_f'_f'_Int_Int_Int_Int_unlockFork1_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d [0]);
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_r  = (\call_f'_f'_Int_Int_Int_Int_goMux1_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork1_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork1_r  = (\call_f'_f'_Int_Int_Int_Int_goMux1_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork1_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intgo_11_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f'_f'_Int_Int_Int_Int_unlockFork2,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5,Pointer_QTree_Int)] > (call_f'_f'_Int_Int_Int_Int_goMux2,Pointer_QTree_Int) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux2_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d [16:1],
                                                  (\call_f'_f'_Int_Int_Int_Int_unlockFork2_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d [0])};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_r  = (\call_f'_f'_Int_Int_Int_Int_goMux2_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork2_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork2_r  = (\call_f'_f'_Int_Int_Int_Int_goMux2_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork2_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intm2ai5_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f'_f'_Int_Int_Int_Int_unlockFork3,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6,MyDTInt_Bool)] > (call_f'_f'_Int_Int_Int_Int_goMux3,MyDTInt_Bool) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux3_d  = (\call_f'_f'_Int_Int_Int_Int_unlockFork3_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d [0]);
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_r  = (\call_f'_f'_Int_Int_Int_Int_goMux3_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork3_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork3_r  = (\call_f'_f'_Int_Int_Int_Int_goMux3_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork3_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_kronai6_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f'_f'_Int_Int_Int_Int_unlockFork4,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7,MyDTInt_Int_Int)] > (call_f'_f'_Int_Int_Int_Int_goMux4,MyDTInt_Int_Int) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux4_d  = (\call_f'_f'_Int_Int_Int_Int_unlockFork4_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d [0]);
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_r  = (\call_f'_f'_Int_Int_Int_Int_goMux4_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork4_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork4_r  = (\call_f'_f'_Int_Int_Int_Int_goMux4_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork4_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intop_kronai7_d [0]));
  
  /* mux (Ty Go,
     Ty Int) : (call_f'_f'_Int_Int_Int_Int_unlockFork5,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8,Int)] > (call_f'_f'_Int_Int_Int_Int_goMux5,Int) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux5_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d [32:1],
                                                  (\call_f'_f'_Int_Int_Int_Int_unlockFork5_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d [0])};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_r  = (\call_f'_f'_Int_Int_Int_Int_goMux5_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork5_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork5_r  = (\call_f'_f'_Int_Int_Int_Int_goMux5_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork5_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intvai8_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f'_f'_Int_Int_Int_Int_unlockFork6,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9,MyDTInt_Bool)] > (call_f'_f'_Int_Int_Int_Int_goMux6,MyDTInt_Bool) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux6_d  = (\call_f'_f'_Int_Int_Int_Int_unlockFork6_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d [0]);
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_r  = (\call_f'_f'_Int_Int_Int_Int_goMux6_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork6_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork6_r  = (\call_f'_f'_Int_Int_Int_Int_goMux6_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork6_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intis_z_mapai9_d [0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int) : (call_f'_f'_Int_Int_Int_Int_unlockFork7,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia,MyDTInt_Int)] > (call_f'_f'_Int_Int_Int_Int_goMux7,MyDTInt_Int) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux7_d  = (\call_f'_f'_Int_Int_Int_Int_unlockFork7_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d [0]);
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_r  = (\call_f'_f'_Int_Int_Int_Int_goMux7_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork7_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork7_r  = (\call_f'_f'_Int_Int_Int_Int_goMux7_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork7_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intf_mapaia_d [0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (call_f'_f'_Int_Int_Int_Int_unlockFork8,Go) [(call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1,Pointer_CTf'_f'_Int_Int_Int_Int)] > (call_f'_f'_Int_Int_Int_Int_goMux8,Pointer_CTf'_f'_Int_Int_Int_Int) */
  assign \call_f'_f'_Int_Int_Int_Int_goMux8_d  = {\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d [16:1],
                                                  (\call_f'_f'_Int_Int_Int_Int_unlockFork8_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d [0])};
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_r  = (\call_f'_f'_Int_Int_Int_Int_goMux8_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork8_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d [0]));
  assign \call_f'_f'_Int_Int_Int_Int_unlockFork8_r  = (\call_f'_f'_Int_Int_Int_Int_goMux8_r  && (\call_f'_f'_Int_Int_Int_Int_unlockFork8_d [0] && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Intsc_0_1_d [0]));
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int) : (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int) > [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12,Go),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ,MyDTInt_Int),
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2,Pointer_CTf_f_Int_Int_Int_Int)] */
  logic [7:0] call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted;
  logic [7:0] call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_done;
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[0]));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[16:1],
                                                                                                                                                                                       (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[1]))};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[32:17],
                                                                                                                                                                                       (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[2]))};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[3]));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[4]));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[5]));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[6]));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[48:33],
                                                                                                                                                                                        (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0] && (! call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted[7]))};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_done = (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted | ({call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d[0],
                                                                                                                                                                                                                                                                                                                                                                         call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d[0]} & {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_r}));
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_r = (& call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted <= 8'd0;
    else
      call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_emitted <= (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_r ? 8'd0 :
                                                                                                                                                                                        call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_done);
  
  /* rbuf (Ty Go) : (call_f_f_Int_Int_Int_Int_goConst,Go) > (call_f_f_Int_Int_Int_Int_initBufi,Go) */
  Go_t call_f_f_Int_Int_Int_Int_goConst_buf;
  assign call_f_f_Int_Int_Int_Int_goConst_r = (! call_f_f_Int_Int_Int_Int_goConst_buf[0]);
  assign call_f_f_Int_Int_Int_Int_initBufi_d = (call_f_f_Int_Int_Int_Int_goConst_buf[0] ? call_f_f_Int_Int_Int_Int_goConst_buf :
                                                call_f_f_Int_Int_Int_Int_goConst_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) call_f_f_Int_Int_Int_Int_goConst_buf <= 1'd0;
    else
      if ((call_f_f_Int_Int_Int_Int_initBufi_r && call_f_f_Int_Int_Int_Int_goConst_buf[0]))
        call_f_f_Int_Int_Int_Int_goConst_buf <= 1'd0;
      else if (((! call_f_f_Int_Int_Int_Int_initBufi_r) && (! call_f_f_Int_Int_Int_Int_goConst_buf[0])))
        call_f_f_Int_Int_Int_Int_goConst_buf <= call_f_f_Int_Int_Int_Int_goConst_d;
  
  /* mergectrl (Ty C5,Ty Go) : [(call_f_f_Int_Int_Int_Int_goMux1,Go),
                           (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf,Go),
                           (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf,Go),
                           (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf,Go),
                           (lizzieLet13_1_4QNode_Int_1_argbuf,Go)] > (go_12_goMux_choice,C5) (go_12_goMux_data,Go) */
  logic [4:0] call_f_f_Int_Int_Int_Int_goMux1_select_d;
  assign call_f_f_Int_Int_Int_Int_goMux1_select_d = ((| call_f_f_Int_Int_Int_Int_goMux1_select_q) ? call_f_f_Int_Int_Int_Int_goMux1_select_q :
                                                     (call_f_f_Int_Int_Int_Int_goMux1_d[0] ? 5'd1 :
                                                      (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_d[0] ? 5'd2 :
                                                       (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_d[0] ? 5'd4 :
                                                        (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_d[0] ? 5'd8 :
                                                         (lizzieLet13_1_4QNode_Int_1_argbuf_d[0] ? 5'd16 :
                                                          5'd0))))));
  logic [4:0] call_f_f_Int_Int_Int_Int_goMux1_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_Int_Int_Int_goMux1_select_q <= 5'd0;
    else
      call_f_f_Int_Int_Int_Int_goMux1_select_q <= (call_f_f_Int_Int_Int_Int_goMux1_done ? 5'd0 :
                                                   call_f_f_Int_Int_Int_Int_goMux1_select_d);
  logic [1:0] call_f_f_Int_Int_Int_Int_goMux1_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_Int_Int_Int_goMux1_emit_q <= 2'd0;
    else
      call_f_f_Int_Int_Int_Int_goMux1_emit_q <= (call_f_f_Int_Int_Int_Int_goMux1_done ? 2'd0 :
                                                 call_f_f_Int_Int_Int_Int_goMux1_emit_d);
  logic [1:0] call_f_f_Int_Int_Int_Int_goMux1_emit_d;
  assign call_f_f_Int_Int_Int_Int_goMux1_emit_d = (call_f_f_Int_Int_Int_Int_goMux1_emit_q | ({go_12_goMux_choice_d[0],
                                                                                              go_12_goMux_data_d[0]} & {go_12_goMux_choice_r,
                                                                                                                        go_12_goMux_data_r}));
  logic call_f_f_Int_Int_Int_Int_goMux1_done;
  assign call_f_f_Int_Int_Int_Int_goMux1_done = (& call_f_f_Int_Int_Int_Int_goMux1_emit_d);
  assign {lizzieLet13_1_4QNode_Int_1_argbuf_r,
          lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_r,
          lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_r,
          lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux1_r} = (call_f_f_Int_Int_Int_Int_goMux1_done ? call_f_f_Int_Int_Int_Int_goMux1_select_d :
                                                5'd0);
  assign go_12_goMux_data_d = ((call_f_f_Int_Int_Int_Int_goMux1_select_d[0] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[0])) ? call_f_f_Int_Int_Int_Int_goMux1_d :
                               ((call_f_f_Int_Int_Int_Int_goMux1_select_d[1] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_d :
                                ((call_f_f_Int_Int_Int_Int_goMux1_select_d[2] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_d :
                                 ((call_f_f_Int_Int_Int_Int_goMux1_select_d[3] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_d :
                                  ((call_f_f_Int_Int_Int_Int_goMux1_select_d[4] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[0])) ? lizzieLet13_1_4QNode_Int_1_argbuf_d :
                                   1'd0)))));
  assign go_12_goMux_choice_d = ((call_f_f_Int_Int_Int_Int_goMux1_select_d[0] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[1])) ? C1_5_dc(1'd1) :
                                 ((call_f_f_Int_Int_Int_Int_goMux1_select_d[1] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[1])) ? C2_5_dc(1'd1) :
                                  ((call_f_f_Int_Int_Int_Int_goMux1_select_d[2] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[1])) ? C3_5_dc(1'd1) :
                                   ((call_f_f_Int_Int_Int_Int_goMux1_select_d[3] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[1])) ? C4_5_dc(1'd1) :
                                    ((call_f_f_Int_Int_Int_Int_goMux1_select_d[4] && (! call_f_f_Int_Int_Int_Int_goMux1_emit_q[1])) ? C5_5_dc(1'd1) :
                                     {3'd0, 1'd0})))));
  
  /* fork (Ty Go) : (call_f_f_Int_Int_Int_Int_initBuf,Go) > [(call_f_f_Int_Int_Int_Int_unlockFork1,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork2,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork3,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork4,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork5,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork6,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork7,Go),
                                                        (call_f_f_Int_Int_Int_Int_unlockFork8,Go)] */
  logic [7:0] call_f_f_Int_Int_Int_Int_initBuf_emitted;
  logic [7:0] call_f_f_Int_Int_Int_Int_initBuf_done;
  assign call_f_f_Int_Int_Int_Int_unlockFork1_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork2_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[1]));
  assign call_f_f_Int_Int_Int_Int_unlockFork3_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[2]));
  assign call_f_f_Int_Int_Int_Int_unlockFork4_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[3]));
  assign call_f_f_Int_Int_Int_Int_unlockFork5_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[4]));
  assign call_f_f_Int_Int_Int_Int_unlockFork6_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[5]));
  assign call_f_f_Int_Int_Int_Int_unlockFork7_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[6]));
  assign call_f_f_Int_Int_Int_Int_unlockFork8_d = (call_f_f_Int_Int_Int_Int_initBuf_d[0] && (! call_f_f_Int_Int_Int_Int_initBuf_emitted[7]));
  assign call_f_f_Int_Int_Int_Int_initBuf_done = (call_f_f_Int_Int_Int_Int_initBuf_emitted | ({call_f_f_Int_Int_Int_Int_unlockFork8_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork7_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork6_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork5_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork4_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork3_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork2_d[0],
                                                                                               call_f_f_Int_Int_Int_Int_unlockFork1_d[0]} & {call_f_f_Int_Int_Int_Int_unlockFork8_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork7_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork6_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork5_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork4_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork3_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork2_r,
                                                                                                                                             call_f_f_Int_Int_Int_Int_unlockFork1_r}));
  assign call_f_f_Int_Int_Int_Int_initBuf_r = (& call_f_f_Int_Int_Int_Int_initBuf_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_Int_Int_Int_initBuf_emitted <= 8'd0;
    else
      call_f_f_Int_Int_Int_Int_initBuf_emitted <= (call_f_f_Int_Int_Int_Int_initBuf_r ? 8'd0 :
                                                   call_f_f_Int_Int_Int_Int_initBuf_done);
  
  /* initbuf (Ty Go,
         Dcon Go) : (call_f_f_Int_Int_Int_Int_initBufi,Go) > (call_f_f_Int_Int_Int_Int_initBuf,Go) */
  assign call_f_f_Int_Int_Int_Int_initBufi_r = ((! call_f_f_Int_Int_Int_Int_initBuf_d[0]) || call_f_f_Int_Int_Int_Int_initBuf_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      call_f_f_Int_Int_Int_Int_initBuf_d <= Go_dc(1'd1);
    else
      if (call_f_f_Int_Int_Int_Int_initBufi_r)
        call_f_f_Int_Int_Int_Int_initBuf_d <= call_f_f_Int_Int_Int_Int_initBufi_d;
  
  /* mux (Ty Go,
     Ty Go) : (call_f_f_Int_Int_Int_Int_unlockFork1,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12,Go)] > (call_f_f_Int_Int_Int_Int_goMux1,Go) */
  assign call_f_f_Int_Int_Int_Int_goMux1_d = (call_f_f_Int_Int_Int_Int_unlockFork1_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d[0]);
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_r = (call_f_f_Int_Int_Int_Int_goMux1_r && (call_f_f_Int_Int_Int_Int_unlockFork1_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork1_r = (call_f_f_Int_Int_Int_Int_goMux1_r && (call_f_f_Int_Int_Int_Int_unlockFork1_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intgo_12_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_Int_Int_Int_unlockFork2,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU,Pointer_QTree_Int)] > (call_f_f_Int_Int_Int_Int_goMux2,Pointer_QTree_Int) */
  assign call_f_f_Int_Int_Int_Int_goMux2_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d[16:1],
                                              (call_f_f_Int_Int_Int_Int_unlockFork2_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d[0])};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_r = (call_f_f_Int_Int_Int_Int_goMux2_r && (call_f_f_Int_Int_Int_Int_unlockFork2_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork2_r = (call_f_f_Int_Int_Int_Int_goMux2_r && (call_f_f_Int_Int_Int_Int_unlockFork2_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm1ahU_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_QTree_Int) : (call_f_f_Int_Int_Int_Int_unlockFork3,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV,Pointer_QTree_Int)] > (call_f_f_Int_Int_Int_Int_goMux3,Pointer_QTree_Int) */
  assign call_f_f_Int_Int_Int_Int_goMux3_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d[16:1],
                                              (call_f_f_Int_Int_Int_Int_unlockFork3_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d[0])};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_r = (call_f_f_Int_Int_Int_Int_goMux3_r && (call_f_f_Int_Int_Int_Int_unlockFork3_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork3_r = (call_f_f_Int_Int_Int_Int_goMux3_r && (call_f_f_Int_Int_Int_Int_unlockFork3_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intm2ahV_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_Int_Int_Int_unlockFork4,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW,MyDTInt_Bool)] > (call_f_f_Int_Int_Int_Int_goMux4,MyDTInt_Bool) */
  assign call_f_f_Int_Int_Int_Int_goMux4_d = (call_f_f_Int_Int_Int_Int_unlockFork4_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d[0]);
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_r = (call_f_f_Int_Int_Int_Int_goMux4_r && (call_f_f_Int_Int_Int_Int_unlockFork4_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork4_r = (call_f_f_Int_Int_Int_Int_goMux4_r && (call_f_f_Int_Int_Int_Int_unlockFork4_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_kronahW_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int_Int) : (call_f_f_Int_Int_Int_Int_unlockFork5,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX,MyDTInt_Int_Int)] > (call_f_f_Int_Int_Int_Int_goMux5,MyDTInt_Int_Int) */
  assign call_f_f_Int_Int_Int_Int_goMux5_d = (call_f_f_Int_Int_Int_Int_unlockFork5_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d[0]);
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_r = (call_f_f_Int_Int_Int_Int_goMux5_r && (call_f_f_Int_Int_Int_Int_unlockFork5_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork5_r = (call_f_f_Int_Int_Int_Int_goMux5_r && (call_f_f_Int_Int_Int_Int_unlockFork5_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intop_kronahX_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Bool) : (call_f_f_Int_Int_Int_Int_unlockFork6,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY,MyDTInt_Bool)] > (call_f_f_Int_Int_Int_Int_goMux6,MyDTInt_Bool) */
  assign call_f_f_Int_Int_Int_Int_goMux6_d = (call_f_f_Int_Int_Int_Int_unlockFork6_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d[0]);
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_r = (call_f_f_Int_Int_Int_Int_goMux6_r && (call_f_f_Int_Int_Int_Int_unlockFork6_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork6_r = (call_f_f_Int_Int_Int_Int_goMux6_r && (call_f_f_Int_Int_Int_Int_unlockFork6_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intis_z_mapahY_d[0]));
  
  /* mux (Ty Go,
     Ty MyDTInt_Int) : (call_f_f_Int_Int_Int_Int_unlockFork7,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ,MyDTInt_Int)] > (call_f_f_Int_Int_Int_Int_goMux7,MyDTInt_Int) */
  assign call_f_f_Int_Int_Int_Int_goMux7_d = (call_f_f_Int_Int_Int_Int_unlockFork7_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d[0]);
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_r = (call_f_f_Int_Int_Int_Int_goMux7_r && (call_f_f_Int_Int_Int_Int_unlockFork7_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork7_r = (call_f_f_Int_Int_Int_Int_goMux7_r && (call_f_f_Int_Int_Int_Int_unlockFork7_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intf_mapahZ_d[0]));
  
  /* mux (Ty Go,
     Ty Pointer_CTf_f_Int_Int_Int_Int) : (call_f_f_Int_Int_Int_Int_unlockFork8,Go) [(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2,Pointer_CTf_f_Int_Int_Int_Int)] > (call_f_f_Int_Int_Int_Int_goMux8,Pointer_CTf_f_Int_Int_Int_Int) */
  assign call_f_f_Int_Int_Int_Int_goMux8_d = {call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d[16:1],
                                              (call_f_f_Int_Int_Int_Int_unlockFork8_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d[0])};
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_r = (call_f_f_Int_Int_Int_Int_goMux8_r && (call_f_f_Int_Int_Int_Int_unlockFork8_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d[0]));
  assign call_f_f_Int_Int_Int_Int_unlockFork8_r = (call_f_f_Int_Int_Int_Int_goMux8_r && (call_f_f_Int_Int_Int_Int_unlockFork8_d[0] && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Intsc_0_2_d[0]));
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_2_1,MyBool) (lizzieLet6_3QVal_Int,MyDTInt_Int) > [(es_2_1MyFalse,MyDTInt_Int),
                                                                               (_41,MyDTInt_Int)] */
  logic [1:0] lizzieLet6_3QVal_Int_onehotd;
  always_comb
    if ((es_2_1_d[0] && lizzieLet6_3QVal_Int_d[0]))
      unique case (es_2_1_d[1:1])
        1'd0: lizzieLet6_3QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet6_3QVal_Int_onehotd = 2'd2;
        default: lizzieLet6_3QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet6_3QVal_Int_onehotd = 2'd0;
  assign es_2_1MyFalse_d = lizzieLet6_3QVal_Int_onehotd[0];
  assign _41_d = lizzieLet6_3QVal_Int_onehotd[1];
  assign lizzieLet6_3QVal_Int_r = (| (lizzieLet6_3QVal_Int_onehotd & {_41_r,
                                                                      es_2_1MyFalse_r}));
  assign es_2_1_r = lizzieLet6_3QVal_Int_r;
  
  /* fork (Ty MyDTInt_Int) : (es_2_1MyFalse,MyDTInt_Int) > [(es_2_1MyFalse_1,MyDTInt_Int),
                                                       (es_2_1MyFalse_2,MyDTInt_Int)] */
  logic [1:0] es_2_1MyFalse_emitted;
  logic [1:0] es_2_1MyFalse_done;
  assign es_2_1MyFalse_1_d = (es_2_1MyFalse_d[0] && (! es_2_1MyFalse_emitted[0]));
  assign es_2_1MyFalse_2_d = (es_2_1MyFalse_d[0] && (! es_2_1MyFalse_emitted[1]));
  assign es_2_1MyFalse_done = (es_2_1MyFalse_emitted | ({es_2_1MyFalse_2_d[0],
                                                         es_2_1MyFalse_1_d[0]} & {es_2_1MyFalse_2_r,
                                                                                  es_2_1MyFalse_1_r}));
  assign es_2_1MyFalse_r = (& es_2_1MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_emitted <= 2'd0;
    else
      es_2_1MyFalse_emitted <= (es_2_1MyFalse_r ? 2'd0 :
                                es_2_1MyFalse_done);
  
  /* buf (Ty MyDTInt_Int) : (es_2_1MyFalse_1,MyDTInt_Int) > (es_2_1MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_2_1MyFalse_1_bufchan_d;
  logic es_2_1MyFalse_1_bufchan_r;
  assign es_2_1MyFalse_1_r = ((! es_2_1MyFalse_1_bufchan_d[0]) || es_2_1MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_2_1MyFalse_1_r)
        es_2_1MyFalse_1_bufchan_d <= es_2_1MyFalse_1_d;
  MyDTInt_Int_t es_2_1MyFalse_1_bufchan_buf;
  assign es_2_1MyFalse_1_bufchan_r = (! es_2_1MyFalse_1_bufchan_buf[0]);
  assign es_2_1MyFalse_1_argbuf_d = (es_2_1MyFalse_1_bufchan_buf[0] ? es_2_1MyFalse_1_bufchan_buf :
                                     es_2_1MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_1MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_2_1MyFalse_1_argbuf_r && es_2_1MyFalse_1_bufchan_buf[0]))
        es_2_1MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_2_1MyFalse_1_argbuf_r) && (! es_2_1MyFalse_1_bufchan_buf[0])))
        es_2_1MyFalse_1_bufchan_buf <= es_2_1MyFalse_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_2_2,MyBool) (lizzieLet6_4QVal_Int_2,Go) > [(es_2_2MyFalse,Go),
                                                               (es_2_2MyTrue,Go)] */
  logic [1:0] lizzieLet6_4QVal_Int_2_onehotd;
  always_comb
    if ((es_2_2_d[0] && lizzieLet6_4QVal_Int_2_d[0]))
      unique case (es_2_2_d[1:1])
        1'd0: lizzieLet6_4QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_4QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_4QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_4QVal_Int_2_onehotd = 2'd0;
  assign es_2_2MyFalse_d = lizzieLet6_4QVal_Int_2_onehotd[0];
  assign es_2_2MyTrue_d = lizzieLet6_4QVal_Int_2_onehotd[1];
  assign lizzieLet6_4QVal_Int_2_r = (| (lizzieLet6_4QVal_Int_2_onehotd & {es_2_2MyTrue_r,
                                                                          es_2_2MyFalse_r}));
  assign es_2_2_r = lizzieLet6_4QVal_Int_2_r;
  
  /* fork (Ty Go) : (es_2_2MyFalse,Go) > [(es_2_2MyFalse_1,Go),
                                     (es_2_2MyFalse_2,Go),
                                     (es_2_2MyFalse_3,Go)] */
  logic [2:0] es_2_2MyFalse_emitted;
  logic [2:0] es_2_2MyFalse_done;
  assign es_2_2MyFalse_1_d = (es_2_2MyFalse_d[0] && (! es_2_2MyFalse_emitted[0]));
  assign es_2_2MyFalse_2_d = (es_2_2MyFalse_d[0] && (! es_2_2MyFalse_emitted[1]));
  assign es_2_2MyFalse_3_d = (es_2_2MyFalse_d[0] && (! es_2_2MyFalse_emitted[2]));
  assign es_2_2MyFalse_done = (es_2_2MyFalse_emitted | ({es_2_2MyFalse_3_d[0],
                                                         es_2_2MyFalse_2_d[0],
                                                         es_2_2MyFalse_1_d[0]} & {es_2_2MyFalse_3_r,
                                                                                  es_2_2MyFalse_2_r,
                                                                                  es_2_2MyFalse_1_r}));
  assign es_2_2MyFalse_r = (& es_2_2MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_emitted <= 3'd0;
    else
      es_2_2MyFalse_emitted <= (es_2_2MyFalse_r ? 3'd0 :
                                es_2_2MyFalse_done);
  
  /* buf (Ty Go) : (es_2_2MyFalse_1,Go) > (es_2_2MyFalse_1_argbuf,Go) */
  Go_t es_2_2MyFalse_1_bufchan_d;
  logic es_2_2MyFalse_1_bufchan_r;
  assign es_2_2MyFalse_1_r = ((! es_2_2MyFalse_1_bufchan_d[0]) || es_2_2MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_2_2MyFalse_1_r)
        es_2_2MyFalse_1_bufchan_d <= es_2_2MyFalse_1_d;
  Go_t es_2_2MyFalse_1_bufchan_buf;
  assign es_2_2MyFalse_1_bufchan_r = (! es_2_2MyFalse_1_bufchan_buf[0]);
  assign es_2_2MyFalse_1_argbuf_d = (es_2_2MyFalse_1_bufchan_buf[0] ? es_2_2MyFalse_1_bufchan_buf :
                                     es_2_2MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyFalse_1_argbuf_r && es_2_2MyFalse_1_bufchan_buf[0]))
        es_2_2MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyFalse_1_argbuf_r) && (! es_2_2MyFalse_1_bufchan_buf[0])))
        es_2_2MyFalse_1_bufchan_buf <= es_2_2MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_2_2MyFalse_1_argbuf,Go),
                                         (es_2_1MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_6_1_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d = TupGo___MyDTInt_Int___Int_dc((& {es_2_2MyFalse_1_argbuf_d[0],
                                                                                          es_2_1MyFalse_1_argbuf_d[0],
                                                                                          es_6_1_1_argbuf_d[0]}), es_2_2MyFalse_1_argbuf_d, es_2_1MyFalse_1_argbuf_d, es_6_1_1_argbuf_d);
  assign {es_2_2MyFalse_1_argbuf_r,
          es_2_1MyFalse_1_argbuf_r,
          es_6_1_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int_1_d[0])}};
  
  /* buf (Ty Go) : (es_2_2MyFalse_2,Go) > (es_2_2MyFalse_2_argbuf,Go) */
  Go_t es_2_2MyFalse_2_bufchan_d;
  logic es_2_2MyFalse_2_bufchan_r;
  assign es_2_2MyFalse_2_r = ((! es_2_2MyFalse_2_bufchan_d[0]) || es_2_2MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_2_2MyFalse_2_r)
        es_2_2MyFalse_2_bufchan_d <= es_2_2MyFalse_2_d;
  Go_t es_2_2MyFalse_2_bufchan_buf;
  assign es_2_2MyFalse_2_bufchan_r = (! es_2_2MyFalse_2_bufchan_buf[0]);
  assign es_2_2MyFalse_2_argbuf_d = (es_2_2MyFalse_2_bufchan_buf[0] ? es_2_2MyFalse_2_bufchan_buf :
                                     es_2_2MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyFalse_2_argbuf_r && es_2_2MyFalse_2_bufchan_buf[0]))
        es_2_2MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyFalse_2_argbuf_r) && (! es_2_2MyFalse_2_bufchan_buf[0])))
        es_2_2MyFalse_2_bufchan_buf <= es_2_2MyFalse_2_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(es_2_2MyFalse_2_argbuf,Go),
                                          (es_2_3MyFalse_1_argbuf,MyDTInt_Bool),
                                          (es_4_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d = TupGo___MyDTInt_Bool___Int_dc((& {es_2_2MyFalse_2_argbuf_d[0],
                                                                                            es_2_3MyFalse_1_argbuf_d[0],
                                                                                            es_4_1_1_argbuf_d[0]}), es_2_2MyFalse_2_argbuf_d, es_2_3MyFalse_1_argbuf_d, es_4_1_1_argbuf_d);
  assign {es_2_2MyFalse_2_argbuf_r,
          es_2_3MyFalse_1_argbuf_r,
          es_4_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int2_d[0])}};
  
  /* fork (Ty Go) : (es_2_2MyTrue,Go) > [(es_2_2MyTrue_1,Go),
                                    (es_2_2MyTrue_2,Go)] */
  logic [1:0] es_2_2MyTrue_emitted;
  logic [1:0] es_2_2MyTrue_done;
  assign es_2_2MyTrue_1_d = (es_2_2MyTrue_d[0] && (! es_2_2MyTrue_emitted[0]));
  assign es_2_2MyTrue_2_d = (es_2_2MyTrue_d[0] && (! es_2_2MyTrue_emitted[1]));
  assign es_2_2MyTrue_done = (es_2_2MyTrue_emitted | ({es_2_2MyTrue_2_d[0],
                                                       es_2_2MyTrue_1_d[0]} & {es_2_2MyTrue_2_r,
                                                                               es_2_2MyTrue_1_r}));
  assign es_2_2MyTrue_r = (& es_2_2MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyTrue_emitted <= 2'd0;
    else
      es_2_2MyTrue_emitted <= (es_2_2MyTrue_r ? 2'd0 :
                               es_2_2MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_2_2MyTrue_1,Go)] > (es_2_2MyTrue_1QNone_Int,QTree_Int) */
  assign es_2_2MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_2_2MyTrue_1_d[0]}), es_2_2MyTrue_1_d);
  assign {es_2_2MyTrue_1_r} = {1 {(es_2_2MyTrue_1QNone_Int_r && es_2_2MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_2_2MyTrue_1QNone_Int,QTree_Int) > (lizzieLet10_1_argbuf,QTree_Int) */
  QTree_Int_t es_2_2MyTrue_1QNone_Int_bufchan_d;
  logic es_2_2MyTrue_1QNone_Int_bufchan_r;
  assign es_2_2MyTrue_1QNone_Int_r = ((! es_2_2MyTrue_1QNone_Int_bufchan_d[0]) || es_2_2MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_2MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_2_2MyTrue_1QNone_Int_r)
        es_2_2MyTrue_1QNone_Int_bufchan_d <= es_2_2MyTrue_1QNone_Int_d;
  QTree_Int_t es_2_2MyTrue_1QNone_Int_bufchan_buf;
  assign es_2_2MyTrue_1QNone_Int_bufchan_r = (! es_2_2MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet10_1_argbuf_d = (es_2_2MyTrue_1QNone_Int_bufchan_buf[0] ? es_2_2MyTrue_1QNone_Int_bufchan_buf :
                                   es_2_2MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_2_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet10_1_argbuf_r && es_2_2MyTrue_1QNone_Int_bufchan_buf[0]))
        es_2_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet10_1_argbuf_r) && (! es_2_2MyTrue_1QNone_Int_bufchan_buf[0])))
        es_2_2MyTrue_1QNone_Int_bufchan_buf <= es_2_2MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_2_2MyTrue_2,Go) > (es_2_2MyTrue_2_argbuf,Go) */
  Go_t es_2_2MyTrue_2_bufchan_d;
  logic es_2_2MyTrue_2_bufchan_r;
  assign es_2_2MyTrue_2_r = ((! es_2_2MyTrue_2_bufchan_d[0]) || es_2_2MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_2_2MyTrue_2_r) es_2_2MyTrue_2_bufchan_d <= es_2_2MyTrue_2_d;
  Go_t es_2_2MyTrue_2_bufchan_buf;
  assign es_2_2MyTrue_2_bufchan_r = (! es_2_2MyTrue_2_bufchan_buf[0]);
  assign es_2_2MyTrue_2_argbuf_d = (es_2_2MyTrue_2_bufchan_buf[0] ? es_2_2MyTrue_2_bufchan_buf :
                                    es_2_2MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_2MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_2_2MyTrue_2_argbuf_r && es_2_2MyTrue_2_bufchan_buf[0]))
        es_2_2MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_2_2MyTrue_2_argbuf_r) && (! es_2_2MyTrue_2_bufchan_buf[0])))
        es_2_2MyTrue_2_bufchan_buf <= es_2_2MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Bool) : (es_2_3,MyBool) (lizzieLet6_6QVal_Int,MyDTInt_Bool) > [(es_2_3MyFalse,MyDTInt_Bool),
                                                                                 (_40,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_6QVal_Int_onehotd;
  always_comb
    if ((es_2_3_d[0] && lizzieLet6_6QVal_Int_d[0]))
      unique case (es_2_3_d[1:1])
        1'd0: lizzieLet6_6QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet6_6QVal_Int_onehotd = 2'd2;
        default: lizzieLet6_6QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet6_6QVal_Int_onehotd = 2'd0;
  assign es_2_3MyFalse_d = lizzieLet6_6QVal_Int_onehotd[0];
  assign _40_d = lizzieLet6_6QVal_Int_onehotd[1];
  assign lizzieLet6_6QVal_Int_r = (| (lizzieLet6_6QVal_Int_onehotd & {_40_r,
                                                                      es_2_3MyFalse_r}));
  assign es_2_3_r = lizzieLet6_6QVal_Int_r;
  
  /* buf (Ty MyDTInt_Bool) : (es_2_3MyFalse,MyDTInt_Bool) > (es_2_3MyFalse_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t es_2_3MyFalse_bufchan_d;
  logic es_2_3MyFalse_bufchan_r;
  assign es_2_3MyFalse_r = ((! es_2_3MyFalse_bufchan_d[0]) || es_2_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_d <= 1'd0;
    else
      if (es_2_3MyFalse_r) es_2_3MyFalse_bufchan_d <= es_2_3MyFalse_d;
  MyDTInt_Bool_t es_2_3MyFalse_bufchan_buf;
  assign es_2_3MyFalse_bufchan_r = (! es_2_3MyFalse_bufchan_buf[0]);
  assign es_2_3MyFalse_1_argbuf_d = (es_2_3MyFalse_bufchan_buf[0] ? es_2_3MyFalse_bufchan_buf :
                                     es_2_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_3MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_2_3MyFalse_1_argbuf_r && es_2_3MyFalse_bufchan_buf[0]))
        es_2_3MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_2_3MyFalse_1_argbuf_r) && (! es_2_3MyFalse_bufchan_buf[0])))
        es_2_3MyFalse_bufchan_buf <= es_2_3MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_2_4,MyBool) (lizzieLet6_7QVal_Int_2,MyDTInt_Int_Int) > [(es_2_4MyFalse,MyDTInt_Int_Int),
                                                                                         (_39,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_7QVal_Int_2_onehotd;
  always_comb
    if ((es_2_4_d[0] && lizzieLet6_7QVal_Int_2_d[0]))
      unique case (es_2_4_d[1:1])
        1'd0: lizzieLet6_7QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_7QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_7QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_7QVal_Int_2_onehotd = 2'd0;
  assign es_2_4MyFalse_d = lizzieLet6_7QVal_Int_2_onehotd[0];
  assign _39_d = lizzieLet6_7QVal_Int_2_onehotd[1];
  assign lizzieLet6_7QVal_Int_2_r = (| (lizzieLet6_7QVal_Int_2_onehotd & {_39_r,
                                                                          es_2_4MyFalse_r}));
  assign es_2_4_r = lizzieLet6_7QVal_Int_2_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (es_2_4MyFalse,MyDTInt_Int_Int) > [(es_2_4MyFalse_1,MyDTInt_Int_Int),
                                                               (es_2_4MyFalse_2,MyDTInt_Int_Int)] */
  logic [1:0] es_2_4MyFalse_emitted;
  logic [1:0] es_2_4MyFalse_done;
  assign es_2_4MyFalse_1_d = (es_2_4MyFalse_d[0] && (! es_2_4MyFalse_emitted[0]));
  assign es_2_4MyFalse_2_d = (es_2_4MyFalse_d[0] && (! es_2_4MyFalse_emitted[1]));
  assign es_2_4MyFalse_done = (es_2_4MyFalse_emitted | ({es_2_4MyFalse_2_d[0],
                                                         es_2_4MyFalse_1_d[0]} & {es_2_4MyFalse_2_r,
                                                                                  es_2_4MyFalse_1_r}));
  assign es_2_4MyFalse_r = (& es_2_4MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_emitted <= 2'd0;
    else
      es_2_4MyFalse_emitted <= (es_2_4MyFalse_r ? 2'd0 :
                                es_2_4MyFalse_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (es_2_4MyFalse_1,MyDTInt_Int_Int) > (es_2_4MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_2_4MyFalse_1_bufchan_d;
  logic es_2_4MyFalse_1_bufchan_r;
  assign es_2_4MyFalse_1_r = ((! es_2_4MyFalse_1_bufchan_d[0]) || es_2_4MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_2_4MyFalse_1_r)
        es_2_4MyFalse_1_bufchan_d <= es_2_4MyFalse_1_d;
  MyDTInt_Int_Int_t es_2_4MyFalse_1_bufchan_buf;
  assign es_2_4MyFalse_1_bufchan_r = (! es_2_4MyFalse_1_bufchan_buf[0]);
  assign es_2_4MyFalse_1_argbuf_d = (es_2_4MyFalse_1_bufchan_buf[0] ? es_2_4MyFalse_1_bufchan_buf :
                                     es_2_4MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_4MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_2_4MyFalse_1_argbuf_r && es_2_4MyFalse_1_bufchan_buf[0]))
        es_2_4MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_2_4MyFalse_1_argbuf_r) && (! es_2_4MyFalse_1_bufchan_buf[0])))
        es_2_4MyFalse_1_bufchan_buf <= es_2_4MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_2_4MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_2_6MyFalse_1_argbuf,Int),
                                              (es_2_7MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_2_4MyFalse_1_argbuf_d[0],
                                                                                                       es_2_6MyFalse_1_argbuf_d[0],
                                                                                                       es_2_7MyFalse_1_argbuf_d[0]}), es_2_4MyFalse_1_argbuf_d, es_2_6MyFalse_1_argbuf_d, es_2_7MyFalse_1_argbuf_d);
  assign {es_2_4MyFalse_1_argbuf_r,
          es_2_6MyFalse_1_argbuf_r,
          es_2_7MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int2_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (es_2_5,MyBool) (lizzieLet6_8QVal_Int,Pointer_CTf'_f'_Int_Int_Int_Int) > [(es_2_5MyFalse,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                       (es_2_5MyTrue,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [1:0] lizzieLet6_8QVal_Int_onehotd;
  always_comb
    if ((es_2_5_d[0] && lizzieLet6_8QVal_Int_d[0]))
      unique case (es_2_5_d[1:1])
        1'd0: lizzieLet6_8QVal_Int_onehotd = 2'd1;
        1'd1: lizzieLet6_8QVal_Int_onehotd = 2'd2;
        default: lizzieLet6_8QVal_Int_onehotd = 2'd0;
      endcase
    else lizzieLet6_8QVal_Int_onehotd = 2'd0;
  assign es_2_5MyFalse_d = {lizzieLet6_8QVal_Int_d[16:1],
                            lizzieLet6_8QVal_Int_onehotd[0]};
  assign es_2_5MyTrue_d = {lizzieLet6_8QVal_Int_d[16:1],
                           lizzieLet6_8QVal_Int_onehotd[1]};
  assign lizzieLet6_8QVal_Int_r = (| (lizzieLet6_8QVal_Int_onehotd & {es_2_5MyTrue_r,
                                                                      es_2_5MyFalse_r}));
  assign es_2_5_r = lizzieLet6_8QVal_Int_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (es_2_5MyTrue,Pointer_CTf'_f'_Int_Int_Int_Int) > (es_2_5MyTrue_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_2_5MyTrue_bufchan_d;
  logic es_2_5MyTrue_bufchan_r;
  assign es_2_5MyTrue_r = ((! es_2_5MyTrue_bufchan_d[0]) || es_2_5MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyTrue_bufchan_d <= {16'd0, 1'd0};
    else if (es_2_5MyTrue_r) es_2_5MyTrue_bufchan_d <= es_2_5MyTrue_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_2_5MyTrue_bufchan_buf;
  assign es_2_5MyTrue_bufchan_r = (! es_2_5MyTrue_bufchan_buf[0]);
  assign es_2_5MyTrue_1_argbuf_d = (es_2_5MyTrue_bufchan_buf[0] ? es_2_5MyTrue_bufchan_buf :
                                    es_2_5MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_5MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_2_5MyTrue_1_argbuf_r && es_2_5MyTrue_bufchan_buf[0]))
        es_2_5MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_2_5MyTrue_1_argbuf_r) && (! es_2_5MyTrue_bufchan_buf[0])))
        es_2_5MyTrue_bufchan_buf <= es_2_5MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_6,MyBool) (lizzieLet6_9QVal_Int_2,Int) > [(es_2_6MyFalse,Int),
                                                                 (_38,Int)] */
  logic [1:0] lizzieLet6_9QVal_Int_2_onehotd;
  always_comb
    if ((es_2_6_d[0] && lizzieLet6_9QVal_Int_2_d[0]))
      unique case (es_2_6_d[1:1])
        1'd0: lizzieLet6_9QVal_Int_2_onehotd = 2'd1;
        1'd1: lizzieLet6_9QVal_Int_2_onehotd = 2'd2;
        default: lizzieLet6_9QVal_Int_2_onehotd = 2'd0;
      endcase
    else lizzieLet6_9QVal_Int_2_onehotd = 2'd0;
  assign es_2_6MyFalse_d = {lizzieLet6_9QVal_Int_2_d[32:1],
                            lizzieLet6_9QVal_Int_2_onehotd[0]};
  assign _38_d = {lizzieLet6_9QVal_Int_2_d[32:1],
                  lizzieLet6_9QVal_Int_2_onehotd[1]};
  assign lizzieLet6_9QVal_Int_2_r = (| (lizzieLet6_9QVal_Int_2_onehotd & {_38_r,
                                                                          es_2_6MyFalse_r}));
  assign es_2_6_r = lizzieLet6_9QVal_Int_2_r;
  
  /* fork (Ty Int) : (es_2_6MyFalse,Int) > [(es_2_6MyFalse_1,Int),
                                       (es_2_6MyFalse_2,Int)] */
  logic [1:0] es_2_6MyFalse_emitted;
  logic [1:0] es_2_6MyFalse_done;
  assign es_2_6MyFalse_1_d = {es_2_6MyFalse_d[32:1],
                              (es_2_6MyFalse_d[0] && (! es_2_6MyFalse_emitted[0]))};
  assign es_2_6MyFalse_2_d = {es_2_6MyFalse_d[32:1],
                              (es_2_6MyFalse_d[0] && (! es_2_6MyFalse_emitted[1]))};
  assign es_2_6MyFalse_done = (es_2_6MyFalse_emitted | ({es_2_6MyFalse_2_d[0],
                                                         es_2_6MyFalse_1_d[0]} & {es_2_6MyFalse_2_r,
                                                                                  es_2_6MyFalse_1_r}));
  assign es_2_6MyFalse_r = (& es_2_6MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_6MyFalse_emitted <= 2'd0;
    else
      es_2_6MyFalse_emitted <= (es_2_6MyFalse_r ? 2'd0 :
                                es_2_6MyFalse_done);
  
  /* buf (Ty Int) : (es_2_6MyFalse_1,Int) > (es_2_6MyFalse_1_argbuf,Int) */
  Int_t es_2_6MyFalse_1_bufchan_d;
  logic es_2_6MyFalse_1_bufchan_r;
  assign es_2_6MyFalse_1_r = ((! es_2_6MyFalse_1_bufchan_d[0]) || es_2_6MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_6MyFalse_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_6MyFalse_1_r)
        es_2_6MyFalse_1_bufchan_d <= es_2_6MyFalse_1_d;
  Int_t es_2_6MyFalse_1_bufchan_buf;
  assign es_2_6MyFalse_1_bufchan_r = (! es_2_6MyFalse_1_bufchan_buf[0]);
  assign es_2_6MyFalse_1_argbuf_d = (es_2_6MyFalse_1_bufchan_buf[0] ? es_2_6MyFalse_1_bufchan_buf :
                                     es_2_6MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_6MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_6MyFalse_1_argbuf_r && es_2_6MyFalse_1_bufchan_buf[0]))
        es_2_6MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_6MyFalse_1_argbuf_r) && (! es_2_6MyFalse_1_bufchan_buf[0])))
        es_2_6MyFalse_1_bufchan_buf <= es_2_6MyFalse_1_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_2_7,MyBool) (v'aib_2,Int) > [(es_2_7MyFalse,Int),
                                                  (_37,Int)] */
  logic [1:0] \v'aib_2_onehotd ;
  always_comb
    if ((es_2_7_d[0] && \v'aib_2_d [0]))
      unique case (es_2_7_d[1:1])
        1'd0: \v'aib_2_onehotd  = 2'd1;
        1'd1: \v'aib_2_onehotd  = 2'd2;
        default: \v'aib_2_onehotd  = 2'd0;
      endcase
    else \v'aib_2_onehotd  = 2'd0;
  assign es_2_7MyFalse_d = {\v'aib_2_d [32:1], \v'aib_2_onehotd [0]};
  assign _37_d = {\v'aib_2_d [32:1], \v'aib_2_onehotd [1]};
  assign \v'aib_2_r  = (| (\v'aib_2_onehotd  & {_37_r,
                                                es_2_7MyFalse_r}));
  assign es_2_7_r = \v'aib_2_r ;
  
  /* fork (Ty Int) : (es_2_7MyFalse,Int) > [(es_2_7MyFalse_1,Int),
                                       (es_2_7MyFalse_2,Int)] */
  logic [1:0] es_2_7MyFalse_emitted;
  logic [1:0] es_2_7MyFalse_done;
  assign es_2_7MyFalse_1_d = {es_2_7MyFalse_d[32:1],
                              (es_2_7MyFalse_d[0] && (! es_2_7MyFalse_emitted[0]))};
  assign es_2_7MyFalse_2_d = {es_2_7MyFalse_d[32:1],
                              (es_2_7MyFalse_d[0] && (! es_2_7MyFalse_emitted[1]))};
  assign es_2_7MyFalse_done = (es_2_7MyFalse_emitted | ({es_2_7MyFalse_2_d[0],
                                                         es_2_7MyFalse_1_d[0]} & {es_2_7MyFalse_2_r,
                                                                                  es_2_7MyFalse_1_r}));
  assign es_2_7MyFalse_r = (& es_2_7MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_7MyFalse_emitted <= 2'd0;
    else
      es_2_7MyFalse_emitted <= (es_2_7MyFalse_r ? 2'd0 :
                                es_2_7MyFalse_done);
  
  /* buf (Ty Int) : (es_2_7MyFalse_1,Int) > (es_2_7MyFalse_1_argbuf,Int) */
  Int_t es_2_7MyFalse_1_bufchan_d;
  logic es_2_7MyFalse_1_bufchan_r;
  assign es_2_7MyFalse_1_r = ((! es_2_7MyFalse_1_bufchan_d[0]) || es_2_7MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_7MyFalse_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_2_7MyFalse_1_r)
        es_2_7MyFalse_1_bufchan_d <= es_2_7MyFalse_1_d;
  Int_t es_2_7MyFalse_1_bufchan_buf;
  assign es_2_7MyFalse_1_bufchan_r = (! es_2_7MyFalse_1_bufchan_buf[0]);
  assign es_2_7MyFalse_1_argbuf_d = (es_2_7MyFalse_1_bufchan_buf[0] ? es_2_7MyFalse_1_bufchan_buf :
                                     es_2_7MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_2_7MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_2_7MyFalse_1_argbuf_r && es_2_7MyFalse_1_bufchan_buf[0]))
        es_2_7MyFalse_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_2_7MyFalse_1_argbuf_r) && (! es_2_7MyFalse_1_bufchan_buf[0])))
        es_2_7MyFalse_1_bufchan_buf <= es_2_7MyFalse_1_bufchan_d;
  
  /* buf (Ty Int#) : (es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32,Int#) > (contRet_0_1_argbuf,Int#) */
  \Int#_t  es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  logic es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_r;
  assign es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_r = ((! es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d[0]) || es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= {32'd0,
                                                                  1'd0};
    else
      if (es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_r)
        es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d <= es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_d;
  \Int#_t  es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf;
  assign es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_r = (! es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]);
  assign contRet_0_1_argbuf_d = (es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0] ? es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf :
                                 es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                    1'd0};
    else
      if ((contRet_0_1_argbuf_r && es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0]))
        es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= {32'd0,
                                                                      1'd0};
      else if (((! contRet_0_1_argbuf_r) && (! es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf[0])))
        es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_buf <= es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_bufchan_d;
  
  /* op_add (Ty Int#) : (es_6_2_1ww2XuO_1_1_Add32,Int#) (lizzieLet19_4Lcall_$wnnz_Int0,Int#) > (es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32,Int#) */
  assign es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_d = {(es_6_2_1ww2XuO_1_1_Add32_d[32:1] + lizzieLet19_4Lcall_$wnnz_Int0_d[32:1]),
                                                            (es_6_2_1ww2XuO_1_1_Add32_d[0] && lizzieLet19_4Lcall_$wnnz_Int0_d[0])};
  assign {es_6_2_1ww2XuO_1_1_Add32_r,
          lizzieLet19_4Lcall_$wnnz_Int0_r} = {2 {(es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_r && es_4_2_1lizzieLet19_4Lcall_$wnnz_Int0_1_Add32_d[0])}};
  
  /* sink (Ty Int) : (es_7_1I#,Int) > */
  assign {\es_7_1I#_r , \es_7_1I#_dout } = {\es_7_1I#_rout ,
                                            \es_7_1I#_d };
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int) : (es_7_1_1,MyBool) (es_2_1MyFalse_2,MyDTInt_Int) > [(es_7_1_1MyFalse,MyDTInt_Int),
                                                                            (_36,MyDTInt_Int)] */
  logic [1:0] es_2_1MyFalse_2_onehotd;
  always_comb
    if ((es_7_1_1_d[0] && es_2_1MyFalse_2_d[0]))
      unique case (es_7_1_1_d[1:1])
        1'd0: es_2_1MyFalse_2_onehotd = 2'd1;
        1'd1: es_2_1MyFalse_2_onehotd = 2'd2;
        default: es_2_1MyFalse_2_onehotd = 2'd0;
      endcase
    else es_2_1MyFalse_2_onehotd = 2'd0;
  assign es_7_1_1MyFalse_d = es_2_1MyFalse_2_onehotd[0];
  assign _36_d = es_2_1MyFalse_2_onehotd[1];
  assign es_2_1MyFalse_2_r = (| (es_2_1MyFalse_2_onehotd & {_36_r,
                                                            es_7_1_1MyFalse_r}));
  assign es_7_1_1_r = es_2_1MyFalse_2_r;
  
  /* buf (Ty MyDTInt_Int) : (es_7_1_1MyFalse,MyDTInt_Int) > (es_7_1_1MyFalse_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t es_7_1_1MyFalse_bufchan_d;
  logic es_7_1_1MyFalse_bufchan_r;
  assign es_7_1_1MyFalse_r = ((! es_7_1_1MyFalse_bufchan_d[0]) || es_7_1_1MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_1MyFalse_bufchan_d <= 1'd0;
    else
      if (es_7_1_1MyFalse_r)
        es_7_1_1MyFalse_bufchan_d <= es_7_1_1MyFalse_d;
  MyDTInt_Int_t es_7_1_1MyFalse_bufchan_buf;
  assign es_7_1_1MyFalse_bufchan_r = (! es_7_1_1MyFalse_bufchan_buf[0]);
  assign es_7_1_1MyFalse_1_argbuf_d = (es_7_1_1MyFalse_bufchan_buf[0] ? es_7_1_1MyFalse_bufchan_buf :
                                       es_7_1_1MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_1MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_7_1_1MyFalse_1_argbuf_r && es_7_1_1MyFalse_bufchan_buf[0]))
        es_7_1_1MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_7_1_1MyFalse_1_argbuf_r) && (! es_7_1_1MyFalse_bufchan_buf[0])))
        es_7_1_1MyFalse_bufchan_buf <= es_7_1_1MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (es_7_1_2,MyBool) (es_2_2MyFalse_3,Go) > [(es_7_1_2MyFalse,Go),
                                                          (es_7_1_2MyTrue,Go)] */
  logic [1:0] es_2_2MyFalse_3_onehotd;
  always_comb
    if ((es_7_1_2_d[0] && es_2_2MyFalse_3_d[0]))
      unique case (es_7_1_2_d[1:1])
        1'd0: es_2_2MyFalse_3_onehotd = 2'd1;
        1'd1: es_2_2MyFalse_3_onehotd = 2'd2;
        default: es_2_2MyFalse_3_onehotd = 2'd0;
      endcase
    else es_2_2MyFalse_3_onehotd = 2'd0;
  assign es_7_1_2MyFalse_d = es_2_2MyFalse_3_onehotd[0];
  assign es_7_1_2MyTrue_d = es_2_2MyFalse_3_onehotd[1];
  assign es_2_2MyFalse_3_r = (| (es_2_2MyFalse_3_onehotd & {es_7_1_2MyTrue_r,
                                                            es_7_1_2MyFalse_r}));
  assign es_7_1_2_r = es_2_2MyFalse_3_r;
  
  /* fork (Ty Go) : (es_7_1_2MyFalse,Go) > [(es_7_1_2MyFalse_1,Go),
                                       (es_7_1_2MyFalse_2,Go)] */
  logic [1:0] es_7_1_2MyFalse_emitted;
  logic [1:0] es_7_1_2MyFalse_done;
  assign es_7_1_2MyFalse_1_d = (es_7_1_2MyFalse_d[0] && (! es_7_1_2MyFalse_emitted[0]));
  assign es_7_1_2MyFalse_2_d = (es_7_1_2MyFalse_d[0] && (! es_7_1_2MyFalse_emitted[1]));
  assign es_7_1_2MyFalse_done = (es_7_1_2MyFalse_emitted | ({es_7_1_2MyFalse_2_d[0],
                                                             es_7_1_2MyFalse_1_d[0]} & {es_7_1_2MyFalse_2_r,
                                                                                        es_7_1_2MyFalse_1_r}));
  assign es_7_1_2MyFalse_r = (& es_7_1_2MyFalse_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyFalse_emitted <= 2'd0;
    else
      es_7_1_2MyFalse_emitted <= (es_7_1_2MyFalse_r ? 2'd0 :
                                  es_7_1_2MyFalse_done);
  
  /* buf (Ty Go) : (es_7_1_2MyFalse_1,Go) > (es_7_1_2MyFalse_1_argbuf,Go) */
  Go_t es_7_1_2MyFalse_1_bufchan_d;
  logic es_7_1_2MyFalse_1_bufchan_r;
  assign es_7_1_2MyFalse_1_r = ((! es_7_1_2MyFalse_1_bufchan_d[0]) || es_7_1_2MyFalse_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyFalse_1_bufchan_d <= 1'd0;
    else
      if (es_7_1_2MyFalse_1_r)
        es_7_1_2MyFalse_1_bufchan_d <= es_7_1_2MyFalse_1_d;
  Go_t es_7_1_2MyFalse_1_bufchan_buf;
  assign es_7_1_2MyFalse_1_bufchan_r = (! es_7_1_2MyFalse_1_bufchan_buf[0]);
  assign es_7_1_2MyFalse_1_argbuf_d = (es_7_1_2MyFalse_1_bufchan_buf[0] ? es_7_1_2MyFalse_1_bufchan_buf :
                                       es_7_1_2MyFalse_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyFalse_1_bufchan_buf <= 1'd0;
    else
      if ((es_7_1_2MyFalse_1_argbuf_r && es_7_1_2MyFalse_1_bufchan_buf[0]))
        es_7_1_2MyFalse_1_bufchan_buf <= 1'd0;
      else if (((! es_7_1_2MyFalse_1_argbuf_r) && (! es_7_1_2MyFalse_1_bufchan_buf[0])))
        es_7_1_2MyFalse_1_bufchan_buf <= es_7_1_2MyFalse_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Int___Int,
      Dcon TupGo___MyDTInt_Int___Int) : [(es_7_1_2MyFalse_1_argbuf,Go),
                                         (es_7_1_1MyFalse_1_argbuf,MyDTInt_Int),
                                         (es_10_1_argbuf,Int)] > (applyfnInt_Int_5TupGo___MyDTInt_Int___Int2,TupGo___MyDTInt_Int___Int) */
  assign applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d = TupGo___MyDTInt_Int___Int_dc((& {es_7_1_2MyFalse_1_argbuf_d[0],
                                                                                         es_7_1_1MyFalse_1_argbuf_d[0],
                                                                                         es_10_1_argbuf_d[0]}), es_7_1_2MyFalse_1_argbuf_d, es_7_1_1MyFalse_1_argbuf_d, es_10_1_argbuf_d);
  assign {es_7_1_2MyFalse_1_argbuf_r,
          es_7_1_1MyFalse_1_argbuf_r,
          es_10_1_argbuf_r} = {3 {(applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_r && applyfnInt_Int_5TupGo___MyDTInt_Int___Int2_d[0])}};
  
  /* buf (Ty Go) : (es_7_1_2MyFalse_2,Go) > (es_7_1_2MyFalse_2_argbuf,Go) */
  Go_t es_7_1_2MyFalse_2_bufchan_d;
  logic es_7_1_2MyFalse_2_bufchan_r;
  assign es_7_1_2MyFalse_2_r = ((! es_7_1_2MyFalse_2_bufchan_d[0]) || es_7_1_2MyFalse_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyFalse_2_bufchan_d <= 1'd0;
    else
      if (es_7_1_2MyFalse_2_r)
        es_7_1_2MyFalse_2_bufchan_d <= es_7_1_2MyFalse_2_d;
  Go_t es_7_1_2MyFalse_2_bufchan_buf;
  assign es_7_1_2MyFalse_2_bufchan_r = (! es_7_1_2MyFalse_2_bufchan_buf[0]);
  assign es_7_1_2MyFalse_2_argbuf_d = (es_7_1_2MyFalse_2_bufchan_buf[0] ? es_7_1_2MyFalse_2_bufchan_buf :
                                       es_7_1_2MyFalse_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyFalse_2_bufchan_buf <= 1'd0;
    else
      if ((es_7_1_2MyFalse_2_argbuf_r && es_7_1_2MyFalse_2_bufchan_buf[0]))
        es_7_1_2MyFalse_2_bufchan_buf <= 1'd0;
      else if (((! es_7_1_2MyFalse_2_argbuf_r) && (! es_7_1_2MyFalse_2_bufchan_buf[0])))
        es_7_1_2MyFalse_2_bufchan_buf <= es_7_1_2MyFalse_2_bufchan_d;
  
  /* fork (Ty Go) : (es_7_1_2MyTrue,Go) > [(es_7_1_2MyTrue_1,Go),
                                      (es_7_1_2MyTrue_2,Go)] */
  logic [1:0] es_7_1_2MyTrue_emitted;
  logic [1:0] es_7_1_2MyTrue_done;
  assign es_7_1_2MyTrue_1_d = (es_7_1_2MyTrue_d[0] && (! es_7_1_2MyTrue_emitted[0]));
  assign es_7_1_2MyTrue_2_d = (es_7_1_2MyTrue_d[0] && (! es_7_1_2MyTrue_emitted[1]));
  assign es_7_1_2MyTrue_done = (es_7_1_2MyTrue_emitted | ({es_7_1_2MyTrue_2_d[0],
                                                           es_7_1_2MyTrue_1_d[0]} & {es_7_1_2MyTrue_2_r,
                                                                                     es_7_1_2MyTrue_1_r}));
  assign es_7_1_2MyTrue_r = (& es_7_1_2MyTrue_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyTrue_emitted <= 2'd0;
    else
      es_7_1_2MyTrue_emitted <= (es_7_1_2MyTrue_r ? 2'd0 :
                                 es_7_1_2MyTrue_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(es_7_1_2MyTrue_1,Go)] > (es_7_1_2MyTrue_1QNone_Int,QTree_Int) */
  assign es_7_1_2MyTrue_1QNone_Int_d = QNone_Int_dc((& {es_7_1_2MyTrue_1_d[0]}), es_7_1_2MyTrue_1_d);
  assign {es_7_1_2MyTrue_1_r} = {1 {(es_7_1_2MyTrue_1QNone_Int_r && es_7_1_2MyTrue_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (es_7_1_2MyTrue_1QNone_Int,QTree_Int) > (lizzieLet9_1_argbuf,QTree_Int) */
  QTree_Int_t es_7_1_2MyTrue_1QNone_Int_bufchan_d;
  logic es_7_1_2MyTrue_1QNone_Int_bufchan_r;
  assign es_7_1_2MyTrue_1QNone_Int_r = ((! es_7_1_2MyTrue_1QNone_Int_bufchan_d[0]) || es_7_1_2MyTrue_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_7_1_2MyTrue_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_7_1_2MyTrue_1QNone_Int_r)
        es_7_1_2MyTrue_1QNone_Int_bufchan_d <= es_7_1_2MyTrue_1QNone_Int_d;
  QTree_Int_t es_7_1_2MyTrue_1QNone_Int_bufchan_buf;
  assign es_7_1_2MyTrue_1QNone_Int_bufchan_r = (! es_7_1_2MyTrue_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet9_1_argbuf_d = (es_7_1_2MyTrue_1QNone_Int_bufchan_buf[0] ? es_7_1_2MyTrue_1QNone_Int_bufchan_buf :
                                  es_7_1_2MyTrue_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      es_7_1_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet9_1_argbuf_r && es_7_1_2MyTrue_1QNone_Int_bufchan_buf[0]))
        es_7_1_2MyTrue_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet9_1_argbuf_r) && (! es_7_1_2MyTrue_1QNone_Int_bufchan_buf[0])))
        es_7_1_2MyTrue_1QNone_Int_bufchan_buf <= es_7_1_2MyTrue_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (es_7_1_2MyTrue_2,Go) > (es_7_1_2MyTrue_2_argbuf,Go) */
  Go_t es_7_1_2MyTrue_2_bufchan_d;
  logic es_7_1_2MyTrue_2_bufchan_r;
  assign es_7_1_2MyTrue_2_r = ((! es_7_1_2MyTrue_2_bufchan_d[0]) || es_7_1_2MyTrue_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyTrue_2_bufchan_d <= 1'd0;
    else
      if (es_7_1_2MyTrue_2_r)
        es_7_1_2MyTrue_2_bufchan_d <= es_7_1_2MyTrue_2_d;
  Go_t es_7_1_2MyTrue_2_bufchan_buf;
  assign es_7_1_2MyTrue_2_bufchan_r = (! es_7_1_2MyTrue_2_bufchan_buf[0]);
  assign es_7_1_2MyTrue_2_argbuf_d = (es_7_1_2MyTrue_2_bufchan_buf[0] ? es_7_1_2MyTrue_2_bufchan_buf :
                                      es_7_1_2MyTrue_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_2MyTrue_2_bufchan_buf <= 1'd0;
    else
      if ((es_7_1_2MyTrue_2_argbuf_r && es_7_1_2MyTrue_2_bufchan_buf[0]))
        es_7_1_2MyTrue_2_bufchan_buf <= 1'd0;
      else if (((! es_7_1_2MyTrue_2_argbuf_r) && (! es_7_1_2MyTrue_2_bufchan_buf[0])))
        es_7_1_2MyTrue_2_bufchan_buf <= es_7_1_2MyTrue_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty MyDTInt_Int_Int) : (es_7_1_3,MyBool) (es_2_4MyFalse_2,MyDTInt_Int_Int) > [(es_7_1_3MyFalse,MyDTInt_Int_Int),
                                                                                    (_35,MyDTInt_Int_Int)] */
  logic [1:0] es_2_4MyFalse_2_onehotd;
  always_comb
    if ((es_7_1_3_d[0] && es_2_4MyFalse_2_d[0]))
      unique case (es_7_1_3_d[1:1])
        1'd0: es_2_4MyFalse_2_onehotd = 2'd1;
        1'd1: es_2_4MyFalse_2_onehotd = 2'd2;
        default: es_2_4MyFalse_2_onehotd = 2'd0;
      endcase
    else es_2_4MyFalse_2_onehotd = 2'd0;
  assign es_7_1_3MyFalse_d = es_2_4MyFalse_2_onehotd[0];
  assign _35_d = es_2_4MyFalse_2_onehotd[1];
  assign es_2_4MyFalse_2_r = (| (es_2_4MyFalse_2_onehotd & {_35_r,
                                                            es_7_1_3MyFalse_r}));
  assign es_7_1_3_r = es_2_4MyFalse_2_r;
  
  /* buf (Ty MyDTInt_Int_Int) : (es_7_1_3MyFalse,MyDTInt_Int_Int) > (es_7_1_3MyFalse_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t es_7_1_3MyFalse_bufchan_d;
  logic es_7_1_3MyFalse_bufchan_r;
  assign es_7_1_3MyFalse_r = ((! es_7_1_3MyFalse_bufchan_d[0]) || es_7_1_3MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_3MyFalse_bufchan_d <= 1'd0;
    else
      if (es_7_1_3MyFalse_r)
        es_7_1_3MyFalse_bufchan_d <= es_7_1_3MyFalse_d;
  MyDTInt_Int_Int_t es_7_1_3MyFalse_bufchan_buf;
  assign es_7_1_3MyFalse_bufchan_r = (! es_7_1_3MyFalse_bufchan_buf[0]);
  assign es_7_1_3MyFalse_1_argbuf_d = (es_7_1_3MyFalse_bufchan_buf[0] ? es_7_1_3MyFalse_bufchan_buf :
                                       es_7_1_3MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_3MyFalse_bufchan_buf <= 1'd0;
    else
      if ((es_7_1_3MyFalse_1_argbuf_r && es_7_1_3MyFalse_bufchan_buf[0]))
        es_7_1_3MyFalse_bufchan_buf <= 1'd0;
      else if (((! es_7_1_3MyFalse_1_argbuf_r) && (! es_7_1_3MyFalse_bufchan_buf[0])))
        es_7_1_3MyFalse_bufchan_buf <= es_7_1_3MyFalse_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(es_7_1_3MyFalse_1_argbuf,MyDTInt_Int_Int),
                                              (es_7_1_5MyFalse_1_argbuf,Int),
                                              (es_7_1_6MyFalse_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d = TupMyDTInt_Int_Int___Int___Int_dc((& {es_7_1_3MyFalse_1_argbuf_d[0],
                                                                                                       es_7_1_5MyFalse_1_argbuf_d[0],
                                                                                                       es_7_1_6MyFalse_1_argbuf_d[0]}), es_7_1_3MyFalse_1_argbuf_d, es_7_1_5MyFalse_1_argbuf_d, es_7_1_6MyFalse_1_argbuf_d);
  assign {es_7_1_3MyFalse_1_argbuf_r,
          es_7_1_5MyFalse_1_argbuf_r,
          es_7_1_6MyFalse_1_argbuf_r} = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int3_d[0])}};
  
  /* demux (Ty MyBool,
       Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (es_7_1_4,MyBool) (es_2_5MyFalse,Pointer_CTf'_f'_Int_Int_Int_Int) > [(es_7_1_4MyFalse,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                  (es_7_1_4MyTrue,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [1:0] es_2_5MyFalse_onehotd;
  always_comb
    if ((es_7_1_4_d[0] && es_2_5MyFalse_d[0]))
      unique case (es_7_1_4_d[1:1])
        1'd0: es_2_5MyFalse_onehotd = 2'd1;
        1'd1: es_2_5MyFalse_onehotd = 2'd2;
        default: es_2_5MyFalse_onehotd = 2'd0;
      endcase
    else es_2_5MyFalse_onehotd = 2'd0;
  assign es_7_1_4MyFalse_d = {es_2_5MyFalse_d[16:1],
                              es_2_5MyFalse_onehotd[0]};
  assign es_7_1_4MyTrue_d = {es_2_5MyFalse_d[16:1],
                             es_2_5MyFalse_onehotd[1]};
  assign es_2_5MyFalse_r = (| (es_2_5MyFalse_onehotd & {es_7_1_4MyTrue_r,
                                                        es_7_1_4MyFalse_r}));
  assign es_7_1_4_r = es_2_5MyFalse_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (es_7_1_4MyFalse,Pointer_CTf'_f'_Int_Int_Int_Int) > (es_7_1_4MyFalse_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyFalse_bufchan_d;
  logic es_7_1_4MyFalse_bufchan_r;
  assign es_7_1_4MyFalse_r = ((! es_7_1_4MyFalse_bufchan_d[0]) || es_7_1_4MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_4MyFalse_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_7_1_4MyFalse_r)
        es_7_1_4MyFalse_bufchan_d <= es_7_1_4MyFalse_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyFalse_bufchan_buf;
  assign es_7_1_4MyFalse_bufchan_r = (! es_7_1_4MyFalse_bufchan_buf[0]);
  assign es_7_1_4MyFalse_1_argbuf_d = (es_7_1_4MyFalse_bufchan_buf[0] ? es_7_1_4MyFalse_bufchan_buf :
                                       es_7_1_4MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_4MyFalse_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_7_1_4MyFalse_1_argbuf_r && es_7_1_4MyFalse_bufchan_buf[0]))
        es_7_1_4MyFalse_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_7_1_4MyFalse_1_argbuf_r) && (! es_7_1_4MyFalse_bufchan_buf[0])))
        es_7_1_4MyFalse_bufchan_buf <= es_7_1_4MyFalse_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (es_7_1_4MyTrue,Pointer_CTf'_f'_Int_Int_Int_Int) > (es_7_1_4MyTrue_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyTrue_bufchan_d;
  logic es_7_1_4MyTrue_bufchan_r;
  assign es_7_1_4MyTrue_r = ((! es_7_1_4MyTrue_bufchan_d[0]) || es_7_1_4MyTrue_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_4MyTrue_bufchan_d <= {16'd0, 1'd0};
    else
      if (es_7_1_4MyTrue_r) es_7_1_4MyTrue_bufchan_d <= es_7_1_4MyTrue_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  es_7_1_4MyTrue_bufchan_buf;
  assign es_7_1_4MyTrue_bufchan_r = (! es_7_1_4MyTrue_bufchan_buf[0]);
  assign es_7_1_4MyTrue_1_argbuf_d = (es_7_1_4MyTrue_bufchan_buf[0] ? es_7_1_4MyTrue_bufchan_buf :
                                      es_7_1_4MyTrue_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_4MyTrue_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_7_1_4MyTrue_1_argbuf_r && es_7_1_4MyTrue_bufchan_buf[0]))
        es_7_1_4MyTrue_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_7_1_4MyTrue_1_argbuf_r) && (! es_7_1_4MyTrue_bufchan_buf[0])))
        es_7_1_4MyTrue_bufchan_buf <= es_7_1_4MyTrue_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_7_1_5,MyBool) (es_2_6MyFalse_2,Int) > [(es_7_1_5MyFalse,Int),
                                                            (_34,Int)] */
  logic [1:0] es_2_6MyFalse_2_onehotd;
  always_comb
    if ((es_7_1_5_d[0] && es_2_6MyFalse_2_d[0]))
      unique case (es_7_1_5_d[1:1])
        1'd0: es_2_6MyFalse_2_onehotd = 2'd1;
        1'd1: es_2_6MyFalse_2_onehotd = 2'd2;
        default: es_2_6MyFalse_2_onehotd = 2'd0;
      endcase
    else es_2_6MyFalse_2_onehotd = 2'd0;
  assign es_7_1_5MyFalse_d = {es_2_6MyFalse_2_d[32:1],
                              es_2_6MyFalse_2_onehotd[0]};
  assign _34_d = {es_2_6MyFalse_2_d[32:1],
                  es_2_6MyFalse_2_onehotd[1]};
  assign es_2_6MyFalse_2_r = (| (es_2_6MyFalse_2_onehotd & {_34_r,
                                                            es_7_1_5MyFalse_r}));
  assign es_7_1_5_r = es_2_6MyFalse_2_r;
  
  /* buf (Ty Int) : (es_7_1_5MyFalse,Int) > (es_7_1_5MyFalse_1_argbuf,Int) */
  Int_t es_7_1_5MyFalse_bufchan_d;
  logic es_7_1_5MyFalse_bufchan_r;
  assign es_7_1_5MyFalse_r = ((! es_7_1_5MyFalse_bufchan_d[0]) || es_7_1_5MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_5MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_7_1_5MyFalse_r)
        es_7_1_5MyFalse_bufchan_d <= es_7_1_5MyFalse_d;
  Int_t es_7_1_5MyFalse_bufchan_buf;
  assign es_7_1_5MyFalse_bufchan_r = (! es_7_1_5MyFalse_bufchan_buf[0]);
  assign es_7_1_5MyFalse_1_argbuf_d = (es_7_1_5MyFalse_bufchan_buf[0] ? es_7_1_5MyFalse_bufchan_buf :
                                       es_7_1_5MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_7_1_5MyFalse_1_argbuf_r && es_7_1_5MyFalse_bufchan_buf[0]))
        es_7_1_5MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_7_1_5MyFalse_1_argbuf_r) && (! es_7_1_5MyFalse_bufchan_buf[0])))
        es_7_1_5MyFalse_bufchan_buf <= es_7_1_5MyFalse_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Int) : (es_7_1_6,MyBool) (es_2_7MyFalse_2,Int) > [(es_7_1_6MyFalse,Int),
                                                            (_33,Int)] */
  logic [1:0] es_2_7MyFalse_2_onehotd;
  always_comb
    if ((es_7_1_6_d[0] && es_2_7MyFalse_2_d[0]))
      unique case (es_7_1_6_d[1:1])
        1'd0: es_2_7MyFalse_2_onehotd = 2'd1;
        1'd1: es_2_7MyFalse_2_onehotd = 2'd2;
        default: es_2_7MyFalse_2_onehotd = 2'd0;
      endcase
    else es_2_7MyFalse_2_onehotd = 2'd0;
  assign es_7_1_6MyFalse_d = {es_2_7MyFalse_2_d[32:1],
                              es_2_7MyFalse_2_onehotd[0]};
  assign _33_d = {es_2_7MyFalse_2_d[32:1],
                  es_2_7MyFalse_2_onehotd[1]};
  assign es_2_7MyFalse_2_r = (| (es_2_7MyFalse_2_onehotd & {_33_r,
                                                            es_7_1_6MyFalse_r}));
  assign es_7_1_6_r = es_2_7MyFalse_2_r;
  
  /* buf (Ty Int) : (es_7_1_6MyFalse,Int) > (es_7_1_6MyFalse_1_argbuf,Int) */
  Int_t es_7_1_6MyFalse_bufchan_d;
  logic es_7_1_6MyFalse_bufchan_r;
  assign es_7_1_6MyFalse_r = ((! es_7_1_6MyFalse_bufchan_d[0]) || es_7_1_6MyFalse_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_6MyFalse_bufchan_d <= {32'd0, 1'd0};
    else
      if (es_7_1_6MyFalse_r)
        es_7_1_6MyFalse_bufchan_d <= es_7_1_6MyFalse_d;
  Int_t es_7_1_6MyFalse_bufchan_buf;
  assign es_7_1_6MyFalse_bufchan_r = (! es_7_1_6MyFalse_bufchan_buf[0]);
  assign es_7_1_6MyFalse_1_argbuf_d = (es_7_1_6MyFalse_bufchan_buf[0] ? es_7_1_6MyFalse_bufchan_buf :
                                       es_7_1_6MyFalse_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_7_1_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((es_7_1_6MyFalse_1_argbuf_r && es_7_1_6MyFalse_bufchan_buf[0]))
        es_7_1_6MyFalse_bufchan_buf <= {32'd0, 1'd0};
      else if (((! es_7_1_6MyFalse_1_argbuf_r) && (! es_7_1_6MyFalse_bufchan_buf[0])))
        es_7_1_6MyFalse_bufchan_buf <= es_7_1_6MyFalse_bufchan_d;
  
  /* buf (Ty QTree_Int) : (es_8_1QVal_Int,QTree_Int) > (lizzieLet8_1_argbuf,QTree_Int) */
  QTree_Int_t es_8_1QVal_Int_bufchan_d;
  logic es_8_1QVal_Int_bufchan_r;
  assign es_8_1QVal_Int_r = ((! es_8_1QVal_Int_bufchan_d[0]) || es_8_1QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_8_1QVal_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (es_8_1QVal_Int_r) es_8_1QVal_Int_bufchan_d <= es_8_1QVal_Int_d;
  QTree_Int_t es_8_1QVal_Int_bufchan_buf;
  assign es_8_1QVal_Int_bufchan_r = (! es_8_1QVal_Int_bufchan_buf[0]);
  assign lizzieLet8_1_argbuf_d = (es_8_1QVal_Int_bufchan_buf[0] ? es_8_1QVal_Int_bufchan_buf :
                                  es_8_1QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) es_8_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet8_1_argbuf_r && es_8_1QVal_Int_bufchan_buf[0]))
        es_8_1QVal_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet8_1_argbuf_r) && (! es_8_1QVal_Int_bufchan_buf[0])))
        es_8_1QVal_Int_bufchan_buf <= es_8_1QVal_Int_bufchan_d;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int,
          Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int) > [(f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13,Go),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1,Int),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                        (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1,MyDTInt_Int)] */
  logic [6:0] \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted ;
  logic [6:0] \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_done ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_d  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [0]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_d  = {\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [16:1],
                                                                                                                                          (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [1]))};
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_d  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [2]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_d  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [3]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_d  = {\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [48:17],
                                                                                                                                         (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [4]))};
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_d  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [5]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_d  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted [6]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_done  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted  | ({\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_d [0],
                                                                                                                                                                                                                                                                           \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0]} & {\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_r ,
                                                                                                                                                                                                                                                                                                                                                                                                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_r }));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_r  = (& \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted  <= 7'd0;
    else
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_emitted  <= (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_r  ? 7'd0 :
                                                                                                                                         \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_done );
  
  /* buf (Ty MyDTInt_Int) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1,MyDTInt_Int) > (f_mapaia_1_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_d ;
  MyDTInt_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf [0]);
  assign f_mapaia_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf  :
                                  \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf  <= 1'd0;
    else
      if ((f_mapaia_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf  <= 1'd0;
      else if (((! f_mapaia_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intf_mapaia_1_bufchan_d ;
  
  /* fork (Ty Go) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13,Go) > [(go_13_1,Go),
                                                                                                                                               (go_13_2,Go)] */
  logic [1:0] \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted ;
  logic [1:0] \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_done ;
  assign go_13_1_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted [0]));
  assign go_13_2_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_d [0] && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted [1]));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_done  = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  | ({go_13_2_d[0],
                                                                                                                                                                                                                                                                                 go_13_1_d[0]} & {go_13_2_r,
                                                                                                                                                                                                                                                                                                  go_13_1_r}));
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_r  = (& \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  <= 2'd0;
    else
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_emitted  <= (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_r  ? 2'd0 :
                                                                                                                                            \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intgo_13_done );
  
  /* buf (Ty MyDTInt_Bool) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1,MyDTInt_Bool) > (is_z_kronai6_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_d ;
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf [0]);
  assign is_z_kronai6_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf  :
                                      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf  <= 1'd0;
    else
      if ((is_z_kronai6_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf  <= 1'd0;
      else if (((! is_z_kronai6_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_kronai6_1_bufchan_d ;
  
  /* buf (Ty MyDTInt_Bool) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1,MyDTInt_Bool) > (is_z_mapai9_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_d ;
  MyDTInt_Bool_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf [0]);
  assign is_z_mapai9_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf  :
                                     \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf  <= 1'd0;
    else
      if ((is_z_mapai9_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf  <= 1'd0;
      else if (((! is_z_mapai9_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intis_z_mapai9_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1,Pointer_QTree_Int) > (m2ai5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d  <= {16'd0,
                                                                                                                                                1'd0};
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_d ;
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf [0]);
  assign m2ai5_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf  :
                               \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf  <= {16'd0,
                                                                                                                                                  1'd0};
    else
      if ((m2ai5_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf  <= {16'd0,
                                                                                                                                                    1'd0};
      else if (((! m2ai5_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intm2ai5_1_bufchan_d ;
  
  /* buf (Ty MyDTInt_Int_Int) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1,MyDTInt_Int_Int) > (op_kronai7_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d  <= 1'd0;
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_d ;
  MyDTInt_Int_Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf [0]);
  assign op_kronai7_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf  :
                                    \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf  <= 1'd0;
    else
      if ((op_kronai7_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf  <= 1'd0;
      else if (((! op_kronai7_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intop_kronai7_1_bufchan_d ;
  
  /* buf (Ty Int) : (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1,Int) > (vai8_1_1_argbuf,Int) */
  Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d ;
  logic \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_r ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_r  = ((! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d [0]) || \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d  <= {32'd0,
                                                                                                                                               1'd0};
    else
      if (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_r )
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_d ;
  Int_t \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_r  = (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf [0]);
  assign vai8_1_1_argbuf_d = (\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf [0] ? \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf  :
                              \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf  <= {32'd0,
                                                                                                                                                 1'd0};
    else
      if ((vai8_1_1_argbuf_r && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf  <= {32'd0,
                                                                                                                                                   1'd0};
      else if (((! vai8_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_buf  <= \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Intvai8_1_bufchan_d ;
  
  /* buf (Ty Pointer_QTree_Int) : (f'_f'_Int_Int_Int_Int_resbuf,Pointer_QTree_Int) > (lizzieLet8_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d ;
  logic \f'_f'_Int_Int_Int_Int_resbuf_bufchan_r ;
  assign \f'_f'_Int_Int_Int_Int_resbuf_r  = ((! \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d [0]) || \f'_f'_Int_Int_Int_Int_resbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d  <= {16'd0, 1'd0};
    else
      if (\f'_f'_Int_Int_Int_Int_resbuf_r )
        \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d  <= \f'_f'_Int_Int_Int_Int_resbuf_d ;
  Pointer_QTree_Int_t \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf ;
  assign \f'_f'_Int_Int_Int_Int_resbuf_bufchan_r  = (! \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf [0]);
  assign lizzieLet8_1_1_argbuf_d = (\f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf [0] ? \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf  :
                                    \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
    else
      if ((lizzieLet8_1_1_argbuf_r && \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf [0]))
        \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf  <= {16'd0, 1'd0};
      else if (((! lizzieLet8_1_1_argbuf_r) && (! \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf [0])))
        \f'_f'_Int_Int_Int_Int_resbuf_bufchan_buf  <= \f'_f'_Int_Int_Int_Int_resbuf_bufchan_d ;
  
  /* destruct (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int,
          Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int) > [(f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14,Go),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1,Pointer_QTree_Int),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1,MyDTInt_Int_Int),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1,MyDTInt_Bool),
                                                                                                                                                                                                                                                                                                                                                                                (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1,MyDTInt_Int)] */
  logic [6:0] f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted;
  logic [6:0] f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_done;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[0]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_d = {f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[16:1],
                                                                                                                                                    (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[1]))};
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_d = {f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[32:17],
                                                                                                                                                    (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[2]))};
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[3]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[4]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[5]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted[6]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_done = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted | ({f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_d[0],
                                                                                                                                                                                                                                                                                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_d[0]} & {f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_r,
                                                                                                                                                                                                                                                                                                                                                                                                                                            f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_r}));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_r = (& f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted <= 7'd0;
    else
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_emitted <= (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_r ? 7'd0 :
                                                                                                                                                   f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_done);
  
  /* buf (Ty MyDTInt_Int) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1,MyDTInt_Int) > (f_mapahZ_1_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_d;
  MyDTInt_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf[0]);
  assign f_mapahZ_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf :
                                  f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf <= 1'd0;
    else
      if ((f_mapahZ_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf <= 1'd0;
      else if (((! f_mapahZ_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intf_mapahZ_1_bufchan_d;
  
  /* fork (Ty Go) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14,Go) > [(go_14_1,Go),
                                                                                                                                                           (go_14_2,Go)] */
  logic [1:0] f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted;
  logic [1:0] f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_done;
  assign go_14_1_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted[0]));
  assign go_14_2_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_d[0] && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted[1]));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_done = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted | ({go_14_2_d[0],
                                                                                                                                                                                                                                                                                                     go_14_1_d[0]} & {go_14_2_r,
                                                                                                                                                                                                                                                                                                                      go_14_1_r}));
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_r = (& f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted <= 2'd0;
    else
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_emitted <= (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_r ? 2'd0 :
                                                                                                                                                      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intgo_14_done);
  
  /* buf (Ty MyDTInt_Bool) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1,MyDTInt_Bool) > (is_z_kronahW_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_d;
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf[0]);
  assign is_z_kronahW_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf :
                                      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronahW_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf <= 1'd0;
      else if (((! is_z_kronahW_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_kronahW_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1,MyDTInt_Bool) > (is_z_mapahY_1_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_d;
  MyDTInt_Bool_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf[0]);
  assign is_z_mapahY_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf :
                                     f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapahY_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf <= 1'd0;
      else if (((! is_z_mapahY_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intis_z_mapahY_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1,Pointer_QTree_Int) > (m1ahU_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d <= {16'd0,
                                                                                                                                                          1'd0};
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_d;
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf[0]);
  assign m1ahU_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf :
                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf <= {16'd0,
                                                                                                                                                            1'd0};
    else
      if ((m1ahU_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf <= {16'd0,
                                                                                                                                                              1'd0};
      else if (((! m1ahU_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm1ahU_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1,Pointer_QTree_Int) > (m2ahV_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d <= {16'd0,
                                                                                                                                                          1'd0};
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_d;
  Pointer_QTree_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf[0]);
  assign m2ahV_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf :
                               f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf <= {16'd0,
                                                                                                                                                            1'd0};
    else
      if ((m2ahV_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf <= {16'd0,
                                                                                                                                                              1'd0};
      else if (((! m2ahV_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intm2ahV_1_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1,MyDTInt_Int_Int) > (op_kronahX_1_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d;
  logic f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_r;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_r = ((! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d[0]) || f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d <= 1'd0;
    else
      if (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_r)
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_d;
  MyDTInt_Int_Int_t f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf;
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_r = (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf[0]);
  assign op_kronahX_1_1_argbuf_d = (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf[0] ? f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf :
                                    f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf <= 1'd0;
    else
      if ((op_kronahX_1_1_argbuf_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf[0]))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf <= 1'd0;
      else if (((! op_kronahX_1_1_argbuf_r) && (! f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf[0])))
        f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_buf <= f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Intop_kronahX_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (f_f_Int_Int_Int_Int_resbuf,Pointer_QTree_Int) > (es_0_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t f_f_Int_Int_Int_Int_resbuf_bufchan_d;
  logic f_f_Int_Int_Int_Int_resbuf_bufchan_r;
  assign f_f_Int_Int_Int_Int_resbuf_r = ((! f_f_Int_Int_Int_Int_resbuf_bufchan_d[0]) || f_f_Int_Int_Int_Int_resbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_Int_resbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (f_f_Int_Int_Int_Int_resbuf_r)
        f_f_Int_Int_Int_Int_resbuf_bufchan_d <= f_f_Int_Int_Int_Int_resbuf_d;
  Pointer_QTree_Int_t f_f_Int_Int_Int_Int_resbuf_bufchan_buf;
  assign f_f_Int_Int_Int_Int_resbuf_bufchan_r = (! f_f_Int_Int_Int_Int_resbuf_bufchan_buf[0]);
  assign es_0_1_argbuf_d = (f_f_Int_Int_Int_Int_resbuf_bufchan_buf[0] ? f_f_Int_Int_Int_Int_resbuf_bufchan_buf :
                            f_f_Int_Int_Int_Int_resbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      f_f_Int_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((es_0_1_argbuf_r && f_f_Int_Int_Int_Int_resbuf_bufchan_buf[0]))
        f_f_Int_Int_Int_Int_resbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! es_0_1_argbuf_r) && (! f_f_Int_Int_Int_Int_resbuf_bufchan_buf[0])))
        f_f_Int_Int_Int_Int_resbuf_bufchan_buf <= f_f_Int_Int_Int_Int_resbuf_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (f_mapahZ_2_2,MyDTInt_Int) > (f_mapahZ_2_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapahZ_2_2_bufchan_d;
  logic f_mapahZ_2_2_bufchan_r;
  assign f_mapahZ_2_2_r = ((! f_mapahZ_2_2_bufchan_d[0]) || f_mapahZ_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_2_2_bufchan_d <= 1'd0;
    else if (f_mapahZ_2_2_r) f_mapahZ_2_2_bufchan_d <= f_mapahZ_2_2_d;
  MyDTInt_Int_t f_mapahZ_2_2_bufchan_buf;
  assign f_mapahZ_2_2_bufchan_r = (! f_mapahZ_2_2_bufchan_buf[0]);
  assign f_mapahZ_2_2_argbuf_d = (f_mapahZ_2_2_bufchan_buf[0] ? f_mapahZ_2_2_bufchan_buf :
                                  f_mapahZ_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_2_2_bufchan_buf <= 1'd0;
    else
      if ((f_mapahZ_2_2_argbuf_r && f_mapahZ_2_2_bufchan_buf[0]))
        f_mapahZ_2_2_bufchan_buf <= 1'd0;
      else if (((! f_mapahZ_2_2_argbuf_r) && (! f_mapahZ_2_2_bufchan_buf[0])))
        f_mapahZ_2_2_bufchan_buf <= f_mapahZ_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (f_mapahZ_2_destruct,MyDTInt_Int) > [(f_mapahZ_2_1,MyDTInt_Int),
                                                             (f_mapahZ_2_2,MyDTInt_Int)] */
  logic [1:0] f_mapahZ_2_destruct_emitted;
  logic [1:0] f_mapahZ_2_destruct_done;
  assign f_mapahZ_2_1_d = (f_mapahZ_2_destruct_d[0] && (! f_mapahZ_2_destruct_emitted[0]));
  assign f_mapahZ_2_2_d = (f_mapahZ_2_destruct_d[0] && (! f_mapahZ_2_destruct_emitted[1]));
  assign f_mapahZ_2_destruct_done = (f_mapahZ_2_destruct_emitted | ({f_mapahZ_2_2_d[0],
                                                                     f_mapahZ_2_1_d[0]} & {f_mapahZ_2_2_r,
                                                                                           f_mapahZ_2_1_r}));
  assign f_mapahZ_2_destruct_r = (& f_mapahZ_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_2_destruct_emitted <= 2'd0;
    else
      f_mapahZ_2_destruct_emitted <= (f_mapahZ_2_destruct_r ? 2'd0 :
                                      f_mapahZ_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (f_mapahZ_3_2,MyDTInt_Int) > (f_mapahZ_3_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapahZ_3_2_bufchan_d;
  logic f_mapahZ_3_2_bufchan_r;
  assign f_mapahZ_3_2_r = ((! f_mapahZ_3_2_bufchan_d[0]) || f_mapahZ_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_3_2_bufchan_d <= 1'd0;
    else if (f_mapahZ_3_2_r) f_mapahZ_3_2_bufchan_d <= f_mapahZ_3_2_d;
  MyDTInt_Int_t f_mapahZ_3_2_bufchan_buf;
  assign f_mapahZ_3_2_bufchan_r = (! f_mapahZ_3_2_bufchan_buf[0]);
  assign f_mapahZ_3_2_argbuf_d = (f_mapahZ_3_2_bufchan_buf[0] ? f_mapahZ_3_2_bufchan_buf :
                                  f_mapahZ_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_3_2_bufchan_buf <= 1'd0;
    else
      if ((f_mapahZ_3_2_argbuf_r && f_mapahZ_3_2_bufchan_buf[0]))
        f_mapahZ_3_2_bufchan_buf <= 1'd0;
      else if (((! f_mapahZ_3_2_argbuf_r) && (! f_mapahZ_3_2_bufchan_buf[0])))
        f_mapahZ_3_2_bufchan_buf <= f_mapahZ_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (f_mapahZ_3_destruct,MyDTInt_Int) > [(f_mapahZ_3_1,MyDTInt_Int),
                                                             (f_mapahZ_3_2,MyDTInt_Int)] */
  logic [1:0] f_mapahZ_3_destruct_emitted;
  logic [1:0] f_mapahZ_3_destruct_done;
  assign f_mapahZ_3_1_d = (f_mapahZ_3_destruct_d[0] && (! f_mapahZ_3_destruct_emitted[0]));
  assign f_mapahZ_3_2_d = (f_mapahZ_3_destruct_d[0] && (! f_mapahZ_3_destruct_emitted[1]));
  assign f_mapahZ_3_destruct_done = (f_mapahZ_3_destruct_emitted | ({f_mapahZ_3_2_d[0],
                                                                     f_mapahZ_3_1_d[0]} & {f_mapahZ_3_2_r,
                                                                                           f_mapahZ_3_1_r}));
  assign f_mapahZ_3_destruct_r = (& f_mapahZ_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_3_destruct_emitted <= 2'd0;
    else
      f_mapahZ_3_destruct_emitted <= (f_mapahZ_3_destruct_r ? 2'd0 :
                                      f_mapahZ_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (f_mapahZ_4_destruct,MyDTInt_Int) > (f_mapahZ_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapahZ_4_destruct_bufchan_d;
  logic f_mapahZ_4_destruct_bufchan_r;
  assign f_mapahZ_4_destruct_r = ((! f_mapahZ_4_destruct_bufchan_d[0]) || f_mapahZ_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_4_destruct_bufchan_d <= 1'd0;
    else
      if (f_mapahZ_4_destruct_r)
        f_mapahZ_4_destruct_bufchan_d <= f_mapahZ_4_destruct_d;
  MyDTInt_Int_t f_mapahZ_4_destruct_bufchan_buf;
  assign f_mapahZ_4_destruct_bufchan_r = (! f_mapahZ_4_destruct_bufchan_buf[0]);
  assign f_mapahZ_4_1_argbuf_d = (f_mapahZ_4_destruct_bufchan_buf[0] ? f_mapahZ_4_destruct_bufchan_buf :
                                  f_mapahZ_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapahZ_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((f_mapahZ_4_1_argbuf_r && f_mapahZ_4_destruct_bufchan_buf[0]))
        f_mapahZ_4_destruct_bufchan_buf <= 1'd0;
      else if (((! f_mapahZ_4_1_argbuf_r) && (! f_mapahZ_4_destruct_bufchan_buf[0])))
        f_mapahZ_4_destruct_bufchan_buf <= f_mapahZ_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (f_mapaia_2_2,MyDTInt_Int) > (f_mapaia_2_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapaia_2_2_bufchan_d;
  logic f_mapaia_2_2_bufchan_r;
  assign f_mapaia_2_2_r = ((! f_mapaia_2_2_bufchan_d[0]) || f_mapaia_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_2_2_bufchan_d <= 1'd0;
    else if (f_mapaia_2_2_r) f_mapaia_2_2_bufchan_d <= f_mapaia_2_2_d;
  MyDTInt_Int_t f_mapaia_2_2_bufchan_buf;
  assign f_mapaia_2_2_bufchan_r = (! f_mapaia_2_2_bufchan_buf[0]);
  assign f_mapaia_2_2_argbuf_d = (f_mapaia_2_2_bufchan_buf[0] ? f_mapaia_2_2_bufchan_buf :
                                  f_mapaia_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_2_2_bufchan_buf <= 1'd0;
    else
      if ((f_mapaia_2_2_argbuf_r && f_mapaia_2_2_bufchan_buf[0]))
        f_mapaia_2_2_bufchan_buf <= 1'd0;
      else if (((! f_mapaia_2_2_argbuf_r) && (! f_mapaia_2_2_bufchan_buf[0])))
        f_mapaia_2_2_bufchan_buf <= f_mapaia_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (f_mapaia_2_destruct,MyDTInt_Int) > [(f_mapaia_2_1,MyDTInt_Int),
                                                             (f_mapaia_2_2,MyDTInt_Int)] */
  logic [1:0] f_mapaia_2_destruct_emitted;
  logic [1:0] f_mapaia_2_destruct_done;
  assign f_mapaia_2_1_d = (f_mapaia_2_destruct_d[0] && (! f_mapaia_2_destruct_emitted[0]));
  assign f_mapaia_2_2_d = (f_mapaia_2_destruct_d[0] && (! f_mapaia_2_destruct_emitted[1]));
  assign f_mapaia_2_destruct_done = (f_mapaia_2_destruct_emitted | ({f_mapaia_2_2_d[0],
                                                                     f_mapaia_2_1_d[0]} & {f_mapaia_2_2_r,
                                                                                           f_mapaia_2_1_r}));
  assign f_mapaia_2_destruct_r = (& f_mapaia_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_2_destruct_emitted <= 2'd0;
    else
      f_mapaia_2_destruct_emitted <= (f_mapaia_2_destruct_r ? 2'd0 :
                                      f_mapaia_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (f_mapaia_3_2,MyDTInt_Int) > (f_mapaia_3_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapaia_3_2_bufchan_d;
  logic f_mapaia_3_2_bufchan_r;
  assign f_mapaia_3_2_r = ((! f_mapaia_3_2_bufchan_d[0]) || f_mapaia_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_3_2_bufchan_d <= 1'd0;
    else if (f_mapaia_3_2_r) f_mapaia_3_2_bufchan_d <= f_mapaia_3_2_d;
  MyDTInt_Int_t f_mapaia_3_2_bufchan_buf;
  assign f_mapaia_3_2_bufchan_r = (! f_mapaia_3_2_bufchan_buf[0]);
  assign f_mapaia_3_2_argbuf_d = (f_mapaia_3_2_bufchan_buf[0] ? f_mapaia_3_2_bufchan_buf :
                                  f_mapaia_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_3_2_bufchan_buf <= 1'd0;
    else
      if ((f_mapaia_3_2_argbuf_r && f_mapaia_3_2_bufchan_buf[0]))
        f_mapaia_3_2_bufchan_buf <= 1'd0;
      else if (((! f_mapaia_3_2_argbuf_r) && (! f_mapaia_3_2_bufchan_buf[0])))
        f_mapaia_3_2_bufchan_buf <= f_mapaia_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int) : (f_mapaia_3_destruct,MyDTInt_Int) > [(f_mapaia_3_1,MyDTInt_Int),
                                                             (f_mapaia_3_2,MyDTInt_Int)] */
  logic [1:0] f_mapaia_3_destruct_emitted;
  logic [1:0] f_mapaia_3_destruct_done;
  assign f_mapaia_3_1_d = (f_mapaia_3_destruct_d[0] && (! f_mapaia_3_destruct_emitted[0]));
  assign f_mapaia_3_2_d = (f_mapaia_3_destruct_d[0] && (! f_mapaia_3_destruct_emitted[1]));
  assign f_mapaia_3_destruct_done = (f_mapaia_3_destruct_emitted | ({f_mapaia_3_2_d[0],
                                                                     f_mapaia_3_1_d[0]} & {f_mapaia_3_2_r,
                                                                                           f_mapaia_3_1_r}));
  assign f_mapaia_3_destruct_r = (& f_mapaia_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_3_destruct_emitted <= 2'd0;
    else
      f_mapaia_3_destruct_emitted <= (f_mapaia_3_destruct_r ? 2'd0 :
                                      f_mapaia_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int) : (f_mapaia_4_destruct,MyDTInt_Int) > (f_mapaia_4_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t f_mapaia_4_destruct_bufchan_d;
  logic f_mapaia_4_destruct_bufchan_r;
  assign f_mapaia_4_destruct_r = ((! f_mapaia_4_destruct_bufchan_d[0]) || f_mapaia_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_4_destruct_bufchan_d <= 1'd0;
    else
      if (f_mapaia_4_destruct_r)
        f_mapaia_4_destruct_bufchan_d <= f_mapaia_4_destruct_d;
  MyDTInt_Int_t f_mapaia_4_destruct_bufchan_buf;
  assign f_mapaia_4_destruct_bufchan_r = (! f_mapaia_4_destruct_bufchan_buf[0]);
  assign f_mapaia_4_1_argbuf_d = (f_mapaia_4_destruct_bufchan_buf[0] ? f_mapaia_4_destruct_bufchan_buf :
                                  f_mapaia_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) f_mapaia_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((f_mapaia_4_1_argbuf_r && f_mapaia_4_destruct_bufchan_buf[0]))
        f_mapaia_4_destruct_bufchan_buf <= 1'd0;
      else if (((! f_mapaia_4_1_argbuf_r) && (! f_mapaia_4_destruct_bufchan_buf[0])))
        f_mapaia_4_destruct_bufchan_buf <= f_mapaia_4_destruct_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int,
      Dcon Dcon_main1) : [(go_1,Go)] > (go_1Dcon_main1,MyDTInt_Int) */
  assign go_1Dcon_main1_d = Dcon_main1_dc((& {go_1_d[0]}), go_1_d);
  assign {go_1_r} = {1 {(go_1Dcon_main1_r && go_1Dcon_main1_d[0])}};
  
  /* fork (Ty C5) : (go_10_goMux_choice,C5) > [(go_10_goMux_choice_1,C5),
                                          (go_10_goMux_choice_2,C5)] */
  logic [1:0] go_10_goMux_choice_emitted;
  logic [1:0] go_10_goMux_choice_done;
  assign go_10_goMux_choice_1_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[0]))};
  assign go_10_goMux_choice_2_d = {go_10_goMux_choice_d[3:1],
                                   (go_10_goMux_choice_d[0] && (! go_10_goMux_choice_emitted[1]))};
  assign go_10_goMux_choice_done = (go_10_goMux_choice_emitted | ({go_10_goMux_choice_2_d[0],
                                                                   go_10_goMux_choice_1_d[0]} & {go_10_goMux_choice_2_r,
                                                                                                 go_10_goMux_choice_1_r}));
  assign go_10_goMux_choice_r = (& go_10_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_10_goMux_choice_emitted <= 2'd0;
    else
      go_10_goMux_choice_emitted <= (go_10_goMux_choice_r ? 2'd0 :
                                     go_10_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_10_goMux_choice_1,C5) [(call_$wnnz_Int_goMux2,Pointer_QTree_Int),
                                                        (q2abX_1_1_argbuf,Pointer_QTree_Int),
                                                        (q3abY_2_1_argbuf,Pointer_QTree_Int),
                                                        (q4abZ_3_1_argbuf,Pointer_QTree_Int),
                                                        (q1abW_1_argbuf,Pointer_QTree_Int)] > (wstH_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] wstH_1_goMux_mux_mux;
  logic [4:0] wstH_1_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_1_d[3:1])
      3'd0:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd1,
                                                           call_$wnnz_Int_goMux2_d};
      3'd1:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd2,
                                                           q2abX_1_1_argbuf_d};
      3'd2:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd4,
                                                           q3abY_2_1_argbuf_d};
      3'd3:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd8,
                                                           q4abZ_3_1_argbuf_d};
      3'd4:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd16,
                                                           q1abW_1_argbuf_d};
      default:
        {wstH_1_goMux_mux_onehot, wstH_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign wstH_1_goMux_mux_d = {wstH_1_goMux_mux_mux[16:1],
                               (wstH_1_goMux_mux_mux[0] && go_10_goMux_choice_1_d[0])};
  assign go_10_goMux_choice_1_r = (wstH_1_goMux_mux_d[0] && wstH_1_goMux_mux_r);
  assign {q1abW_1_argbuf_r,
          q4abZ_3_1_argbuf_r,
          q3abY_2_1_argbuf_r,
          q2abX_1_1_argbuf_r,
          call_$wnnz_Int_goMux2_r} = (go_10_goMux_choice_1_r ? wstH_1_goMux_mux_onehot :
                                      5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CT$wnnz_Int) : (go_10_goMux_choice_2,C5) [(call_$wnnz_Int_goMux3,Pointer_CT$wnnz_Int),
                                                          (sca2_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca1_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca0_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sca3_1_argbuf,Pointer_CT$wnnz_Int)] > (sc_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] sc_0_goMux_mux_mux;
  logic [4:0] sc_0_goMux_mux_onehot;
  always_comb
    unique case (go_10_goMux_choice_2_d[3:1])
      3'd0:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd1,
                                                       call_$wnnz_Int_goMux3_d};
      3'd1:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd2,
                                                       sca2_1_argbuf_d};
      3'd2:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd4,
                                                       sca1_1_argbuf_d};
      3'd3:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd8,
                                                       sca0_1_argbuf_d};
      3'd4:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd16,
                                                       sca3_1_argbuf_d};
      default:
        {sc_0_goMux_mux_onehot, sc_0_goMux_mux_mux} = {5'd0,
                                                       {16'd0, 1'd0}};
    endcase
  assign sc_0_goMux_mux_d = {sc_0_goMux_mux_mux[16:1],
                             (sc_0_goMux_mux_mux[0] && go_10_goMux_choice_2_d[0])};
  assign go_10_goMux_choice_2_r = (sc_0_goMux_mux_d[0] && sc_0_goMux_mux_r);
  assign {sca3_1_argbuf_r,
          sca0_1_argbuf_r,
          sca1_1_argbuf_r,
          sca2_1_argbuf_r,
          call_$wnnz_Int_goMux3_r} = (go_10_goMux_choice_2_r ? sc_0_goMux_mux_onehot :
                                      5'd0);
  
  /* fork (Ty C5) : (go_11_goMux_choice,C5) > [(go_11_goMux_choice_1,C5),
                                          (go_11_goMux_choice_2,C5),
                                          (go_11_goMux_choice_3,C5),
                                          (go_11_goMux_choice_4,C5),
                                          (go_11_goMux_choice_5,C5),
                                          (go_11_goMux_choice_6,C5),
                                          (go_11_goMux_choice_7,C5)] */
  logic [6:0] go_11_goMux_choice_emitted;
  logic [6:0] go_11_goMux_choice_done;
  assign go_11_goMux_choice_1_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[0]))};
  assign go_11_goMux_choice_2_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[1]))};
  assign go_11_goMux_choice_3_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[2]))};
  assign go_11_goMux_choice_4_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[3]))};
  assign go_11_goMux_choice_5_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[4]))};
  assign go_11_goMux_choice_6_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[5]))};
  assign go_11_goMux_choice_7_d = {go_11_goMux_choice_d[3:1],
                                   (go_11_goMux_choice_d[0] && (! go_11_goMux_choice_emitted[6]))};
  assign go_11_goMux_choice_done = (go_11_goMux_choice_emitted | ({go_11_goMux_choice_7_d[0],
                                                                   go_11_goMux_choice_6_d[0],
                                                                   go_11_goMux_choice_5_d[0],
                                                                   go_11_goMux_choice_4_d[0],
                                                                   go_11_goMux_choice_3_d[0],
                                                                   go_11_goMux_choice_2_d[0],
                                                                   go_11_goMux_choice_1_d[0]} & {go_11_goMux_choice_7_r,
                                                                                                 go_11_goMux_choice_6_r,
                                                                                                 go_11_goMux_choice_5_r,
                                                                                                 go_11_goMux_choice_4_r,
                                                                                                 go_11_goMux_choice_3_r,
                                                                                                 go_11_goMux_choice_2_r,
                                                                                                 go_11_goMux_choice_1_r}));
  assign go_11_goMux_choice_r = (& go_11_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_11_goMux_choice_emitted <= 7'd0;
    else
      go_11_goMux_choice_emitted <= (go_11_goMux_choice_r ? 7'd0 :
                                     go_11_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_11_goMux_choice_1,C5) [(call_f'_f'_Int_Int_Int_Int_goMux2,Pointer_QTree_Int),
                                                        (q3aie_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2aid_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1aic_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4aif_1_argbuf,Pointer_QTree_Int)] > (m2ai5_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2ai5_goMux_mux_mux;
  logic [4:0] m2ai5_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_1_d[3:1])
      3'd0:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd1,
                                                         \call_f'_f'_Int_Int_Int_Int_goMux2_d };
      3'd1:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd2,
                                                         q3aie_1_1_argbuf_d};
      3'd2:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd4,
                                                         q2aid_2_1_argbuf_d};
      3'd3:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd8,
                                                         q1aic_3_1_argbuf_d};
      3'd4:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd16,
                                                         q4aif_1_argbuf_d};
      default:
        {m2ai5_goMux_mux_onehot, m2ai5_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ai5_goMux_mux_d = {m2ai5_goMux_mux_mux[16:1],
                              (m2ai5_goMux_mux_mux[0] && go_11_goMux_choice_1_d[0])};
  assign go_11_goMux_choice_1_r = (m2ai5_goMux_mux_d[0] && m2ai5_goMux_mux_r);
  assign {q4aif_1_argbuf_r,
          q1aic_3_1_argbuf_r,
          q2aid_2_1_argbuf_r,
          q3aie_1_1_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux2_r } = (go_11_goMux_choice_1_r ? m2ai5_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_11_goMux_choice_2,C5) [(call_f'_f'_Int_Int_Int_Int_goMux3,MyDTInt_Bool),
                                                   (is_z_kronai6_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_kronai6_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_kronai6_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_kronai6_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_kronai6_goMux_mux_mux;
  logic [4:0] is_z_kronai6_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_2_d[3:1])
      3'd0:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd1,
                                        \call_f'_f'_Int_Int_Int_Int_goMux3_d };
      3'd1:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd2, is_z_kronai6_2_2_argbuf_d};
      3'd2:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd4, is_z_kronai6_3_2_argbuf_d};
      3'd3:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd8, is_z_kronai6_4_1_argbuf_d};
      3'd4:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd16,
                                        lizzieLet6_5QNode_Int_2_argbuf_d};
      default:
        {is_z_kronai6_goMux_mux_onehot,
         is_z_kronai6_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_z_kronai6_goMux_mux_d = (is_z_kronai6_goMux_mux_mux[0] && go_11_goMux_choice_2_d[0]);
  assign go_11_goMux_choice_2_r = (is_z_kronai6_goMux_mux_d[0] && is_z_kronai6_goMux_mux_r);
  assign {lizzieLet6_5QNode_Int_2_argbuf_r,
          is_z_kronai6_4_1_argbuf_r,
          is_z_kronai6_3_2_argbuf_r,
          is_z_kronai6_2_2_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux3_r } = (go_11_goMux_choice_2_r ? is_z_kronai6_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_11_goMux_choice_3,C5) [(call_f'_f'_Int_Int_Int_Int_goMux4,MyDTInt_Int_Int),
                                                      (op_kronai7_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_kronai7_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_kronai7_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet6_7QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_kronai7_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_kronai7_goMux_mux_mux;
  logic [4:0] op_kronai7_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_3_d[3:1])
      3'd0:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd1,
                                                                   \call_f'_f'_Int_Int_Int_Int_goMux4_d };
      3'd1:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd2,
                                                                   op_kronai7_2_2_argbuf_d};
      3'd2:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd4,
                                                                   op_kronai7_3_2_argbuf_d};
      3'd3:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd8,
                                                                   op_kronai7_4_1_argbuf_d};
      3'd4:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet6_7QNode_Int_2_argbuf_d};
      default:
        {op_kronai7_goMux_mux_onehot, op_kronai7_goMux_mux_mux} = {5'd0,
                                                                   1'd0};
    endcase
  assign op_kronai7_goMux_mux_d = (op_kronai7_goMux_mux_mux[0] && go_11_goMux_choice_3_d[0]);
  assign go_11_goMux_choice_3_r = (op_kronai7_goMux_mux_d[0] && op_kronai7_goMux_mux_r);
  assign {lizzieLet6_7QNode_Int_2_argbuf_r,
          op_kronai7_4_1_argbuf_r,
          op_kronai7_3_2_argbuf_r,
          op_kronai7_2_2_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux4_r } = (go_11_goMux_choice_3_r ? op_kronai7_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty Int) : (go_11_goMux_choice_4,C5) [(call_f'_f'_Int_Int_Int_Int_goMux5,Int),
                                          (vai8_2_2_argbuf,Int),
                                          (vai8_3_2_argbuf,Int),
                                          (vai8_4_1_argbuf,Int),
                                          (lizzieLet6_9QNode_Int_2_argbuf,Int)] > (vai8_goMux_mux,Int) */
  logic [32:0] vai8_goMux_mux_mux;
  logic [4:0] vai8_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_4_d[3:1])
      3'd0:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd1,
                                                       \call_f'_f'_Int_Int_Int_Int_goMux5_d };
      3'd1:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd2,
                                                       vai8_2_2_argbuf_d};
      3'd2:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd4,
                                                       vai8_3_2_argbuf_d};
      3'd3:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd8,
                                                       vai8_4_1_argbuf_d};
      3'd4:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd16,
                                                       lizzieLet6_9QNode_Int_2_argbuf_d};
      default:
        {vai8_goMux_mux_onehot, vai8_goMux_mux_mux} = {5'd0,
                                                       {32'd0, 1'd0}};
    endcase
  assign vai8_goMux_mux_d = {vai8_goMux_mux_mux[32:1],
                             (vai8_goMux_mux_mux[0] && go_11_goMux_choice_4_d[0])};
  assign go_11_goMux_choice_4_r = (vai8_goMux_mux_d[0] && vai8_goMux_mux_r);
  assign {lizzieLet6_9QNode_Int_2_argbuf_r,
          vai8_4_1_argbuf_r,
          vai8_3_2_argbuf_r,
          vai8_2_2_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux5_r } = (go_11_goMux_choice_4_r ? vai8_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_11_goMux_choice_5,C5) [(call_f'_f'_Int_Int_Int_Int_goMux6,MyDTInt_Bool),
                                                   (is_z_mapai9_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapai9_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapai9_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet6_6QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_mapai9_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_mapai9_goMux_mux_mux;
  logic [4:0] is_z_mapai9_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_5_d[3:1])
      3'd0:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd1,
                                                                     \call_f'_f'_Int_Int_Int_Int_goMux6_d };
      3'd1:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd2,
                                                                     is_z_mapai9_2_2_argbuf_d};
      3'd2:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd4,
                                                                     is_z_mapai9_3_2_argbuf_d};
      3'd3:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd8,
                                                                     is_z_mapai9_4_1_argbuf_d};
      3'd4:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd16,
                                                                     lizzieLet6_6QNode_Int_2_argbuf_d};
      default:
        {is_z_mapai9_goMux_mux_onehot, is_z_mapai9_goMux_mux_mux} = {5'd0,
                                                                     1'd0};
    endcase
  assign is_z_mapai9_goMux_mux_d = (is_z_mapai9_goMux_mux_mux[0] && go_11_goMux_choice_5_d[0]);
  assign go_11_goMux_choice_5_r = (is_z_mapai9_goMux_mux_d[0] && is_z_mapai9_goMux_mux_r);
  assign {lizzieLet6_6QNode_Int_2_argbuf_r,
          is_z_mapai9_4_1_argbuf_r,
          is_z_mapai9_3_2_argbuf_r,
          is_z_mapai9_2_2_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux6_r } = (go_11_goMux_choice_5_r ? is_z_mapai9_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int) : (go_11_goMux_choice_6,C5) [(call_f'_f'_Int_Int_Int_Int_goMux7,MyDTInt_Int),
                                                  (f_mapaia_2_2_argbuf,MyDTInt_Int),
                                                  (f_mapaia_3_2_argbuf,MyDTInt_Int),
                                                  (f_mapaia_4_1_argbuf,MyDTInt_Int),
                                                  (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int)] > (f_mapaia_goMux_mux,MyDTInt_Int) */
  logic [0:0] f_mapaia_goMux_mux_mux;
  logic [4:0] f_mapaia_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_6_d[3:1])
      3'd0:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd1,
                                                               \call_f'_f'_Int_Int_Int_Int_goMux7_d };
      3'd1:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd2,
                                                               f_mapaia_2_2_argbuf_d};
      3'd2:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd4,
                                                               f_mapaia_3_2_argbuf_d};
      3'd3:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd8,
                                                               f_mapaia_4_1_argbuf_d};
      3'd4:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd16,
                                                               lizzieLet6_3QNode_Int_2_argbuf_d};
      default:
        {f_mapaia_goMux_mux_onehot, f_mapaia_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign f_mapaia_goMux_mux_d = (f_mapaia_goMux_mux_mux[0] && go_11_goMux_choice_6_d[0]);
  assign go_11_goMux_choice_6_r = (f_mapaia_goMux_mux_d[0] && f_mapaia_goMux_mux_r);
  assign {lizzieLet6_3QNode_Int_2_argbuf_r,
          f_mapaia_4_1_argbuf_r,
          f_mapaia_3_2_argbuf_r,
          f_mapaia_2_2_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux7_r } = (go_11_goMux_choice_6_r ? f_mapaia_goMux_mux_onehot :
                                                    5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (go_11_goMux_choice_7,C5) [(call_f'_f'_Int_Int_Int_Int_goMux8,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (sca2_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (sca1_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (sca0_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (sca3_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int)] > (sc_0_1_goMux_mux,Pointer_CTf'_f'_Int_Int_Int_Int) */
  logic [16:0] sc_0_1_goMux_mux_mux;
  logic [4:0] sc_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_11_goMux_choice_7_d[3:1])
      3'd0:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd1,
                                                           \call_f'_f'_Int_Int_Int_Int_goMux8_d };
      3'd1:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd2,
                                                           sca2_1_1_argbuf_d};
      3'd2:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd4,
                                                           sca1_1_1_argbuf_d};
      3'd3:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd8,
                                                           sca0_1_1_argbuf_d};
      3'd4:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd16,
                                                           sca3_1_1_argbuf_d};
      default:
        {sc_0_1_goMux_mux_onehot, sc_0_1_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_1_goMux_mux_d = {sc_0_1_goMux_mux_mux[16:1],
                               (sc_0_1_goMux_mux_mux[0] && go_11_goMux_choice_7_d[0])};
  assign go_11_goMux_choice_7_r = (sc_0_1_goMux_mux_d[0] && sc_0_1_goMux_mux_r);
  assign {sca3_1_1_argbuf_r,
          sca0_1_1_argbuf_r,
          sca1_1_1_argbuf_r,
          sca2_1_1_argbuf_r,
          \call_f'_f'_Int_Int_Int_Int_goMux8_r } = (go_11_goMux_choice_7_r ? sc_0_1_goMux_mux_onehot :
                                                    5'd0);
  
  /* fork (Ty C5) : (go_12_goMux_choice,C5) > [(go_12_goMux_choice_1,C5),
                                          (go_12_goMux_choice_2,C5),
                                          (go_12_goMux_choice_3,C5),
                                          (go_12_goMux_choice_4,C5),
                                          (go_12_goMux_choice_5,C5),
                                          (go_12_goMux_choice_6,C5),
                                          (go_12_goMux_choice_7,C5)] */
  logic [6:0] go_12_goMux_choice_emitted;
  logic [6:0] go_12_goMux_choice_done;
  assign go_12_goMux_choice_1_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[0]))};
  assign go_12_goMux_choice_2_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[1]))};
  assign go_12_goMux_choice_3_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[2]))};
  assign go_12_goMux_choice_4_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[3]))};
  assign go_12_goMux_choice_5_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[4]))};
  assign go_12_goMux_choice_6_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[5]))};
  assign go_12_goMux_choice_7_d = {go_12_goMux_choice_d[3:1],
                                   (go_12_goMux_choice_d[0] && (! go_12_goMux_choice_emitted[6]))};
  assign go_12_goMux_choice_done = (go_12_goMux_choice_emitted | ({go_12_goMux_choice_7_d[0],
                                                                   go_12_goMux_choice_6_d[0],
                                                                   go_12_goMux_choice_5_d[0],
                                                                   go_12_goMux_choice_4_d[0],
                                                                   go_12_goMux_choice_3_d[0],
                                                                   go_12_goMux_choice_2_d[0],
                                                                   go_12_goMux_choice_1_d[0]} & {go_12_goMux_choice_7_r,
                                                                                                 go_12_goMux_choice_6_r,
                                                                                                 go_12_goMux_choice_5_r,
                                                                                                 go_12_goMux_choice_4_r,
                                                                                                 go_12_goMux_choice_3_r,
                                                                                                 go_12_goMux_choice_2_r,
                                                                                                 go_12_goMux_choice_1_r}));
  assign go_12_goMux_choice_r = (& go_12_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_12_goMux_choice_emitted <= 7'd0;
    else
      go_12_goMux_choice_emitted <= (go_12_goMux_choice_r ? 7'd0 :
                                     go_12_goMux_choice_done);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_1,C5) [(call_f_f_Int_Int_Int_Int_goMux2,Pointer_QTree_Int),
                                                        (q3ai3_1_1_argbuf,Pointer_QTree_Int),
                                                        (q2ai2_2_1_argbuf,Pointer_QTree_Int),
                                                        (q1ai1_3_1_argbuf,Pointer_QTree_Int),
                                                        (q4ai4_1_argbuf,Pointer_QTree_Int)] > (m1ahU_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m1ahU_goMux_mux_mux;
  logic [4:0] m1ahU_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_1_d[3:1])
      3'd0:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_Int_Int_Int_goMux2_d};
      3'd1:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd2,
                                                         q3ai3_1_1_argbuf_d};
      3'd2:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd4,
                                                         q2ai2_2_1_argbuf_d};
      3'd3:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd8,
                                                         q1ai1_3_1_argbuf_d};
      3'd4:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd16,
                                                         q4ai4_1_argbuf_d};
      default:
        {m1ahU_goMux_mux_onehot, m1ahU_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m1ahU_goMux_mux_d = {m1ahU_goMux_mux_mux[16:1],
                              (m1ahU_goMux_mux_mux[0] && go_12_goMux_choice_1_d[0])};
  assign go_12_goMux_choice_1_r = (m1ahU_goMux_mux_d[0] && m1ahU_goMux_mux_r);
  assign {q4ai4_1_argbuf_r,
          q1ai1_3_1_argbuf_r,
          q2ai2_2_1_argbuf_r,
          q3ai3_1_1_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux2_r} = (go_12_goMux_choice_1_r ? m1ahU_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_QTree_Int) : (go_12_goMux_choice_2,C5) [(call_f_f_Int_Int_Int_Int_goMux3,Pointer_QTree_Int),
                                                        (m2ahV_2_2_argbuf,Pointer_QTree_Int),
                                                        (m2ahV_3_2_argbuf,Pointer_QTree_Int),
                                                        (m2ahV_4_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet13_1_7QNode_Int_2_argbuf,Pointer_QTree_Int)] > (m2ahV_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] m2ahV_goMux_mux_mux;
  logic [4:0] m2ahV_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_2_d[3:1])
      3'd0:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd1,
                                                         call_f_f_Int_Int_Int_Int_goMux3_d};
      3'd1:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd2,
                                                         m2ahV_2_2_argbuf_d};
      3'd2:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd4,
                                                         m2ahV_3_2_argbuf_d};
      3'd3:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd8,
                                                         m2ahV_4_1_argbuf_d};
      3'd4:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd16,
                                                         lizzieLet13_1_7QNode_Int_2_argbuf_d};
      default:
        {m2ahV_goMux_mux_onehot, m2ahV_goMux_mux_mux} = {5'd0,
                                                         {16'd0, 1'd0}};
    endcase
  assign m2ahV_goMux_mux_d = {m2ahV_goMux_mux_mux[16:1],
                              (m2ahV_goMux_mux_mux[0] && go_12_goMux_choice_2_d[0])};
  assign go_12_goMux_choice_2_r = (m2ahV_goMux_mux_d[0] && m2ahV_goMux_mux_r);
  assign {lizzieLet13_1_7QNode_Int_2_argbuf_r,
          m2ahV_4_1_argbuf_r,
          m2ahV_3_2_argbuf_r,
          m2ahV_2_2_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux3_r} = (go_12_goMux_choice_2_r ? m2ahV_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_12_goMux_choice_3,C5) [(call_f_f_Int_Int_Int_Int_goMux4,MyDTInt_Bool),
                                                   (is_z_kronahW_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_kronahW_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_kronahW_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet13_1_5QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_kronahW_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_kronahW_goMux_mux_mux;
  logic [4:0] is_z_kronahW_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_3_d[3:1])
      3'd0:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd1,
                                        call_f_f_Int_Int_Int_Int_goMux4_d};
      3'd1:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd2, is_z_kronahW_2_2_argbuf_d};
      3'd2:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd4, is_z_kronahW_3_2_argbuf_d};
      3'd3:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd8, is_z_kronahW_4_1_argbuf_d};
      3'd4:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd16,
                                        lizzieLet13_1_5QNode_Int_2_argbuf_d};
      default:
        {is_z_kronahW_goMux_mux_onehot,
         is_z_kronahW_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign is_z_kronahW_goMux_mux_d = (is_z_kronahW_goMux_mux_mux[0] && go_12_goMux_choice_3_d[0]);
  assign go_12_goMux_choice_3_r = (is_z_kronahW_goMux_mux_d[0] && is_z_kronahW_goMux_mux_r);
  assign {lizzieLet13_1_5QNode_Int_2_argbuf_r,
          is_z_kronahW_4_1_argbuf_r,
          is_z_kronahW_3_2_argbuf_r,
          is_z_kronahW_2_2_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux4_r} = (go_12_goMux_choice_3_r ? is_z_kronahW_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int_Int) : (go_12_goMux_choice_4,C5) [(call_f_f_Int_Int_Int_Int_goMux5,MyDTInt_Int_Int),
                                                      (op_kronahX_2_2_argbuf,MyDTInt_Int_Int),
                                                      (op_kronahX_3_2_argbuf,MyDTInt_Int_Int),
                                                      (op_kronahX_4_1_argbuf,MyDTInt_Int_Int),
                                                      (lizzieLet13_1_8QNode_Int_2_argbuf,MyDTInt_Int_Int)] > (op_kronahX_goMux_mux,MyDTInt_Int_Int) */
  logic [0:0] op_kronahX_goMux_mux_mux;
  logic [4:0] op_kronahX_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_4_d[3:1])
      3'd0:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd1,
                                                                   call_f_f_Int_Int_Int_Int_goMux5_d};
      3'd1:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd2,
                                                                   op_kronahX_2_2_argbuf_d};
      3'd2:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd4,
                                                                   op_kronahX_3_2_argbuf_d};
      3'd3:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd8,
                                                                   op_kronahX_4_1_argbuf_d};
      3'd4:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd16,
                                                                   lizzieLet13_1_8QNode_Int_2_argbuf_d};
      default:
        {op_kronahX_goMux_mux_onehot, op_kronahX_goMux_mux_mux} = {5'd0,
                                                                   1'd0};
    endcase
  assign op_kronahX_goMux_mux_d = (op_kronahX_goMux_mux_mux[0] && go_12_goMux_choice_4_d[0]);
  assign go_12_goMux_choice_4_r = (op_kronahX_goMux_mux_d[0] && op_kronahX_goMux_mux_r);
  assign {lizzieLet13_1_8QNode_Int_2_argbuf_r,
          op_kronahX_4_1_argbuf_r,
          op_kronahX_3_2_argbuf_r,
          op_kronahX_2_2_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux5_r} = (go_12_goMux_choice_4_r ? op_kronahX_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Bool) : (go_12_goMux_choice_5,C5) [(call_f_f_Int_Int_Int_Int_goMux6,MyDTInt_Bool),
                                                   (is_z_mapahY_2_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapahY_3_2_argbuf,MyDTInt_Bool),
                                                   (is_z_mapahY_4_1_argbuf,MyDTInt_Bool),
                                                   (lizzieLet13_1_6QNode_Int_2_argbuf,MyDTInt_Bool)] > (is_z_mapahY_goMux_mux,MyDTInt_Bool) */
  logic [0:0] is_z_mapahY_goMux_mux_mux;
  logic [4:0] is_z_mapahY_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_5_d[3:1])
      3'd0:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd1,
                                                                     call_f_f_Int_Int_Int_Int_goMux6_d};
      3'd1:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd2,
                                                                     is_z_mapahY_2_2_argbuf_d};
      3'd2:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd4,
                                                                     is_z_mapahY_3_2_argbuf_d};
      3'd3:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd8,
                                                                     is_z_mapahY_4_1_argbuf_d};
      3'd4:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd16,
                                                                     lizzieLet13_1_6QNode_Int_2_argbuf_d};
      default:
        {is_z_mapahY_goMux_mux_onehot, is_z_mapahY_goMux_mux_mux} = {5'd0,
                                                                     1'd0};
    endcase
  assign is_z_mapahY_goMux_mux_d = (is_z_mapahY_goMux_mux_mux[0] && go_12_goMux_choice_5_d[0]);
  assign go_12_goMux_choice_5_r = (is_z_mapahY_goMux_mux_d[0] && is_z_mapahY_goMux_mux_r);
  assign {lizzieLet13_1_6QNode_Int_2_argbuf_r,
          is_z_mapahY_4_1_argbuf_r,
          is_z_mapahY_3_2_argbuf_r,
          is_z_mapahY_2_2_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux6_r} = (go_12_goMux_choice_5_r ? is_z_mapahY_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty MyDTInt_Int) : (go_12_goMux_choice_6,C5) [(call_f_f_Int_Int_Int_Int_goMux7,MyDTInt_Int),
                                                  (f_mapahZ_2_2_argbuf,MyDTInt_Int),
                                                  (f_mapahZ_3_2_argbuf,MyDTInt_Int),
                                                  (f_mapahZ_4_1_argbuf,MyDTInt_Int),
                                                  (lizzieLet13_1_3QNode_Int_2_argbuf,MyDTInt_Int)] > (f_mapahZ_goMux_mux,MyDTInt_Int) */
  logic [0:0] f_mapahZ_goMux_mux_mux;
  logic [4:0] f_mapahZ_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_6_d[3:1])
      3'd0:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd1,
                                                               call_f_f_Int_Int_Int_Int_goMux7_d};
      3'd1:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd2,
                                                               f_mapahZ_2_2_argbuf_d};
      3'd2:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd4,
                                                               f_mapahZ_3_2_argbuf_d};
      3'd3:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd8,
                                                               f_mapahZ_4_1_argbuf_d};
      3'd4:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd16,
                                                               lizzieLet13_1_3QNode_Int_2_argbuf_d};
      default:
        {f_mapahZ_goMux_mux_onehot, f_mapahZ_goMux_mux_mux} = {5'd0, 1'd0};
    endcase
  assign f_mapahZ_goMux_mux_d = (f_mapahZ_goMux_mux_mux[0] && go_12_goMux_choice_6_d[0]);
  assign go_12_goMux_choice_6_r = (f_mapahZ_goMux_mux_d[0] && f_mapahZ_goMux_mux_r);
  assign {lizzieLet13_1_3QNode_Int_2_argbuf_r,
          f_mapahZ_4_1_argbuf_r,
          f_mapahZ_3_2_argbuf_r,
          f_mapahZ_2_2_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux7_r} = (go_12_goMux_choice_6_r ? f_mapahZ_goMux_mux_onehot :
                                                5'd0);
  
  /* mux (Ty C5,
     Ty Pointer_CTf_f_Int_Int_Int_Int) : (go_12_goMux_choice_7,C5) [(call_f_f_Int_Int_Int_Int_goMux8,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (sca2_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (sca1_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (sca0_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (sca3_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int)] > (sc_0_2_goMux_mux,Pointer_CTf_f_Int_Int_Int_Int) */
  logic [16:0] sc_0_2_goMux_mux_mux;
  logic [4:0] sc_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_12_goMux_choice_7_d[3:1])
      3'd0:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd1,
                                                           call_f_f_Int_Int_Int_Int_goMux8_d};
      3'd1:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd2,
                                                           sca2_2_1_argbuf_d};
      3'd2:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd4,
                                                           sca1_2_1_argbuf_d};
      3'd3:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd8,
                                                           sca0_2_1_argbuf_d};
      3'd4:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd16,
                                                           sca3_2_1_argbuf_d};
      default:
        {sc_0_2_goMux_mux_onehot, sc_0_2_goMux_mux_mux} = {5'd0,
                                                           {16'd0, 1'd0}};
    endcase
  assign sc_0_2_goMux_mux_d = {sc_0_2_goMux_mux_mux[16:1],
                               (sc_0_2_goMux_mux_mux[0] && go_12_goMux_choice_7_d[0])};
  assign go_12_goMux_choice_7_r = (sc_0_2_goMux_mux_d[0] && sc_0_2_goMux_mux_r);
  assign {sca3_2_1_argbuf_r,
          sca0_2_1_argbuf_r,
          sca1_2_1_argbuf_r,
          sca2_2_1_argbuf_r,
          call_f_f_Int_Int_Int_Int_goMux8_r} = (go_12_goMux_choice_7_r ? sc_0_2_goMux_mux_onehot :
                                                5'd0);
  
  /* dcon (Ty CTf'_f'_Int_Int_Int_Int,
      Dcon Lf'_f'_Int_Int_Int_Intsbos) : [(go_13_1,Go)] > (go_13_1Lf'_f'_Int_Int_Int_Intsbos,CTf'_f'_Int_Int_Int_Int) */
  assign \go_13_1Lf'_f'_Int_Int_Int_Intsbos_d  = \Lf'_f'_Int_Int_Int_Intsbos_dc ((& {go_13_1_d[0]}), go_13_1_d);
  assign {go_13_1_r} = {1 {(\go_13_1Lf'_f'_Int_Int_Int_Intsbos_r  && \go_13_1Lf'_f'_Int_Int_Int_Intsbos_d [0])}};
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (go_13_1Lf'_f'_Int_Int_Int_Intsbos,CTf'_f'_Int_Int_Int_Int) > (lizzieLet17_1_argbuf,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d ;
  logic \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_r ;
  assign \go_13_1Lf'_f'_Int_Int_Int_Intsbos_r  = ((! \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d [0]) || \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d  <= {99'd0, 1'd0};
    else
      if (\go_13_1Lf'_f'_Int_Int_Int_Intsbos_r )
        \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d  <= \go_13_1Lf'_f'_Int_Int_Int_Intsbos_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf ;
  assign \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_r  = (! \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf [0]);
  assign lizzieLet17_1_argbuf_d = (\go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf [0] ? \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf  :
                                   \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
    else
      if ((lizzieLet17_1_argbuf_r && \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf [0]))
        \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf  <= {99'd0, 1'd0};
      else if (((! lizzieLet17_1_argbuf_r) && (! \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf [0])))
        \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_buf  <= \go_13_1Lf'_f'_Int_Int_Int_Intsbos_bufchan_d ;
  
  /* buf (Ty Go) : (go_13_2,Go) > (go_13_2_argbuf,Go) */
  Go_t go_13_2_bufchan_d;
  logic go_13_2_bufchan_r;
  assign go_13_2_r = ((! go_13_2_bufchan_d[0]) || go_13_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_d <= 1'd0;
    else if (go_13_2_r) go_13_2_bufchan_d <= go_13_2_d;
  Go_t go_13_2_bufchan_buf;
  assign go_13_2_bufchan_r = (! go_13_2_bufchan_buf[0]);
  assign go_13_2_argbuf_d = (go_13_2_bufchan_buf[0] ? go_13_2_bufchan_buf :
                             go_13_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_13_2_bufchan_buf <= 1'd0;
    else
      if ((go_13_2_argbuf_r && go_13_2_bufchan_buf[0]))
        go_13_2_bufchan_buf <= 1'd0;
      else if (((! go_13_2_argbuf_r) && (! go_13_2_bufchan_buf[0])))
        go_13_2_bufchan_buf <= go_13_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int) : [(go_13_2_argbuf,Go),
                                                                                                                                               (m2ai5_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                               (is_z_kronai6_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                               (op_kronai7_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                               (vai8_1_1_argbuf,Int),
                                                                                                                                               (is_z_mapai9_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                               (f_mapaia_1_1_argbuf,MyDTInt_Int),
                                                                                                                                               (lizzieLet6_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int)] > (call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int) */
  assign \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d  = \TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_dc ((& {go_13_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    m2ai5_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    is_z_kronai6_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    op_kronai7_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    vai8_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    is_z_mapai9_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    f_mapaia_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                    lizzieLet6_1_1_argbuf_d[0]}), go_13_2_argbuf_d, m2ai5_1_1_argbuf_d, is_z_kronai6_1_1_argbuf_d, op_kronai7_1_1_argbuf_d, vai8_1_1_argbuf_d, is_z_mapai9_1_1_argbuf_d, f_mapaia_1_1_argbuf_d, lizzieLet6_1_1_argbuf_d);
  assign {go_13_2_argbuf_r,
          m2ai5_1_1_argbuf_r,
          is_z_kronai6_1_1_argbuf_r,
          op_kronai7_1_1_argbuf_r,
          vai8_1_1_argbuf_r,
          is_z_mapai9_1_1_argbuf_r,
          f_mapaia_1_1_argbuf_r,
          lizzieLet6_1_1_argbuf_r} = {8 {(\call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_r  && \call_f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf'_f'_Int_Int_Int_Int_1_d [0])}};
  
  /* dcon (Ty CTf_f_Int_Int_Int_Int,
      Dcon Lf_f_Int_Int_Int_Intsbos) : [(go_14_1,Go)] > (go_14_1Lf_f_Int_Int_Int_Intsbos,CTf_f_Int_Int_Int_Int) */
  assign go_14_1Lf_f_Int_Int_Int_Intsbos_d = Lf_f_Int_Int_Int_Intsbos_dc((& {go_14_1_d[0]}), go_14_1_d);
  assign {go_14_1_r} = {1 {(go_14_1Lf_f_Int_Int_Int_Intsbos_r && go_14_1Lf_f_Int_Int_Int_Intsbos_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (go_14_1Lf_f_Int_Int_Int_Intsbos,CTf_f_Int_Int_Int_Int) > (lizzieLet18_1_argbuf,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d;
  logic go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_r;
  assign go_14_1Lf_f_Int_Int_Int_Intsbos_r = ((! go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d[0]) || go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d <= {83'd0, 1'd0};
    else
      if (go_14_1Lf_f_Int_Int_Int_Intsbos_r)
        go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d <= go_14_1Lf_f_Int_Int_Int_Intsbos_d;
  CTf_f_Int_Int_Int_Int_t go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf;
  assign go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_r = (! go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf[0]);
  assign lizzieLet18_1_argbuf_d = (go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf[0] ? go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf :
                                   go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
    else
      if ((lizzieLet18_1_argbuf_r && go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf[0]))
        go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf <= {83'd0, 1'd0};
      else if (((! lizzieLet18_1_argbuf_r) && (! go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf[0])))
        go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_buf <= go_14_1Lf_f_Int_Int_Int_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_14_2,Go) > (go_14_2_argbuf,Go) */
  Go_t go_14_2_bufchan_d;
  logic go_14_2_bufchan_r;
  assign go_14_2_r = ((! go_14_2_bufchan_d[0]) || go_14_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_d <= 1'd0;
    else if (go_14_2_r) go_14_2_bufchan_d <= go_14_2_d;
  Go_t go_14_2_bufchan_buf;
  assign go_14_2_bufchan_r = (! go_14_2_bufchan_buf[0]);
  assign go_14_2_argbuf_d = (go_14_2_bufchan_buf[0] ? go_14_2_bufchan_buf :
                             go_14_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_14_2_bufchan_buf <= 1'd0;
    else
      if ((go_14_2_argbuf_r && go_14_2_bufchan_buf[0]))
        go_14_2_bufchan_buf <= 1'd0;
      else if (((! go_14_2_argbuf_r) && (! go_14_2_bufchan_buf[0])))
        go_14_2_bufchan_buf <= go_14_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int) : [(go_14_2_argbuf,Go),
                                                                                                                                                           (m1ahU_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                                           (m2ahV_1_1_argbuf,Pointer_QTree_Int),
                                                                                                                                                           (is_z_kronahW_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                                           (op_kronahX_1_1_argbuf,MyDTInt_Int_Int),
                                                                                                                                                           (is_z_mapahY_1_1_argbuf,MyDTInt_Bool),
                                                                                                                                                           (f_mapahZ_1_1_argbuf,MyDTInt_Int),
                                                                                                                                                           (lizzieLet10_1_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int)] > (call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int) */
  assign call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_dc((& {go_14_2_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      m1ahU_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      m2ahV_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      is_z_kronahW_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      op_kronahX_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      is_z_mapahY_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      f_mapahZ_1_1_argbuf_d[0],
                                                                                                                                                                                                                                                                                                                                      lizzieLet10_1_1_argbuf_d[0]}), go_14_2_argbuf_d, m1ahU_1_1_argbuf_d, m2ahV_1_1_argbuf_d, is_z_kronahW_1_1_argbuf_d, op_kronahX_1_1_argbuf_d, is_z_mapahY_1_1_argbuf_d, f_mapahZ_1_1_argbuf_d, lizzieLet10_1_1_argbuf_d);
  assign {go_14_2_argbuf_r,
          m1ahU_1_1_argbuf_r,
          m2ahV_1_1_argbuf_r,
          is_z_kronahW_1_1_argbuf_r,
          op_kronahX_1_1_argbuf_r,
          is_z_mapahY_1_1_argbuf_r,
          f_mapahZ_1_1_argbuf_r,
          lizzieLet10_1_1_argbuf_r} = {8 {(call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_r && call_f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int___Pointer_CTf_f_Int_Int_Int_Int_1_d[0])}};
  
  /* fork (Ty C4) : (go_15_goMux_choice,C4) > [(go_15_goMux_choice_1,C4),
                                          (go_15_goMux_choice_2,C4)] */
  logic [1:0] go_15_goMux_choice_emitted;
  logic [1:0] go_15_goMux_choice_done;
  assign go_15_goMux_choice_1_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[0]))};
  assign go_15_goMux_choice_2_d = {go_15_goMux_choice_d[2:1],
                                   (go_15_goMux_choice_d[0] && (! go_15_goMux_choice_emitted[1]))};
  assign go_15_goMux_choice_done = (go_15_goMux_choice_emitted | ({go_15_goMux_choice_2_d[0],
                                                                   go_15_goMux_choice_1_d[0]} & {go_15_goMux_choice_2_r,
                                                                                                 go_15_goMux_choice_1_r}));
  assign go_15_goMux_choice_r = (& go_15_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_15_goMux_choice_emitted <= 2'd0;
    else
      go_15_goMux_choice_emitted <= (go_15_goMux_choice_r ? 2'd0 :
                                     go_15_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Int#) : (go_15_goMux_choice_1,C4) [(lizzieLet11_1_argbuf,Int#),
                                           (contRet_0_1_argbuf,Int#),
                                           (lizzieLet12_1_argbuf,Int#),
                                           (lizzieLet11_1_1_argbuf,Int#)] > (srtarg_0_goMux_mux,Int#) */
  logic [32:0] srtarg_0_goMux_mux_mux;
  logic [3:0] srtarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet11_1_argbuf_d};
      2'd1:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd2,
                                                               contRet_0_1_argbuf_d};
      2'd2:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet12_1_argbuf_d};
      2'd3:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet11_1_1_argbuf_d};
      default:
        {srtarg_0_goMux_mux_onehot, srtarg_0_goMux_mux_mux} = {4'd0,
                                                               {32'd0, 1'd0}};
    endcase
  assign srtarg_0_goMux_mux_d = {srtarg_0_goMux_mux_mux[32:1],
                                 (srtarg_0_goMux_mux_mux[0] && go_15_goMux_choice_1_d[0])};
  assign go_15_goMux_choice_1_r = (srtarg_0_goMux_mux_d[0] && srtarg_0_goMux_mux_r);
  assign {lizzieLet11_1_1_argbuf_r,
          lizzieLet12_1_argbuf_r,
          contRet_0_1_argbuf_r,
          lizzieLet11_1_argbuf_r} = (go_15_goMux_choice_1_r ? srtarg_0_goMux_mux_onehot :
                                     4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CT$wnnz_Int) : (go_15_goMux_choice_2,C4) [(lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (sc_0_6_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int),
                                                          (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int)] > (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) */
  logic [16:0] scfarg_0_goMux_mux_mux;
  logic [3:0] scfarg_0_goMux_mux_onehot;
  always_comb
    unique case (go_15_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd1,
                                                               lizzieLet4_4QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd2,
                                                               sc_0_6_1_argbuf_d};
      2'd2:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd4,
                                                               lizzieLet4_4QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd8,
                                                               lizzieLet4_4QError_Int_1_argbuf_d};
      default:
        {scfarg_0_goMux_mux_onehot, scfarg_0_goMux_mux_mux} = {4'd0,
                                                               {16'd0, 1'd0}};
    endcase
  assign scfarg_0_goMux_mux_d = {scfarg_0_goMux_mux_mux[16:1],
                                 (scfarg_0_goMux_mux_mux[0] && go_15_goMux_choice_2_d[0])};
  assign go_15_goMux_choice_2_r = (scfarg_0_goMux_mux_d[0] && scfarg_0_goMux_mux_r);
  assign {lizzieLet4_4QError_Int_1_argbuf_r,
          lizzieLet4_4QVal_Int_1_argbuf_r,
          sc_0_6_1_argbuf_r,
          lizzieLet4_4QNone_Int_1_argbuf_r} = (go_15_goMux_choice_2_r ? scfarg_0_goMux_mux_onehot :
                                               4'd0);
  
  /* fork (Ty C6) : (go_16_goMux_choice,C6) > [(go_16_goMux_choice_1,C6),
                                          (go_16_goMux_choice_2,C6)] */
  logic [1:0] go_16_goMux_choice_emitted;
  logic [1:0] go_16_goMux_choice_done;
  assign go_16_goMux_choice_1_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[0]))};
  assign go_16_goMux_choice_2_d = {go_16_goMux_choice_d[3:1],
                                   (go_16_goMux_choice_d[0] && (! go_16_goMux_choice_emitted[1]))};
  assign go_16_goMux_choice_done = (go_16_goMux_choice_emitted | ({go_16_goMux_choice_2_d[0],
                                                                   go_16_goMux_choice_1_d[0]} & {go_16_goMux_choice_2_r,
                                                                                                 go_16_goMux_choice_1_r}));
  assign go_16_goMux_choice_r = (& go_16_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_16_goMux_choice_emitted <= 2'd0;
    else
      go_16_goMux_choice_emitted <= (go_16_goMux_choice_r ? 2'd0 :
                                     go_16_goMux_choice_done);
  
  /* mux (Ty C6,
     Ty Pointer_QTree_Int) : (go_16_goMux_choice_1,C6) [(lizzieLet1_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet2_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet3_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet4_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet5_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_1_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_1_goMux_mux_mux;
  logic [5:0] srtarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_1_d[3:1])
      3'd0:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet1_1_1_argbuf_d};
      3'd1:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   contRet_0_1_1_argbuf_d};
      3'd2:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   lizzieLet2_1_1_argbuf_d};
      3'd3:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   lizzieLet3_1_1_argbuf_d};
      3'd4:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   lizzieLet4_1_1_argbuf_d};
      3'd5:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet5_1_1_argbuf_d};
      default:
        {srtarg_0_1_goMux_mux_onehot, srtarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_1_goMux_mux_d = {srtarg_0_1_goMux_mux_mux[16:1],
                                   (srtarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_1_d[0])};
  assign go_16_goMux_choice_1_r = (srtarg_0_1_goMux_mux_d[0] && srtarg_0_1_goMux_mux_r);
  assign {lizzieLet5_1_1_argbuf_r,
          lizzieLet4_1_1_argbuf_r,
          lizzieLet3_1_1_argbuf_r,
          lizzieLet2_1_1_argbuf_r,
          contRet_0_1_1_argbuf_r,
          lizzieLet1_1_1_argbuf_r} = (go_16_goMux_choice_1_r ? srtarg_0_1_goMux_mux_onehot :
                                      6'd0);
  
  /* mux (Ty C6,
     Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (go_16_goMux_choice_2,C6) [(lizzieLet6_8QNone_Int_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (sc_0_10_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (es_7_1_4MyFalse_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (es_7_1_4MyTrue_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (es_2_5MyTrue_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                      (lizzieLet6_8QError_Int_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int)] > (scfarg_0_1_goMux_mux,Pointer_CTf'_f'_Int_Int_Int_Int) */
  logic [16:0] scfarg_0_1_goMux_mux_mux;
  logic [5:0] scfarg_0_1_goMux_mux_onehot;
  always_comb
    unique case (go_16_goMux_choice_2_d[3:1])
      3'd0:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd1,
                                                                   lizzieLet6_8QNone_Int_1_argbuf_d};
      3'd1:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd2,
                                                                   sc_0_10_1_argbuf_d};
      3'd2:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd4,
                                                                   es_7_1_4MyFalse_1_argbuf_d};
      3'd3:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd8,
                                                                   es_7_1_4MyTrue_1_argbuf_d};
      3'd4:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd16,
                                                                   es_2_5MyTrue_1_argbuf_d};
      3'd5:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd32,
                                                                   lizzieLet6_8QError_Int_1_argbuf_d};
      default:
        {scfarg_0_1_goMux_mux_onehot, scfarg_0_1_goMux_mux_mux} = {6'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_1_goMux_mux_d = {scfarg_0_1_goMux_mux_mux[16:1],
                                   (scfarg_0_1_goMux_mux_mux[0] && go_16_goMux_choice_2_d[0])};
  assign go_16_goMux_choice_2_r = (scfarg_0_1_goMux_mux_d[0] && scfarg_0_1_goMux_mux_r);
  assign {lizzieLet6_8QError_Int_1_argbuf_r,
          es_2_5MyTrue_1_argbuf_r,
          es_7_1_4MyTrue_1_argbuf_r,
          es_7_1_4MyFalse_1_argbuf_r,
          sc_0_10_1_argbuf_r,
          lizzieLet6_8QNone_Int_1_argbuf_r} = (go_16_goMux_choice_2_r ? scfarg_0_1_goMux_mux_onehot :
                                               6'd0);
  
  /* fork (Ty C4) : (go_17_goMux_choice,C4) > [(go_17_goMux_choice_1,C4),
                                          (go_17_goMux_choice_2,C4)] */
  logic [1:0] go_17_goMux_choice_emitted;
  logic [1:0] go_17_goMux_choice_done;
  assign go_17_goMux_choice_1_d = {go_17_goMux_choice_d[2:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[0]))};
  assign go_17_goMux_choice_2_d = {go_17_goMux_choice_d[2:1],
                                   (go_17_goMux_choice_d[0] && (! go_17_goMux_choice_emitted[1]))};
  assign go_17_goMux_choice_done = (go_17_goMux_choice_emitted | ({go_17_goMux_choice_2_d[0],
                                                                   go_17_goMux_choice_1_d[0]} & {go_17_goMux_choice_2_r,
                                                                                                 go_17_goMux_choice_1_r}));
  assign go_17_goMux_choice_r = (& go_17_goMux_choice_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_17_goMux_choice_emitted <= 2'd0;
    else
      go_17_goMux_choice_emitted <= (go_17_goMux_choice_r ? 2'd0 :
                                     go_17_goMux_choice_done);
  
  /* mux (Ty C4,
     Ty Pointer_QTree_Int) : (go_17_goMux_choice_1,C4) [(lizzieLet7_1_1_argbuf,Pointer_QTree_Int),
                                                        (contRet_0_2_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet8_1_1_argbuf,Pointer_QTree_Int),
                                                        (lizzieLet9_1_1_argbuf,Pointer_QTree_Int)] > (srtarg_0_2_goMux_mux,Pointer_QTree_Int) */
  logic [16:0] srtarg_0_2_goMux_mux_mux;
  logic [3:0] srtarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_1_d[2:1])
      2'd0:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet7_1_1_argbuf_d};
      2'd1:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {4'd2,
                                                                   contRet_0_2_1_argbuf_d};
      2'd2:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet8_1_1_argbuf_d};
      2'd3:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet9_1_1_argbuf_d};
      default:
        {srtarg_0_2_goMux_mux_onehot, srtarg_0_2_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign srtarg_0_2_goMux_mux_d = {srtarg_0_2_goMux_mux_mux[16:1],
                                   (srtarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_1_d[0])};
  assign go_17_goMux_choice_1_r = (srtarg_0_2_goMux_mux_d[0] && srtarg_0_2_goMux_mux_r);
  assign {lizzieLet9_1_1_argbuf_r,
          lizzieLet8_1_1_argbuf_r,
          contRet_0_2_1_argbuf_r,
          lizzieLet7_1_1_argbuf_r} = (go_17_goMux_choice_1_r ? srtarg_0_2_goMux_mux_onehot :
                                      4'd0);
  
  /* mux (Ty C4,
     Ty Pointer_CTf_f_Int_Int_Int_Int) : (go_17_goMux_choice_2,C4) [(lizzieLet13_1_9QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (sc_0_14_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (lizzieLet13_1_9QVal_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int),
                                                                    (lizzieLet13_1_9QError_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int)] > (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int_Int_Int_Int) */
  logic [16:0] scfarg_0_2_goMux_mux_mux;
  logic [3:0] scfarg_0_2_goMux_mux_onehot;
  always_comb
    unique case (go_17_goMux_choice_2_d[2:1])
      2'd0:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {4'd1,
                                                                   lizzieLet13_1_9QNone_Int_1_argbuf_d};
      2'd1:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {4'd2,
                                                                   sc_0_14_1_argbuf_d};
      2'd2:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {4'd4,
                                                                   lizzieLet13_1_9QVal_Int_1_argbuf_d};
      2'd3:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {4'd8,
                                                                   lizzieLet13_1_9QError_Int_1_argbuf_d};
      default:
        {scfarg_0_2_goMux_mux_onehot, scfarg_0_2_goMux_mux_mux} = {4'd0,
                                                                   {16'd0, 1'd0}};
    endcase
  assign scfarg_0_2_goMux_mux_d = {scfarg_0_2_goMux_mux_mux[16:1],
                                   (scfarg_0_2_goMux_mux_mux[0] && go_17_goMux_choice_2_d[0])};
  assign go_17_goMux_choice_2_r = (scfarg_0_2_goMux_mux_d[0] && scfarg_0_2_goMux_mux_r);
  assign {lizzieLet13_1_9QError_Int_1_argbuf_r,
          lizzieLet13_1_9QVal_Int_1_argbuf_r,
          sc_0_14_1_argbuf_r,
          lizzieLet13_1_9QNone_Int_1_argbuf_r} = (go_17_goMux_choice_2_r ? scfarg_0_2_goMux_mux_onehot :
                                                  4'd0);
  
  /* buf (Ty MyDTInt_Int) : (go_1Dcon_main1,MyDTInt_Int) > (es_6_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t go_1Dcon_main1_bufchan_d;
  logic go_1Dcon_main1_bufchan_r;
  assign go_1Dcon_main1_r = ((! go_1Dcon_main1_bufchan_d[0]) || go_1Dcon_main1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1Dcon_main1_bufchan_d <= 1'd0;
    else
      if (go_1Dcon_main1_r) go_1Dcon_main1_bufchan_d <= go_1Dcon_main1_d;
  MyDTInt_Int_t go_1Dcon_main1_bufchan_buf;
  assign go_1Dcon_main1_bufchan_r = (! go_1Dcon_main1_bufchan_buf[0]);
  assign es_6_1_argbuf_d = (go_1Dcon_main1_bufchan_buf[0] ? go_1Dcon_main1_bufchan_buf :
                            go_1Dcon_main1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_1Dcon_main1_bufchan_buf <= 1'd0;
    else
      if ((es_6_1_argbuf_r && go_1Dcon_main1_bufchan_buf[0]))
        go_1Dcon_main1_bufchan_buf <= 1'd0;
      else if (((! es_6_1_argbuf_r) && (! go_1Dcon_main1_bufchan_buf[0])))
        go_1Dcon_main1_bufchan_buf <= go_1Dcon_main1_bufchan_d;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_eqZero) : [(go_2,Go)] > (go_2Dcon_eqZero,MyDTInt_Bool) */
  assign go_2Dcon_eqZero_d = Dcon_eqZero_dc((& {go_2_d[0]}), go_2_d);
  assign {go_2_r} = {1 {(go_2Dcon_eqZero_r && go_2Dcon_eqZero_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_2Dcon_eqZero,MyDTInt_Bool) > (es_5_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_2Dcon_eqZero_bufchan_d;
  logic go_2Dcon_eqZero_bufchan_r;
  assign go_2Dcon_eqZero_r = ((! go_2Dcon_eqZero_bufchan_d[0]) || go_2Dcon_eqZero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_eqZero_bufchan_d <= 1'd0;
    else
      if (go_2Dcon_eqZero_r)
        go_2Dcon_eqZero_bufchan_d <= go_2Dcon_eqZero_d;
  MyDTInt_Bool_t go_2Dcon_eqZero_bufchan_buf;
  assign go_2Dcon_eqZero_bufchan_r = (! go_2Dcon_eqZero_bufchan_buf[0]);
  assign es_5_1_argbuf_d = (go_2Dcon_eqZero_bufchan_buf[0] ? go_2Dcon_eqZero_bufchan_buf :
                            go_2Dcon_eqZero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_2Dcon_eqZero_bufchan_buf <= 1'd0;
    else
      if ((es_5_1_argbuf_r && go_2Dcon_eqZero_bufchan_buf[0]))
        go_2Dcon_eqZero_bufchan_buf <= 1'd0;
      else if (((! es_5_1_argbuf_r) && (! go_2Dcon_eqZero_bufchan_buf[0])))
        go_2Dcon_eqZero_bufchan_buf <= go_2Dcon_eqZero_bufchan_d;
  
  /* dcon (Ty MyDTInt_Int_Int,
      Dcon Dcon_$fNumInt_$c*) : [(go_3,Go)] > (go_3Dcon_$fNumInt_$c*,MyDTInt_Int_Int) */
  assign \go_3Dcon_$fNumInt_$ctimes_d  = \Dcon_$fNumInt_$ctimes_dc ((& {go_3_d[0]}), go_3_d);
  assign {go_3_r} = {1 {(\go_3Dcon_$fNumInt_$ctimes_r  && \go_3Dcon_$fNumInt_$ctimes_d [0])}};
  
  /* buf (Ty MyDTInt_Int_Int) : (go_3Dcon_$fNumInt_$c*,MyDTInt_Int_Int) > (es_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t \go_3Dcon_$fNumInt_$ctimes_bufchan_d ;
  logic \go_3Dcon_$fNumInt_$ctimes_bufchan_r ;
  assign \go_3Dcon_$fNumInt_$ctimes_r  = ((! \go_3Dcon_$fNumInt_$ctimes_bufchan_d [0]) || \go_3Dcon_$fNumInt_$ctimes_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \go_3Dcon_$fNumInt_$ctimes_bufchan_d  <= 1'd0;
    else
      if (\go_3Dcon_$fNumInt_$ctimes_r )
        \go_3Dcon_$fNumInt_$ctimes_bufchan_d  <= \go_3Dcon_$fNumInt_$ctimes_d ;
  MyDTInt_Int_Int_t \go_3Dcon_$fNumInt_$ctimes_bufchan_buf ;
  assign \go_3Dcon_$fNumInt_$ctimes_bufchan_r  = (! \go_3Dcon_$fNumInt_$ctimes_bufchan_buf [0]);
  assign es_4_1_argbuf_d = (\go_3Dcon_$fNumInt_$ctimes_bufchan_buf [0] ? \go_3Dcon_$fNumInt_$ctimes_bufchan_buf  :
                            \go_3Dcon_$fNumInt_$ctimes_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \go_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
    else
      if ((es_4_1_argbuf_r && \go_3Dcon_$fNumInt_$ctimes_bufchan_buf [0]))
        \go_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= 1'd0;
      else if (((! es_4_1_argbuf_r) && (! \go_3Dcon_$fNumInt_$ctimes_bufchan_buf [0])))
        \go_3Dcon_$fNumInt_$ctimes_bufchan_buf  <= \go_3Dcon_$fNumInt_$ctimes_bufchan_d ;
  
  /* dcon (Ty MyDTInt_Bool,
      Dcon Dcon_eqZero) : [(go_4,Go)] > (go_4Dcon_eqZero,MyDTInt_Bool) */
  assign go_4Dcon_eqZero_d = Dcon_eqZero_dc((& {go_4_d[0]}), go_4_d);
  assign {go_4_r} = {1 {(go_4Dcon_eqZero_r && go_4Dcon_eqZero_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (go_4Dcon_eqZero,MyDTInt_Bool) > (es_3_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t go_4Dcon_eqZero_bufchan_d;
  logic go_4Dcon_eqZero_bufchan_r;
  assign go_4Dcon_eqZero_r = ((! go_4Dcon_eqZero_bufchan_d[0]) || go_4Dcon_eqZero_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_eqZero_bufchan_d <= 1'd0;
    else
      if (go_4Dcon_eqZero_r)
        go_4Dcon_eqZero_bufchan_d <= go_4Dcon_eqZero_d;
  MyDTInt_Bool_t go_4Dcon_eqZero_bufchan_buf;
  assign go_4Dcon_eqZero_bufchan_r = (! go_4Dcon_eqZero_bufchan_buf[0]);
  assign es_3_1_argbuf_d = (go_4Dcon_eqZero_bufchan_buf[0] ? go_4Dcon_eqZero_bufchan_buf :
                            go_4Dcon_eqZero_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_4Dcon_eqZero_bufchan_buf <= 1'd0;
    else
      if ((es_3_1_argbuf_r && go_4Dcon_eqZero_bufchan_buf[0]))
        go_4Dcon_eqZero_bufchan_buf <= 1'd0;
      else if (((! es_3_1_argbuf_r) && (! go_4Dcon_eqZero_bufchan_buf[0])))
        go_4Dcon_eqZero_bufchan_buf <= go_4Dcon_eqZero_bufchan_d;
  
  /* buf (Ty Go) : (go_5,Go) > (go_5_argbuf,Go) */
  Go_t go_5_bufchan_d;
  logic go_5_bufchan_r;
  assign go_5_r = ((! go_5_bufchan_d[0]) || go_5_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_d <= 1'd0;
    else if (go_5_r) go_5_bufchan_d <= go_5_d;
  Go_t go_5_bufchan_buf;
  assign go_5_bufchan_r = (! go_5_bufchan_buf[0]);
  assign go_5_argbuf_d = (go_5_bufchan_buf[0] ? go_5_bufchan_buf :
                          go_5_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_5_bufchan_buf <= 1'd0;
    else
      if ((go_5_argbuf_r && go_5_bufchan_buf[0]))
        go_5_bufchan_buf <= 1'd0;
      else if (((! go_5_argbuf_r) && (! go_5_bufchan_buf[0])))
        go_5_bufchan_buf <= go_5_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int) : [(go_5_argbuf,Go),
                                                                                                                           (m1ahS_0,Pointer_QTree_Int),
                                                                                                                           (m2ahT_1,Pointer_QTree_Int),
                                                                                                                           (es_3_1_argbuf,MyDTInt_Bool),
                                                                                                                           (es_4_1_argbuf,MyDTInt_Int_Int),
                                                                                                                           (es_5_1_argbuf,MyDTInt_Bool),
                                                                                                                           (es_6_1_argbuf,MyDTInt_Int)] > (f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int) */
  assign f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_dc((& {go_5_argbuf_d[0],
                                                                                                                                                                                                                                                                 m1ahS_0_d[0],
                                                                                                                                                                                                                                                                 m2ahT_1_d[0],
                                                                                                                                                                                                                                                                 es_3_1_argbuf_d[0],
                                                                                                                                                                                                                                                                 es_4_1_argbuf_d[0],
                                                                                                                                                                                                                                                                 es_5_1_argbuf_d[0],
                                                                                                                                                                                                                                                                 es_6_1_argbuf_d[0]}), go_5_argbuf_d, m1ahS_0_d, m2ahT_1_d, es_3_1_argbuf_d, es_4_1_argbuf_d, es_5_1_argbuf_d, es_6_1_argbuf_d);
  assign {go_5_argbuf_r,
          m1ahS_0_r,
          m2ahT_1_r,
          es_3_1_argbuf_r,
          es_4_1_argbuf_r,
          es_5_1_argbuf_r,
          es_6_1_argbuf_r} = {7 {(f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_r && f_f_Int_Int_Int_IntTupGo___Pointer_QTree_Int___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___MyDTInt_Bool___MyDTInt_Int_1_d[0])}};
  
  /* buf (Ty Go) : (go_6,Go) > (go_6_argbuf,Go) */
  Go_t go_6_bufchan_d;
  logic go_6_bufchan_r;
  assign go_6_r = ((! go_6_bufchan_d[0]) || go_6_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_d <= 1'd0;
    else if (go_6_r) go_6_bufchan_d <= go_6_d;
  Go_t go_6_bufchan_buf;
  assign go_6_bufchan_r = (! go_6_bufchan_buf[0]);
  assign go_6_argbuf_d = (go_6_bufchan_buf[0] ? go_6_bufchan_buf :
                          go_6_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_6_bufchan_buf <= 1'd0;
    else
      if ((go_6_argbuf_r && go_6_bufchan_buf[0]))
        go_6_bufchan_buf <= 1'd0;
      else if (((! go_6_argbuf_r) && (! go_6_bufchan_buf[0])))
        go_6_bufchan_buf <= go_6_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int,
      Dcon TupGo___Pointer_QTree_Int) : [(go_6_argbuf,Go),
                                         (es_0_1_argbuf,Pointer_QTree_Int)] > ($wnnz_IntTupGo___Pointer_QTree_Int_1,TupGo___Pointer_QTree_Int) */
  assign \$wnnz_IntTupGo___Pointer_QTree_Int_1_d  = TupGo___Pointer_QTree_Int_dc((& {go_6_argbuf_d[0],
                                                                                     es_0_1_argbuf_d[0]}), go_6_argbuf_d, es_0_1_argbuf_d);
  assign {go_6_argbuf_r,
          es_0_1_argbuf_r} = {2 {(\$wnnz_IntTupGo___Pointer_QTree_Int_1_r  && \$wnnz_IntTupGo___Pointer_QTree_Int_1_d [0])}};
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon L$wnnz_Intsbos) : [(go_7_1,Go)] > (go_7_1L$wnnz_Intsbos,CT$wnnz_Int) */
  assign go_7_1L$wnnz_Intsbos_d = L$wnnz_Intsbos_dc((& {go_7_1_d[0]}), go_7_1_d);
  assign {go_7_1_r} = {1 {(go_7_1L$wnnz_Intsbos_r && go_7_1L$wnnz_Intsbos_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (go_7_1L$wnnz_Intsbos,CT$wnnz_Int) > (lizzieLet0_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t go_7_1L$wnnz_Intsbos_bufchan_d;
  logic go_7_1L$wnnz_Intsbos_bufchan_r;
  assign go_7_1L$wnnz_Intsbos_r = ((! go_7_1L$wnnz_Intsbos_bufchan_d[0]) || go_7_1L$wnnz_Intsbos_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_7_1L$wnnz_Intsbos_bufchan_d <= {115'd0, 1'd0};
    else
      if (go_7_1L$wnnz_Intsbos_r)
        go_7_1L$wnnz_Intsbos_bufchan_d <= go_7_1L$wnnz_Intsbos_d;
  CT$wnnz_Int_t go_7_1L$wnnz_Intsbos_bufchan_buf;
  assign go_7_1L$wnnz_Intsbos_bufchan_r = (! go_7_1L$wnnz_Intsbos_bufchan_buf[0]);
  assign lizzieLet0_1_argbuf_d = (go_7_1L$wnnz_Intsbos_bufchan_buf[0] ? go_7_1L$wnnz_Intsbos_bufchan_buf :
                                  go_7_1L$wnnz_Intsbos_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      go_7_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
    else
      if ((lizzieLet0_1_argbuf_r && go_7_1L$wnnz_Intsbos_bufchan_buf[0]))
        go_7_1L$wnnz_Intsbos_bufchan_buf <= {115'd0, 1'd0};
      else if (((! lizzieLet0_1_argbuf_r) && (! go_7_1L$wnnz_Intsbos_bufchan_buf[0])))
        go_7_1L$wnnz_Intsbos_bufchan_buf <= go_7_1L$wnnz_Intsbos_bufchan_d;
  
  /* buf (Ty Go) : (go_7_2,Go) > (go_7_2_argbuf,Go) */
  Go_t go_7_2_bufchan_d;
  logic go_7_2_bufchan_r;
  assign go_7_2_r = ((! go_7_2_bufchan_d[0]) || go_7_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_d <= 1'd0;
    else if (go_7_2_r) go_7_2_bufchan_d <= go_7_2_d;
  Go_t go_7_2_bufchan_buf;
  assign go_7_2_bufchan_r = (! go_7_2_bufchan_buf[0]);
  assign go_7_2_argbuf_d = (go_7_2_bufchan_buf[0] ? go_7_2_bufchan_buf :
                            go_7_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) go_7_2_bufchan_buf <= 1'd0;
    else
      if ((go_7_2_argbuf_r && go_7_2_bufchan_buf[0]))
        go_7_2_bufchan_buf <= 1'd0;
      else if (((! go_7_2_argbuf_r) && (! go_7_2_bufchan_buf[0])))
        go_7_2_bufchan_buf <= go_7_2_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int,
      Dcon TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) : [(go_7_2_argbuf,Go),
                                                               (wstH_1_argbuf,Pointer_QTree_Int),
                                                               (lizzieLet13_1_argbuf,Pointer_CT$wnnz_Int)] > (call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1,TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int) */
  assign call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d = TupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_dc((& {go_7_2_argbuf_d[0],
                                                                                                                                    wstH_1_argbuf_d[0],
                                                                                                                                    lizzieLet13_1_argbuf_d[0]}), go_7_2_argbuf_d, wstH_1_argbuf_d, lizzieLet13_1_argbuf_d);
  assign {go_7_2_argbuf_r,
          wstH_1_argbuf_r,
          lizzieLet13_1_argbuf_r} = {3 {(call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_r && call_$wnnz_IntTupGo___Pointer_QTree_Int___Pointer_CT$wnnz_Int_1_d[0])}};
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronahW_2_2,MyDTInt_Bool) > (is_z_kronahW_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronahW_2_2_bufchan_d;
  logic is_z_kronahW_2_2_bufchan_r;
  assign is_z_kronahW_2_2_r = ((! is_z_kronahW_2_2_bufchan_d[0]) || is_z_kronahW_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_kronahW_2_2_r)
        is_z_kronahW_2_2_bufchan_d <= is_z_kronahW_2_2_d;
  MyDTInt_Bool_t is_z_kronahW_2_2_bufchan_buf;
  assign is_z_kronahW_2_2_bufchan_r = (! is_z_kronahW_2_2_bufchan_buf[0]);
  assign is_z_kronahW_2_2_argbuf_d = (is_z_kronahW_2_2_bufchan_buf[0] ? is_z_kronahW_2_2_bufchan_buf :
                                      is_z_kronahW_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronahW_2_2_argbuf_r && is_z_kronahW_2_2_bufchan_buf[0]))
        is_z_kronahW_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_kronahW_2_2_argbuf_r) && (! is_z_kronahW_2_2_bufchan_buf[0])))
        is_z_kronahW_2_2_bufchan_buf <= is_z_kronahW_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_kronahW_2_destruct,MyDTInt_Bool) > [(is_z_kronahW_2_1,MyDTInt_Bool),
                                                                   (is_z_kronahW_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_kronahW_2_destruct_emitted;
  logic [1:0] is_z_kronahW_2_destruct_done;
  assign is_z_kronahW_2_1_d = (is_z_kronahW_2_destruct_d[0] && (! is_z_kronahW_2_destruct_emitted[0]));
  assign is_z_kronahW_2_2_d = (is_z_kronahW_2_destruct_d[0] && (! is_z_kronahW_2_destruct_emitted[1]));
  assign is_z_kronahW_2_destruct_done = (is_z_kronahW_2_destruct_emitted | ({is_z_kronahW_2_2_d[0],
                                                                             is_z_kronahW_2_1_d[0]} & {is_z_kronahW_2_2_r,
                                                                                                       is_z_kronahW_2_1_r}));
  assign is_z_kronahW_2_destruct_r = (& is_z_kronahW_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_2_destruct_emitted <= 2'd0;
    else
      is_z_kronahW_2_destruct_emitted <= (is_z_kronahW_2_destruct_r ? 2'd0 :
                                          is_z_kronahW_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronahW_3_2,MyDTInt_Bool) > (is_z_kronahW_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronahW_3_2_bufchan_d;
  logic is_z_kronahW_3_2_bufchan_r;
  assign is_z_kronahW_3_2_r = ((! is_z_kronahW_3_2_bufchan_d[0]) || is_z_kronahW_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_kronahW_3_2_r)
        is_z_kronahW_3_2_bufchan_d <= is_z_kronahW_3_2_d;
  MyDTInt_Bool_t is_z_kronahW_3_2_bufchan_buf;
  assign is_z_kronahW_3_2_bufchan_r = (! is_z_kronahW_3_2_bufchan_buf[0]);
  assign is_z_kronahW_3_2_argbuf_d = (is_z_kronahW_3_2_bufchan_buf[0] ? is_z_kronahW_3_2_bufchan_buf :
                                      is_z_kronahW_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronahW_3_2_argbuf_r && is_z_kronahW_3_2_bufchan_buf[0]))
        is_z_kronahW_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_kronahW_3_2_argbuf_r) && (! is_z_kronahW_3_2_bufchan_buf[0])))
        is_z_kronahW_3_2_bufchan_buf <= is_z_kronahW_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_kronahW_3_destruct,MyDTInt_Bool) > [(is_z_kronahW_3_1,MyDTInt_Bool),
                                                                   (is_z_kronahW_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_kronahW_3_destruct_emitted;
  logic [1:0] is_z_kronahW_3_destruct_done;
  assign is_z_kronahW_3_1_d = (is_z_kronahW_3_destruct_d[0] && (! is_z_kronahW_3_destruct_emitted[0]));
  assign is_z_kronahW_3_2_d = (is_z_kronahW_3_destruct_d[0] && (! is_z_kronahW_3_destruct_emitted[1]));
  assign is_z_kronahW_3_destruct_done = (is_z_kronahW_3_destruct_emitted | ({is_z_kronahW_3_2_d[0],
                                                                             is_z_kronahW_3_1_d[0]} & {is_z_kronahW_3_2_r,
                                                                                                       is_z_kronahW_3_1_r}));
  assign is_z_kronahW_3_destruct_r = (& is_z_kronahW_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_3_destruct_emitted <= 2'd0;
    else
      is_z_kronahW_3_destruct_emitted <= (is_z_kronahW_3_destruct_r ? 2'd0 :
                                          is_z_kronahW_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronahW_4_destruct,MyDTInt_Bool) > (is_z_kronahW_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronahW_4_destruct_bufchan_d;
  logic is_z_kronahW_4_destruct_bufchan_r;
  assign is_z_kronahW_4_destruct_r = ((! is_z_kronahW_4_destruct_bufchan_d[0]) || is_z_kronahW_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_kronahW_4_destruct_r)
        is_z_kronahW_4_destruct_bufchan_d <= is_z_kronahW_4_destruct_d;
  MyDTInt_Bool_t is_z_kronahW_4_destruct_bufchan_buf;
  assign is_z_kronahW_4_destruct_bufchan_r = (! is_z_kronahW_4_destruct_bufchan_buf[0]);
  assign is_z_kronahW_4_1_argbuf_d = (is_z_kronahW_4_destruct_bufchan_buf[0] ? is_z_kronahW_4_destruct_bufchan_buf :
                                      is_z_kronahW_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronahW_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronahW_4_1_argbuf_r && is_z_kronahW_4_destruct_bufchan_buf[0]))
        is_z_kronahW_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_kronahW_4_1_argbuf_r) && (! is_z_kronahW_4_destruct_bufchan_buf[0])))
        is_z_kronahW_4_destruct_bufchan_buf <= is_z_kronahW_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronai6_2_2,MyDTInt_Bool) > (is_z_kronai6_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronai6_2_2_bufchan_d;
  logic is_z_kronai6_2_2_bufchan_r;
  assign is_z_kronai6_2_2_r = ((! is_z_kronai6_2_2_bufchan_d[0]) || is_z_kronai6_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_kronai6_2_2_r)
        is_z_kronai6_2_2_bufchan_d <= is_z_kronai6_2_2_d;
  MyDTInt_Bool_t is_z_kronai6_2_2_bufchan_buf;
  assign is_z_kronai6_2_2_bufchan_r = (! is_z_kronai6_2_2_bufchan_buf[0]);
  assign is_z_kronai6_2_2_argbuf_d = (is_z_kronai6_2_2_bufchan_buf[0] ? is_z_kronai6_2_2_bufchan_buf :
                                      is_z_kronai6_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronai6_2_2_argbuf_r && is_z_kronai6_2_2_bufchan_buf[0]))
        is_z_kronai6_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_kronai6_2_2_argbuf_r) && (! is_z_kronai6_2_2_bufchan_buf[0])))
        is_z_kronai6_2_2_bufchan_buf <= is_z_kronai6_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_kronai6_2_destruct,MyDTInt_Bool) > [(is_z_kronai6_2_1,MyDTInt_Bool),
                                                                   (is_z_kronai6_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_kronai6_2_destruct_emitted;
  logic [1:0] is_z_kronai6_2_destruct_done;
  assign is_z_kronai6_2_1_d = (is_z_kronai6_2_destruct_d[0] && (! is_z_kronai6_2_destruct_emitted[0]));
  assign is_z_kronai6_2_2_d = (is_z_kronai6_2_destruct_d[0] && (! is_z_kronai6_2_destruct_emitted[1]));
  assign is_z_kronai6_2_destruct_done = (is_z_kronai6_2_destruct_emitted | ({is_z_kronai6_2_2_d[0],
                                                                             is_z_kronai6_2_1_d[0]} & {is_z_kronai6_2_2_r,
                                                                                                       is_z_kronai6_2_1_r}));
  assign is_z_kronai6_2_destruct_r = (& is_z_kronai6_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_2_destruct_emitted <= 2'd0;
    else
      is_z_kronai6_2_destruct_emitted <= (is_z_kronai6_2_destruct_r ? 2'd0 :
                                          is_z_kronai6_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronai6_3_2,MyDTInt_Bool) > (is_z_kronai6_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronai6_3_2_bufchan_d;
  logic is_z_kronai6_3_2_bufchan_r;
  assign is_z_kronai6_3_2_r = ((! is_z_kronai6_3_2_bufchan_d[0]) || is_z_kronai6_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_kronai6_3_2_r)
        is_z_kronai6_3_2_bufchan_d <= is_z_kronai6_3_2_d;
  MyDTInt_Bool_t is_z_kronai6_3_2_bufchan_buf;
  assign is_z_kronai6_3_2_bufchan_r = (! is_z_kronai6_3_2_bufchan_buf[0]);
  assign is_z_kronai6_3_2_argbuf_d = (is_z_kronai6_3_2_bufchan_buf[0] ? is_z_kronai6_3_2_bufchan_buf :
                                      is_z_kronai6_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronai6_3_2_argbuf_r && is_z_kronai6_3_2_bufchan_buf[0]))
        is_z_kronai6_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_kronai6_3_2_argbuf_r) && (! is_z_kronai6_3_2_bufchan_buf[0])))
        is_z_kronai6_3_2_bufchan_buf <= is_z_kronai6_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_kronai6_3_destruct,MyDTInt_Bool) > [(is_z_kronai6_3_1,MyDTInt_Bool),
                                                                   (is_z_kronai6_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_kronai6_3_destruct_emitted;
  logic [1:0] is_z_kronai6_3_destruct_done;
  assign is_z_kronai6_3_1_d = (is_z_kronai6_3_destruct_d[0] && (! is_z_kronai6_3_destruct_emitted[0]));
  assign is_z_kronai6_3_2_d = (is_z_kronai6_3_destruct_d[0] && (! is_z_kronai6_3_destruct_emitted[1]));
  assign is_z_kronai6_3_destruct_done = (is_z_kronai6_3_destruct_emitted | ({is_z_kronai6_3_2_d[0],
                                                                             is_z_kronai6_3_1_d[0]} & {is_z_kronai6_3_2_r,
                                                                                                       is_z_kronai6_3_1_r}));
  assign is_z_kronai6_3_destruct_r = (& is_z_kronai6_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_3_destruct_emitted <= 2'd0;
    else
      is_z_kronai6_3_destruct_emitted <= (is_z_kronai6_3_destruct_r ? 2'd0 :
                                          is_z_kronai6_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_kronai6_4_destruct,MyDTInt_Bool) > (is_z_kronai6_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_kronai6_4_destruct_bufchan_d;
  logic is_z_kronai6_4_destruct_bufchan_r;
  assign is_z_kronai6_4_destruct_r = ((! is_z_kronai6_4_destruct_bufchan_d[0]) || is_z_kronai6_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_kronai6_4_destruct_r)
        is_z_kronai6_4_destruct_bufchan_d <= is_z_kronai6_4_destruct_d;
  MyDTInt_Bool_t is_z_kronai6_4_destruct_bufchan_buf;
  assign is_z_kronai6_4_destruct_bufchan_r = (! is_z_kronai6_4_destruct_bufchan_buf[0]);
  assign is_z_kronai6_4_1_argbuf_d = (is_z_kronai6_4_destruct_bufchan_buf[0] ? is_z_kronai6_4_destruct_bufchan_buf :
                                      is_z_kronai6_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_kronai6_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_kronai6_4_1_argbuf_r && is_z_kronai6_4_destruct_bufchan_buf[0]))
        is_z_kronai6_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_kronai6_4_1_argbuf_r) && (! is_z_kronai6_4_destruct_bufchan_buf[0])))
        is_z_kronai6_4_destruct_bufchan_buf <= is_z_kronai6_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapahY_2_2,MyDTInt_Bool) > (is_z_mapahY_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapahY_2_2_bufchan_d;
  logic is_z_mapahY_2_2_bufchan_r;
  assign is_z_mapahY_2_2_r = ((! is_z_mapahY_2_2_bufchan_d[0]) || is_z_mapahY_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapahY_2_2_r)
        is_z_mapahY_2_2_bufchan_d <= is_z_mapahY_2_2_d;
  MyDTInt_Bool_t is_z_mapahY_2_2_bufchan_buf;
  assign is_z_mapahY_2_2_bufchan_r = (! is_z_mapahY_2_2_bufchan_buf[0]);
  assign is_z_mapahY_2_2_argbuf_d = (is_z_mapahY_2_2_bufchan_buf[0] ? is_z_mapahY_2_2_bufchan_buf :
                                     is_z_mapahY_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapahY_2_2_argbuf_r && is_z_mapahY_2_2_bufchan_buf[0]))
        is_z_mapahY_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapahY_2_2_argbuf_r) && (! is_z_mapahY_2_2_bufchan_buf[0])))
        is_z_mapahY_2_2_bufchan_buf <= is_z_mapahY_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapahY_2_destruct,MyDTInt_Bool) > [(is_z_mapahY_2_1,MyDTInt_Bool),
                                                                  (is_z_mapahY_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapahY_2_destruct_emitted;
  logic [1:0] is_z_mapahY_2_destruct_done;
  assign is_z_mapahY_2_1_d = (is_z_mapahY_2_destruct_d[0] && (! is_z_mapahY_2_destruct_emitted[0]));
  assign is_z_mapahY_2_2_d = (is_z_mapahY_2_destruct_d[0] && (! is_z_mapahY_2_destruct_emitted[1]));
  assign is_z_mapahY_2_destruct_done = (is_z_mapahY_2_destruct_emitted | ({is_z_mapahY_2_2_d[0],
                                                                           is_z_mapahY_2_1_d[0]} & {is_z_mapahY_2_2_r,
                                                                                                    is_z_mapahY_2_1_r}));
  assign is_z_mapahY_2_destruct_r = (& is_z_mapahY_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_2_destruct_emitted <= 2'd0;
    else
      is_z_mapahY_2_destruct_emitted <= (is_z_mapahY_2_destruct_r ? 2'd0 :
                                         is_z_mapahY_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapahY_3_2,MyDTInt_Bool) > (is_z_mapahY_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapahY_3_2_bufchan_d;
  logic is_z_mapahY_3_2_bufchan_r;
  assign is_z_mapahY_3_2_r = ((! is_z_mapahY_3_2_bufchan_d[0]) || is_z_mapahY_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapahY_3_2_r)
        is_z_mapahY_3_2_bufchan_d <= is_z_mapahY_3_2_d;
  MyDTInt_Bool_t is_z_mapahY_3_2_bufchan_buf;
  assign is_z_mapahY_3_2_bufchan_r = (! is_z_mapahY_3_2_bufchan_buf[0]);
  assign is_z_mapahY_3_2_argbuf_d = (is_z_mapahY_3_2_bufchan_buf[0] ? is_z_mapahY_3_2_bufchan_buf :
                                     is_z_mapahY_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapahY_3_2_argbuf_r && is_z_mapahY_3_2_bufchan_buf[0]))
        is_z_mapahY_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapahY_3_2_argbuf_r) && (! is_z_mapahY_3_2_bufchan_buf[0])))
        is_z_mapahY_3_2_bufchan_buf <= is_z_mapahY_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapahY_3_destruct,MyDTInt_Bool) > [(is_z_mapahY_3_1,MyDTInt_Bool),
                                                                  (is_z_mapahY_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapahY_3_destruct_emitted;
  logic [1:0] is_z_mapahY_3_destruct_done;
  assign is_z_mapahY_3_1_d = (is_z_mapahY_3_destruct_d[0] && (! is_z_mapahY_3_destruct_emitted[0]));
  assign is_z_mapahY_3_2_d = (is_z_mapahY_3_destruct_d[0] && (! is_z_mapahY_3_destruct_emitted[1]));
  assign is_z_mapahY_3_destruct_done = (is_z_mapahY_3_destruct_emitted | ({is_z_mapahY_3_2_d[0],
                                                                           is_z_mapahY_3_1_d[0]} & {is_z_mapahY_3_2_r,
                                                                                                    is_z_mapahY_3_1_r}));
  assign is_z_mapahY_3_destruct_r = (& is_z_mapahY_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_3_destruct_emitted <= 2'd0;
    else
      is_z_mapahY_3_destruct_emitted <= (is_z_mapahY_3_destruct_r ? 2'd0 :
                                         is_z_mapahY_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapahY_4_destruct,MyDTInt_Bool) > (is_z_mapahY_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapahY_4_destruct_bufchan_d;
  logic is_z_mapahY_4_destruct_bufchan_r;
  assign is_z_mapahY_4_destruct_r = ((! is_z_mapahY_4_destruct_bufchan_d[0]) || is_z_mapahY_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_mapahY_4_destruct_r)
        is_z_mapahY_4_destruct_bufchan_d <= is_z_mapahY_4_destruct_d;
  MyDTInt_Bool_t is_z_mapahY_4_destruct_bufchan_buf;
  assign is_z_mapahY_4_destruct_bufchan_r = (! is_z_mapahY_4_destruct_bufchan_buf[0]);
  assign is_z_mapahY_4_1_argbuf_d = (is_z_mapahY_4_destruct_bufchan_buf[0] ? is_z_mapahY_4_destruct_bufchan_buf :
                                     is_z_mapahY_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapahY_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapahY_4_1_argbuf_r && is_z_mapahY_4_destruct_bufchan_buf[0]))
        is_z_mapahY_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_mapahY_4_1_argbuf_r) && (! is_z_mapahY_4_destruct_bufchan_buf[0])))
        is_z_mapahY_4_destruct_bufchan_buf <= is_z_mapahY_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapai9_2_2,MyDTInt_Bool) > (is_z_mapai9_2_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapai9_2_2_bufchan_d;
  logic is_z_mapai9_2_2_bufchan_r;
  assign is_z_mapai9_2_2_r = ((! is_z_mapai9_2_2_bufchan_d[0]) || is_z_mapai9_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_2_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapai9_2_2_r)
        is_z_mapai9_2_2_bufchan_d <= is_z_mapai9_2_2_d;
  MyDTInt_Bool_t is_z_mapai9_2_2_bufchan_buf;
  assign is_z_mapai9_2_2_bufchan_r = (! is_z_mapai9_2_2_bufchan_buf[0]);
  assign is_z_mapai9_2_2_argbuf_d = (is_z_mapai9_2_2_bufchan_buf[0] ? is_z_mapai9_2_2_bufchan_buf :
                                     is_z_mapai9_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_2_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapai9_2_2_argbuf_r && is_z_mapai9_2_2_bufchan_buf[0]))
        is_z_mapai9_2_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapai9_2_2_argbuf_r) && (! is_z_mapai9_2_2_bufchan_buf[0])))
        is_z_mapai9_2_2_bufchan_buf <= is_z_mapai9_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapai9_2_destruct,MyDTInt_Bool) > [(is_z_mapai9_2_1,MyDTInt_Bool),
                                                                  (is_z_mapai9_2_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapai9_2_destruct_emitted;
  logic [1:0] is_z_mapai9_2_destruct_done;
  assign is_z_mapai9_2_1_d = (is_z_mapai9_2_destruct_d[0] && (! is_z_mapai9_2_destruct_emitted[0]));
  assign is_z_mapai9_2_2_d = (is_z_mapai9_2_destruct_d[0] && (! is_z_mapai9_2_destruct_emitted[1]));
  assign is_z_mapai9_2_destruct_done = (is_z_mapai9_2_destruct_emitted | ({is_z_mapai9_2_2_d[0],
                                                                           is_z_mapai9_2_1_d[0]} & {is_z_mapai9_2_2_r,
                                                                                                    is_z_mapai9_2_1_r}));
  assign is_z_mapai9_2_destruct_r = (& is_z_mapai9_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_2_destruct_emitted <= 2'd0;
    else
      is_z_mapai9_2_destruct_emitted <= (is_z_mapai9_2_destruct_r ? 2'd0 :
                                         is_z_mapai9_2_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapai9_3_2,MyDTInt_Bool) > (is_z_mapai9_3_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapai9_3_2_bufchan_d;
  logic is_z_mapai9_3_2_bufchan_r;
  assign is_z_mapai9_3_2_r = ((! is_z_mapai9_3_2_bufchan_d[0]) || is_z_mapai9_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_3_2_bufchan_d <= 1'd0;
    else
      if (is_z_mapai9_3_2_r)
        is_z_mapai9_3_2_bufchan_d <= is_z_mapai9_3_2_d;
  MyDTInt_Bool_t is_z_mapai9_3_2_bufchan_buf;
  assign is_z_mapai9_3_2_bufchan_r = (! is_z_mapai9_3_2_bufchan_buf[0]);
  assign is_z_mapai9_3_2_argbuf_d = (is_z_mapai9_3_2_bufchan_buf[0] ? is_z_mapai9_3_2_bufchan_buf :
                                     is_z_mapai9_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_3_2_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapai9_3_2_argbuf_r && is_z_mapai9_3_2_bufchan_buf[0]))
        is_z_mapai9_3_2_bufchan_buf <= 1'd0;
      else if (((! is_z_mapai9_3_2_argbuf_r) && (! is_z_mapai9_3_2_bufchan_buf[0])))
        is_z_mapai9_3_2_bufchan_buf <= is_z_mapai9_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Bool) : (is_z_mapai9_3_destruct,MyDTInt_Bool) > [(is_z_mapai9_3_1,MyDTInt_Bool),
                                                                  (is_z_mapai9_3_2,MyDTInt_Bool)] */
  logic [1:0] is_z_mapai9_3_destruct_emitted;
  logic [1:0] is_z_mapai9_3_destruct_done;
  assign is_z_mapai9_3_1_d = (is_z_mapai9_3_destruct_d[0] && (! is_z_mapai9_3_destruct_emitted[0]));
  assign is_z_mapai9_3_2_d = (is_z_mapai9_3_destruct_d[0] && (! is_z_mapai9_3_destruct_emitted[1]));
  assign is_z_mapai9_3_destruct_done = (is_z_mapai9_3_destruct_emitted | ({is_z_mapai9_3_2_d[0],
                                                                           is_z_mapai9_3_1_d[0]} & {is_z_mapai9_3_2_r,
                                                                                                    is_z_mapai9_3_1_r}));
  assign is_z_mapai9_3_destruct_r = (& is_z_mapai9_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_3_destruct_emitted <= 2'd0;
    else
      is_z_mapai9_3_destruct_emitted <= (is_z_mapai9_3_destruct_r ? 2'd0 :
                                         is_z_mapai9_3_destruct_done);
  
  /* buf (Ty MyDTInt_Bool) : (is_z_mapai9_4_destruct,MyDTInt_Bool) > (is_z_mapai9_4_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t is_z_mapai9_4_destruct_bufchan_d;
  logic is_z_mapai9_4_destruct_bufchan_r;
  assign is_z_mapai9_4_destruct_r = ((! is_z_mapai9_4_destruct_bufchan_d[0]) || is_z_mapai9_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_4_destruct_bufchan_d <= 1'd0;
    else
      if (is_z_mapai9_4_destruct_r)
        is_z_mapai9_4_destruct_bufchan_d <= is_z_mapai9_4_destruct_d;
  MyDTInt_Bool_t is_z_mapai9_4_destruct_bufchan_buf;
  assign is_z_mapai9_4_destruct_bufchan_r = (! is_z_mapai9_4_destruct_bufchan_buf[0]);
  assign is_z_mapai9_4_1_argbuf_d = (is_z_mapai9_4_destruct_bufchan_buf[0] ? is_z_mapai9_4_destruct_bufchan_buf :
                                     is_z_mapai9_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) is_z_mapai9_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((is_z_mapai9_4_1_argbuf_r && is_z_mapai9_4_destruct_bufchan_buf[0]))
        is_z_mapai9_4_destruct_bufchan_buf <= 1'd0;
      else if (((! is_z_mapai9_4_1_argbuf_r) && (! is_z_mapai9_4_destruct_bufchan_buf[0])))
        is_z_mapai9_4_destruct_bufchan_buf <= is_z_mapai9_4_destruct_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet13_1_1QNode_Int,QTree_Int) > [(q1ai1_destruct,Pointer_QTree_Int),
                                                                    (q2ai2_destruct,Pointer_QTree_Int),
                                                                    (q3ai3_destruct,Pointer_QTree_Int),
                                                                    (q4ai4_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet13_1_1QNode_Int_emitted;
  logic [3:0] lizzieLet13_1_1QNode_Int_done;
  assign q1ai1_destruct_d = {lizzieLet13_1_1QNode_Int_d[18:3],
                             (lizzieLet13_1_1QNode_Int_d[0] && (! lizzieLet13_1_1QNode_Int_emitted[0]))};
  assign q2ai2_destruct_d = {lizzieLet13_1_1QNode_Int_d[34:19],
                             (lizzieLet13_1_1QNode_Int_d[0] && (! lizzieLet13_1_1QNode_Int_emitted[1]))};
  assign q3ai3_destruct_d = {lizzieLet13_1_1QNode_Int_d[50:35],
                             (lizzieLet13_1_1QNode_Int_d[0] && (! lizzieLet13_1_1QNode_Int_emitted[2]))};
  assign q4ai4_destruct_d = {lizzieLet13_1_1QNode_Int_d[66:51],
                             (lizzieLet13_1_1QNode_Int_d[0] && (! lizzieLet13_1_1QNode_Int_emitted[3]))};
  assign lizzieLet13_1_1QNode_Int_done = (lizzieLet13_1_1QNode_Int_emitted | ({q4ai4_destruct_d[0],
                                                                               q3ai3_destruct_d[0],
                                                                               q2ai2_destruct_d[0],
                                                                               q1ai1_destruct_d[0]} & {q4ai4_destruct_r,
                                                                                                       q3ai3_destruct_r,
                                                                                                       q2ai2_destruct_r,
                                                                                                       q1ai1_destruct_r}));
  assign lizzieLet13_1_1QNode_Int_r = (& lizzieLet13_1_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet13_1_1QNode_Int_emitted <= (lizzieLet13_1_1QNode_Int_r ? 4'd0 :
                                           lizzieLet13_1_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet13_1_1QVal_Int,QTree_Int) > [(vai0_destruct,Int)] */
  assign vai0_destruct_d = {lizzieLet13_1_1QVal_Int_d[34:3],
                            lizzieLet13_1_1QVal_Int_d[0]};
  assign lizzieLet13_1_1QVal_Int_r = vai0_destruct_r;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet13_1_2,QTree_Int) (lizzieLet13_1_1,QTree_Int) > [(_32,QTree_Int),
                                                                                  (lizzieLet13_1_1QVal_Int,QTree_Int),
                                                                                  (lizzieLet13_1_1QNode_Int,QTree_Int),
                                                                                  (_31,QTree_Int)] */
  logic [3:0] lizzieLet13_1_1_onehotd;
  always_comb
    if ((lizzieLet13_1_2_d[0] && lizzieLet13_1_1_d[0]))
      unique case (lizzieLet13_1_2_d[2:1])
        2'd0: lizzieLet13_1_1_onehotd = 4'd1;
        2'd1: lizzieLet13_1_1_onehotd = 4'd2;
        2'd2: lizzieLet13_1_1_onehotd = 4'd4;
        2'd3: lizzieLet13_1_1_onehotd = 4'd8;
        default: lizzieLet13_1_1_onehotd = 4'd0;
      endcase
    else lizzieLet13_1_1_onehotd = 4'd0;
  assign _32_d = {lizzieLet13_1_1_d[66:1],
                  lizzieLet13_1_1_onehotd[0]};
  assign lizzieLet13_1_1QVal_Int_d = {lizzieLet13_1_1_d[66:1],
                                      lizzieLet13_1_1_onehotd[1]};
  assign lizzieLet13_1_1QNode_Int_d = {lizzieLet13_1_1_d[66:1],
                                       lizzieLet13_1_1_onehotd[2]};
  assign _31_d = {lizzieLet13_1_1_d[66:1],
                  lizzieLet13_1_1_onehotd[3]};
  assign lizzieLet13_1_1_r = (| (lizzieLet13_1_1_onehotd & {_31_r,
                                                            lizzieLet13_1_1QNode_Int_r,
                                                            lizzieLet13_1_1QVal_Int_r,
                                                            _32_r}));
  assign lizzieLet13_1_2_r = lizzieLet13_1_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet13_1_3,QTree_Int) (f_mapahZ_goMux_mux,MyDTInt_Int) > [(_30,MyDTInt_Int),
                                                                                         (lizzieLet13_1_3QVal_Int,MyDTInt_Int),
                                                                                         (lizzieLet13_1_3QNode_Int,MyDTInt_Int),
                                                                                         (_29,MyDTInt_Int)] */
  logic [3:0] f_mapahZ_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_3_d[0] && f_mapahZ_goMux_mux_d[0]))
      unique case (lizzieLet13_1_3_d[2:1])
        2'd0: f_mapahZ_goMux_mux_onehotd = 4'd1;
        2'd1: f_mapahZ_goMux_mux_onehotd = 4'd2;
        2'd2: f_mapahZ_goMux_mux_onehotd = 4'd4;
        2'd3: f_mapahZ_goMux_mux_onehotd = 4'd8;
        default: f_mapahZ_goMux_mux_onehotd = 4'd0;
      endcase
    else f_mapahZ_goMux_mux_onehotd = 4'd0;
  assign _30_d = f_mapahZ_goMux_mux_onehotd[0];
  assign lizzieLet13_1_3QVal_Int_d = f_mapahZ_goMux_mux_onehotd[1];
  assign lizzieLet13_1_3QNode_Int_d = f_mapahZ_goMux_mux_onehotd[2];
  assign _29_d = f_mapahZ_goMux_mux_onehotd[3];
  assign f_mapahZ_goMux_mux_r = (| (f_mapahZ_goMux_mux_onehotd & {_29_r,
                                                                  lizzieLet13_1_3QNode_Int_r,
                                                                  lizzieLet13_1_3QVal_Int_r,
                                                                  _30_r}));
  assign lizzieLet13_1_3_r = f_mapahZ_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet13_1_3QNode_Int,MyDTInt_Int) > [(lizzieLet13_1_3QNode_Int_1,MyDTInt_Int),
                                                                  (lizzieLet13_1_3QNode_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet13_1_3QNode_Int_emitted;
  logic [1:0] lizzieLet13_1_3QNode_Int_done;
  assign lizzieLet13_1_3QNode_Int_1_d = (lizzieLet13_1_3QNode_Int_d[0] && (! lizzieLet13_1_3QNode_Int_emitted[0]));
  assign lizzieLet13_1_3QNode_Int_2_d = (lizzieLet13_1_3QNode_Int_d[0] && (! lizzieLet13_1_3QNode_Int_emitted[1]));
  assign lizzieLet13_1_3QNode_Int_done = (lizzieLet13_1_3QNode_Int_emitted | ({lizzieLet13_1_3QNode_Int_2_d[0],
                                                                               lizzieLet13_1_3QNode_Int_1_d[0]} & {lizzieLet13_1_3QNode_Int_2_r,
                                                                                                                   lizzieLet13_1_3QNode_Int_1_r}));
  assign lizzieLet13_1_3QNode_Int_r = (& lizzieLet13_1_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_3QNode_Int_emitted <= (lizzieLet13_1_3QNode_Int_r ? 2'd0 :
                                           lizzieLet13_1_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet13_1_3QNode_Int_2,MyDTInt_Int) > (lizzieLet13_1_3QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_2_bufchan_d;
  logic lizzieLet13_1_3QNode_Int_2_bufchan_r;
  assign lizzieLet13_1_3QNode_Int_2_r = ((! lizzieLet13_1_3QNode_Int_2_bufchan_d[0]) || lizzieLet13_1_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_3QNode_Int_2_r)
        lizzieLet13_1_3QNode_Int_2_bufchan_d <= lizzieLet13_1_3QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet13_1_3QNode_Int_2_bufchan_buf;
  assign lizzieLet13_1_3QNode_Int_2_bufchan_r = (! lizzieLet13_1_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_3QNode_Int_2_argbuf_d = (lizzieLet13_1_3QNode_Int_2_bufchan_buf[0] ? lizzieLet13_1_3QNode_Int_2_bufchan_buf :
                                                lizzieLet13_1_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_3QNode_Int_2_argbuf_r && lizzieLet13_1_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_1_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_3QNode_Int_2_argbuf_r) && (! lizzieLet13_1_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_1_3QNode_Int_2_bufchan_buf <= lizzieLet13_1_3QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet13_1_3QVal_Int,MyDTInt_Int) > (lizzieLet13_1_3QVal_Int_1_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet13_1_3QVal_Int_bufchan_d;
  logic lizzieLet13_1_3QVal_Int_bufchan_r;
  assign lizzieLet13_1_3QVal_Int_r = ((! lizzieLet13_1_3QVal_Int_bufchan_d[0]) || lizzieLet13_1_3QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_3QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_3QVal_Int_r)
        lizzieLet13_1_3QVal_Int_bufchan_d <= lizzieLet13_1_3QVal_Int_d;
  MyDTInt_Int_t lizzieLet13_1_3QVal_Int_bufchan_buf;
  assign lizzieLet13_1_3QVal_Int_bufchan_r = (! lizzieLet13_1_3QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_3QVal_Int_1_argbuf_d = (lizzieLet13_1_3QVal_Int_bufchan_buf[0] ? lizzieLet13_1_3QVal_Int_bufchan_buf :
                                               lizzieLet13_1_3QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_3QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_3QVal_Int_1_argbuf_r && lizzieLet13_1_3QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_3QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_3QVal_Int_1_argbuf_r) && (! lizzieLet13_1_3QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_3QVal_Int_bufchan_buf <= lizzieLet13_1_3QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet13_1_4,QTree_Int) (go_12_goMux_data,Go) > [(lizzieLet13_1_4QNone_Int,Go),
                                                                     (lizzieLet13_1_4QVal_Int,Go),
                                                                     (lizzieLet13_1_4QNode_Int,Go),
                                                                     (lizzieLet13_1_4QError_Int,Go)] */
  logic [3:0] go_12_goMux_data_onehotd;
  always_comb
    if ((lizzieLet13_1_4_d[0] && go_12_goMux_data_d[0]))
      unique case (lizzieLet13_1_4_d[2:1])
        2'd0: go_12_goMux_data_onehotd = 4'd1;
        2'd1: go_12_goMux_data_onehotd = 4'd2;
        2'd2: go_12_goMux_data_onehotd = 4'd4;
        2'd3: go_12_goMux_data_onehotd = 4'd8;
        default: go_12_goMux_data_onehotd = 4'd0;
      endcase
    else go_12_goMux_data_onehotd = 4'd0;
  assign lizzieLet13_1_4QNone_Int_d = go_12_goMux_data_onehotd[0];
  assign lizzieLet13_1_4QVal_Int_d = go_12_goMux_data_onehotd[1];
  assign lizzieLet13_1_4QNode_Int_d = go_12_goMux_data_onehotd[2];
  assign lizzieLet13_1_4QError_Int_d = go_12_goMux_data_onehotd[3];
  assign go_12_goMux_data_r = (| (go_12_goMux_data_onehotd & {lizzieLet13_1_4QError_Int_r,
                                                              lizzieLet13_1_4QNode_Int_r,
                                                              lizzieLet13_1_4QVal_Int_r,
                                                              lizzieLet13_1_4QNone_Int_r}));
  assign lizzieLet13_1_4_r = go_12_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet13_1_4QError_Int,Go) > [(lizzieLet13_1_4QError_Int_1,Go),
                                                 (lizzieLet13_1_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet13_1_4QError_Int_emitted;
  logic [1:0] lizzieLet13_1_4QError_Int_done;
  assign lizzieLet13_1_4QError_Int_1_d = (lizzieLet13_1_4QError_Int_d[0] && (! lizzieLet13_1_4QError_Int_emitted[0]));
  assign lizzieLet13_1_4QError_Int_2_d = (lizzieLet13_1_4QError_Int_d[0] && (! lizzieLet13_1_4QError_Int_emitted[1]));
  assign lizzieLet13_1_4QError_Int_done = (lizzieLet13_1_4QError_Int_emitted | ({lizzieLet13_1_4QError_Int_2_d[0],
                                                                                 lizzieLet13_1_4QError_Int_1_d[0]} & {lizzieLet13_1_4QError_Int_2_r,
                                                                                                                      lizzieLet13_1_4QError_Int_1_r}));
  assign lizzieLet13_1_4QError_Int_r = (& lizzieLet13_1_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_4QError_Int_emitted <= (lizzieLet13_1_4QError_Int_r ? 2'd0 :
                                            lizzieLet13_1_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet13_1_4QError_Int_1,Go)] > (lizzieLet13_1_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet13_1_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet13_1_4QError_Int_1_d[0]}), lizzieLet13_1_4QError_Int_1_d);
  assign {lizzieLet13_1_4QError_Int_1_r} = {1 {(lizzieLet13_1_4QError_Int_1QError_Int_r && lizzieLet13_1_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_1_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet16_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet13_1_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet13_1_4QError_Int_1QError_Int_r = ((! lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet13_1_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet13_1_4QError_Int_1QError_Int_r)
        lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d <= lizzieLet13_1_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet13_1_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet16_1_argbuf_d = (lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf :
                                   lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet16_1_argbuf_r && lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet16_1_argbuf_r) && (! lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet13_1_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet13_1_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_1_4QError_Int_2,Go) > (lizzieLet13_1_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet13_1_4QError_Int_2_bufchan_d;
  logic lizzieLet13_1_4QError_Int_2_bufchan_r;
  assign lizzieLet13_1_4QError_Int_2_r = ((! lizzieLet13_1_4QError_Int_2_bufchan_d[0]) || lizzieLet13_1_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_4QError_Int_2_r)
        lizzieLet13_1_4QError_Int_2_bufchan_d <= lizzieLet13_1_4QError_Int_2_d;
  Go_t lizzieLet13_1_4QError_Int_2_bufchan_buf;
  assign lizzieLet13_1_4QError_Int_2_bufchan_r = (! lizzieLet13_1_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_4QError_Int_2_argbuf_d = (lizzieLet13_1_4QError_Int_2_bufchan_buf[0] ? lizzieLet13_1_4QError_Int_2_bufchan_buf :
                                                 lizzieLet13_1_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_4QError_Int_2_argbuf_r && lizzieLet13_1_4QError_Int_2_bufchan_buf[0]))
        lizzieLet13_1_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_4QError_Int_2_argbuf_r) && (! lizzieLet13_1_4QError_Int_2_bufchan_buf[0])))
        lizzieLet13_1_4QError_Int_2_bufchan_buf <= lizzieLet13_1_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_1_4QNode_Int,Go) > (lizzieLet13_1_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet13_1_4QNode_Int_bufchan_d;
  logic lizzieLet13_1_4QNode_Int_bufchan_r;
  assign lizzieLet13_1_4QNode_Int_r = ((! lizzieLet13_1_4QNode_Int_bufchan_d[0]) || lizzieLet13_1_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_4QNode_Int_r)
        lizzieLet13_1_4QNode_Int_bufchan_d <= lizzieLet13_1_4QNode_Int_d;
  Go_t lizzieLet13_1_4QNode_Int_bufchan_buf;
  assign lizzieLet13_1_4QNode_Int_bufchan_r = (! lizzieLet13_1_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet13_1_4QNode_Int_1_argbuf_d = (lizzieLet13_1_4QNode_Int_bufchan_buf[0] ? lizzieLet13_1_4QNode_Int_bufchan_buf :
                                                lizzieLet13_1_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_4QNode_Int_1_argbuf_r && lizzieLet13_1_4QNode_Int_bufchan_buf[0]))
        lizzieLet13_1_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_4QNode_Int_1_argbuf_r) && (! lizzieLet13_1_4QNode_Int_bufchan_buf[0])))
        lizzieLet13_1_4QNode_Int_bufchan_buf <= lizzieLet13_1_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet13_1_4QNone_Int,Go) > [(lizzieLet13_1_4QNone_Int_1,Go),
                                                (lizzieLet13_1_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet13_1_4QNone_Int_emitted;
  logic [1:0] lizzieLet13_1_4QNone_Int_done;
  assign lizzieLet13_1_4QNone_Int_1_d = (lizzieLet13_1_4QNone_Int_d[0] && (! lizzieLet13_1_4QNone_Int_emitted[0]));
  assign lizzieLet13_1_4QNone_Int_2_d = (lizzieLet13_1_4QNone_Int_d[0] && (! lizzieLet13_1_4QNone_Int_emitted[1]));
  assign lizzieLet13_1_4QNone_Int_done = (lizzieLet13_1_4QNone_Int_emitted | ({lizzieLet13_1_4QNone_Int_2_d[0],
                                                                               lizzieLet13_1_4QNone_Int_1_d[0]} & {lizzieLet13_1_4QNone_Int_2_r,
                                                                                                                   lizzieLet13_1_4QNone_Int_1_r}));
  assign lizzieLet13_1_4QNone_Int_r = (& lizzieLet13_1_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_4QNone_Int_emitted <= (lizzieLet13_1_4QNone_Int_r ? 2'd0 :
                                           lizzieLet13_1_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet13_1_4QNone_Int_1,Go)] > (lizzieLet13_1_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet13_1_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet13_1_4QNone_Int_1_d[0]}), lizzieLet13_1_4QNone_Int_1_d);
  assign {lizzieLet13_1_4QNone_Int_1_r} = {1 {(lizzieLet13_1_4QNone_Int_1QNone_Int_r && lizzieLet13_1_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet13_1_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet14_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet13_1_4QNone_Int_1QNone_Int_r = ((! lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet13_1_4QNone_Int_1QNone_Int_r)
        lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet13_1_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet14_1_argbuf_d = (lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf :
                                   lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet14_1_argbuf_r && lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet14_1_argbuf_r) && (! lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet13_1_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet13_1_4QNone_Int_2,Go) > (lizzieLet13_1_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet13_1_4QNone_Int_2_bufchan_d;
  logic lizzieLet13_1_4QNone_Int_2_bufchan_r;
  assign lizzieLet13_1_4QNone_Int_2_r = ((! lizzieLet13_1_4QNone_Int_2_bufchan_d[0]) || lizzieLet13_1_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_4QNone_Int_2_r)
        lizzieLet13_1_4QNone_Int_2_bufchan_d <= lizzieLet13_1_4QNone_Int_2_d;
  Go_t lizzieLet13_1_4QNone_Int_2_bufchan_buf;
  assign lizzieLet13_1_4QNone_Int_2_bufchan_r = (! lizzieLet13_1_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_4QNone_Int_2_argbuf_d = (lizzieLet13_1_4QNone_Int_2_bufchan_buf[0] ? lizzieLet13_1_4QNone_Int_2_bufchan_buf :
                                                lizzieLet13_1_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_4QNone_Int_2_argbuf_r && lizzieLet13_1_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet13_1_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_4QNone_Int_2_argbuf_r) && (! lizzieLet13_1_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet13_1_4QNone_Int_2_bufchan_buf <= lizzieLet13_1_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet13_1_4QNone_Int_2_argbuf,Go),
                           (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf,Go),
                           (lizzieLet13_1_4QVal_Int_2_argbuf,Go),
                           (lizzieLet13_1_4QError_Int_2_argbuf,Go)] > (go_17_goMux_choice,C4) (go_17_goMux_data,Go) */
  logic [3:0] lizzieLet13_1_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet13_1_4QNone_Int_2_argbuf_select_d = ((| lizzieLet13_1_4QNone_Int_2_argbuf_select_q) ? lizzieLet13_1_4QNone_Int_2_argbuf_select_q :
                                                       (lizzieLet13_1_4QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                        (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_d[0] ? 4'd2 :
                                                         (lizzieLet13_1_4QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                          (lizzieLet13_1_4QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                           4'd0)))));
  logic [3:0] lizzieLet13_1_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet13_1_4QNone_Int_2_argbuf_select_q <= (lizzieLet13_1_4QNone_Int_2_argbuf_done ? 4'd0 :
                                                     lizzieLet13_1_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet13_1_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet13_1_4QNone_Int_2_argbuf_emit_q <= (lizzieLet13_1_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                   lizzieLet13_1_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet13_1_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet13_1_4QNone_Int_2_argbuf_emit_d = (lizzieLet13_1_4QNone_Int_2_argbuf_emit_q | ({go_17_goMux_choice_d[0],
                                                                                                  go_17_goMux_data_d[0]} & {go_17_goMux_choice_r,
                                                                                                                            go_17_goMux_data_r}));
  logic lizzieLet13_1_4QNone_Int_2_argbuf_done;
  assign lizzieLet13_1_4QNone_Int_2_argbuf_done = (& lizzieLet13_1_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet13_1_4QError_Int_2_argbuf_r,
          lizzieLet13_1_4QVal_Int_2_argbuf_r,
          lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_r,
          lizzieLet13_1_4QNone_Int_2_argbuf_r} = (lizzieLet13_1_4QNone_Int_2_argbuf_done ? lizzieLet13_1_4QNone_Int_2_argbuf_select_d :
                                                  4'd0);
  assign go_17_goMux_data_d = ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet13_1_4QNone_Int_2_argbuf_d :
                               ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_d :
                                ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet13_1_4QVal_Int_2_argbuf_d :
                                 ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet13_1_4QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_17_goMux_choice_d = ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet13_1_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet13_1_4QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet13_1_4QVal_Int,Go) > [(lizzieLet13_1_4QVal_Int_1,Go),
                                               (lizzieLet13_1_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet13_1_4QVal_Int_emitted;
  logic [1:0] lizzieLet13_1_4QVal_Int_done;
  assign lizzieLet13_1_4QVal_Int_1_d = (lizzieLet13_1_4QVal_Int_d[0] && (! lizzieLet13_1_4QVal_Int_emitted[0]));
  assign lizzieLet13_1_4QVal_Int_2_d = (lizzieLet13_1_4QVal_Int_d[0] && (! lizzieLet13_1_4QVal_Int_emitted[1]));
  assign lizzieLet13_1_4QVal_Int_done = (lizzieLet13_1_4QVal_Int_emitted | ({lizzieLet13_1_4QVal_Int_2_d[0],
                                                                             lizzieLet13_1_4QVal_Int_1_d[0]} & {lizzieLet13_1_4QVal_Int_2_r,
                                                                                                                lizzieLet13_1_4QVal_Int_1_r}));
  assign lizzieLet13_1_4QVal_Int_r = (& lizzieLet13_1_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_4QVal_Int_emitted <= (lizzieLet13_1_4QVal_Int_r ? 2'd0 :
                                          lizzieLet13_1_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet13_1_4QVal_Int_1,Go) > (lizzieLet13_1_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet13_1_4QVal_Int_1_bufchan_d;
  logic lizzieLet13_1_4QVal_Int_1_bufchan_r;
  assign lizzieLet13_1_4QVal_Int_1_r = ((! lizzieLet13_1_4QVal_Int_1_bufchan_d[0]) || lizzieLet13_1_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_4QVal_Int_1_r)
        lizzieLet13_1_4QVal_Int_1_bufchan_d <= lizzieLet13_1_4QVal_Int_1_d;
  Go_t lizzieLet13_1_4QVal_Int_1_bufchan_buf;
  assign lizzieLet13_1_4QVal_Int_1_bufchan_r = (! lizzieLet13_1_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet13_1_4QVal_Int_1_argbuf_d = (lizzieLet13_1_4QVal_Int_1_bufchan_buf[0] ? lizzieLet13_1_4QVal_Int_1_bufchan_buf :
                                               lizzieLet13_1_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_4QVal_Int_1_argbuf_r && lizzieLet13_1_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet13_1_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_4QVal_Int_1_argbuf_r) && (! lizzieLet13_1_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet13_1_4QVal_Int_1_bufchan_buf <= lizzieLet13_1_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int,
      Dcon TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int) : [(lizzieLet13_1_4QVal_Int_1_argbuf,Go),
                                                                                                             (lizzieLet13_1_7QVal_Int_1_argbuf,Pointer_QTree_Int),
                                                                                                             (lizzieLet13_1_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                                                                                             (lizzieLet13_1_8QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                                                                                             (vai0_1_argbuf,Int),
                                                                                                             (lizzieLet13_1_6QVal_Int_1_argbuf,MyDTInt_Bool),
                                                                                                             (lizzieLet13_1_3QVal_Int_1_argbuf,MyDTInt_Int)] > (f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1,TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int) */
  assign \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d  = TupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_dc((& {lizzieLet13_1_4QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                                                                         lizzieLet13_1_7QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                                                                         lizzieLet13_1_5QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                                                                         lizzieLet13_1_8QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                                                                         vai0_1_argbuf_d[0],
                                                                                                                                                                                                                                         lizzieLet13_1_6QVal_Int_1_argbuf_d[0],
                                                                                                                                                                                                                                         lizzieLet13_1_3QVal_Int_1_argbuf_d[0]}), lizzieLet13_1_4QVal_Int_1_argbuf_d, lizzieLet13_1_7QVal_Int_1_argbuf_d, lizzieLet13_1_5QVal_Int_1_argbuf_d, lizzieLet13_1_8QVal_Int_1_argbuf_d, vai0_1_argbuf_d, lizzieLet13_1_6QVal_Int_1_argbuf_d, lizzieLet13_1_3QVal_Int_1_argbuf_d);
  assign {lizzieLet13_1_4QVal_Int_1_argbuf_r,
          lizzieLet13_1_7QVal_Int_1_argbuf_r,
          lizzieLet13_1_5QVal_Int_1_argbuf_r,
          lizzieLet13_1_8QVal_Int_1_argbuf_r,
          vai0_1_argbuf_r,
          lizzieLet13_1_6QVal_Int_1_argbuf_r,
          lizzieLet13_1_3QVal_Int_1_argbuf_r} = {7 {(\f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_r  && \f'_f'_Int_Int_Int_IntTupGo___Pointer_QTree_Int___MyDTInt_Bool___MyDTInt_Int_Int___Int___MyDTInt_Bool___MyDTInt_Int_1_d [0])}};
  
  /* buf (Ty Go) : (lizzieLet13_1_4QVal_Int_2,Go) > (lizzieLet13_1_4QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet13_1_4QVal_Int_2_bufchan_d;
  logic lizzieLet13_1_4QVal_Int_2_bufchan_r;
  assign lizzieLet13_1_4QVal_Int_2_r = ((! lizzieLet13_1_4QVal_Int_2_bufchan_d[0]) || lizzieLet13_1_4QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_4QVal_Int_2_r)
        lizzieLet13_1_4QVal_Int_2_bufchan_d <= lizzieLet13_1_4QVal_Int_2_d;
  Go_t lizzieLet13_1_4QVal_Int_2_bufchan_buf;
  assign lizzieLet13_1_4QVal_Int_2_bufchan_r = (! lizzieLet13_1_4QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_4QVal_Int_2_argbuf_d = (lizzieLet13_1_4QVal_Int_2_bufchan_buf[0] ? lizzieLet13_1_4QVal_Int_2_bufchan_buf :
                                               lizzieLet13_1_4QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_4QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_4QVal_Int_2_argbuf_r && lizzieLet13_1_4QVal_Int_2_bufchan_buf[0]))
        lizzieLet13_1_4QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_4QVal_Int_2_argbuf_r) && (! lizzieLet13_1_4QVal_Int_2_bufchan_buf[0])))
        lizzieLet13_1_4QVal_Int_2_bufchan_buf <= lizzieLet13_1_4QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet13_1_5,QTree_Int) (is_z_kronahW_goMux_mux,MyDTInt_Bool) > [(_28,MyDTInt_Bool),
                                                                                               (lizzieLet13_1_5QVal_Int,MyDTInt_Bool),
                                                                                               (lizzieLet13_1_5QNode_Int,MyDTInt_Bool),
                                                                                               (_27,MyDTInt_Bool)] */
  logic [3:0] is_z_kronahW_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_5_d[0] && is_z_kronahW_goMux_mux_d[0]))
      unique case (lizzieLet13_1_5_d[2:1])
        2'd0: is_z_kronahW_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_kronahW_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_kronahW_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_kronahW_goMux_mux_onehotd = 4'd8;
        default: is_z_kronahW_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_kronahW_goMux_mux_onehotd = 4'd0;
  assign _28_d = is_z_kronahW_goMux_mux_onehotd[0];
  assign lizzieLet13_1_5QVal_Int_d = is_z_kronahW_goMux_mux_onehotd[1];
  assign lizzieLet13_1_5QNode_Int_d = is_z_kronahW_goMux_mux_onehotd[2];
  assign _27_d = is_z_kronahW_goMux_mux_onehotd[3];
  assign is_z_kronahW_goMux_mux_r = (| (is_z_kronahW_goMux_mux_onehotd & {_27_r,
                                                                          lizzieLet13_1_5QNode_Int_r,
                                                                          lizzieLet13_1_5QVal_Int_r,
                                                                          _28_r}));
  assign lizzieLet13_1_5_r = is_z_kronahW_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet13_1_5QNode_Int,MyDTInt_Bool) > [(lizzieLet13_1_5QNode_Int_1,MyDTInt_Bool),
                                                                    (lizzieLet13_1_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet13_1_5QNode_Int_emitted;
  logic [1:0] lizzieLet13_1_5QNode_Int_done;
  assign lizzieLet13_1_5QNode_Int_1_d = (lizzieLet13_1_5QNode_Int_d[0] && (! lizzieLet13_1_5QNode_Int_emitted[0]));
  assign lizzieLet13_1_5QNode_Int_2_d = (lizzieLet13_1_5QNode_Int_d[0] && (! lizzieLet13_1_5QNode_Int_emitted[1]));
  assign lizzieLet13_1_5QNode_Int_done = (lizzieLet13_1_5QNode_Int_emitted | ({lizzieLet13_1_5QNode_Int_2_d[0],
                                                                               lizzieLet13_1_5QNode_Int_1_d[0]} & {lizzieLet13_1_5QNode_Int_2_r,
                                                                                                                   lizzieLet13_1_5QNode_Int_1_r}));
  assign lizzieLet13_1_5QNode_Int_r = (& lizzieLet13_1_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_5QNode_Int_emitted <= (lizzieLet13_1_5QNode_Int_r ? 2'd0 :
                                           lizzieLet13_1_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_1_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet13_1_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_2_bufchan_d;
  logic lizzieLet13_1_5QNode_Int_2_bufchan_r;
  assign lizzieLet13_1_5QNode_Int_2_r = ((! lizzieLet13_1_5QNode_Int_2_bufchan_d[0]) || lizzieLet13_1_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_5QNode_Int_2_r)
        lizzieLet13_1_5QNode_Int_2_bufchan_d <= lizzieLet13_1_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet13_1_5QNode_Int_2_bufchan_buf;
  assign lizzieLet13_1_5QNode_Int_2_bufchan_r = (! lizzieLet13_1_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_5QNode_Int_2_argbuf_d = (lizzieLet13_1_5QNode_Int_2_bufchan_buf[0] ? lizzieLet13_1_5QNode_Int_2_bufchan_buf :
                                                lizzieLet13_1_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_5QNode_Int_2_argbuf_r && lizzieLet13_1_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_1_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_5QNode_Int_2_argbuf_r) && (! lizzieLet13_1_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_1_5QNode_Int_2_bufchan_buf <= lizzieLet13_1_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_1_5QVal_Int,MyDTInt_Bool) > (lizzieLet13_1_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_1_5QVal_Int_bufchan_d;
  logic lizzieLet13_1_5QVal_Int_bufchan_r;
  assign lizzieLet13_1_5QVal_Int_r = ((! lizzieLet13_1_5QVal_Int_bufchan_d[0]) || lizzieLet13_1_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_5QVal_Int_r)
        lizzieLet13_1_5QVal_Int_bufchan_d <= lizzieLet13_1_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet13_1_5QVal_Int_bufchan_buf;
  assign lizzieLet13_1_5QVal_Int_bufchan_r = (! lizzieLet13_1_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_5QVal_Int_1_argbuf_d = (lizzieLet13_1_5QVal_Int_bufchan_buf[0] ? lizzieLet13_1_5QVal_Int_bufchan_buf :
                                               lizzieLet13_1_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_5QVal_Int_1_argbuf_r && lizzieLet13_1_5QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_5QVal_Int_1_argbuf_r) && (! lizzieLet13_1_5QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_5QVal_Int_bufchan_buf <= lizzieLet13_1_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet13_1_6,QTree_Int) (is_z_mapahY_goMux_mux,MyDTInt_Bool) > [(_26,MyDTInt_Bool),
                                                                                              (lizzieLet13_1_6QVal_Int,MyDTInt_Bool),
                                                                                              (lizzieLet13_1_6QNode_Int,MyDTInt_Bool),
                                                                                              (_25,MyDTInt_Bool)] */
  logic [3:0] is_z_mapahY_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_6_d[0] && is_z_mapahY_goMux_mux_d[0]))
      unique case (lizzieLet13_1_6_d[2:1])
        2'd0: is_z_mapahY_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_mapahY_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_mapahY_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_mapahY_goMux_mux_onehotd = 4'd8;
        default: is_z_mapahY_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_mapahY_goMux_mux_onehotd = 4'd0;
  assign _26_d = is_z_mapahY_goMux_mux_onehotd[0];
  assign lizzieLet13_1_6QVal_Int_d = is_z_mapahY_goMux_mux_onehotd[1];
  assign lizzieLet13_1_6QNode_Int_d = is_z_mapahY_goMux_mux_onehotd[2];
  assign _25_d = is_z_mapahY_goMux_mux_onehotd[3];
  assign is_z_mapahY_goMux_mux_r = (| (is_z_mapahY_goMux_mux_onehotd & {_25_r,
                                                                        lizzieLet13_1_6QNode_Int_r,
                                                                        lizzieLet13_1_6QVal_Int_r,
                                                                        _26_r}));
  assign lizzieLet13_1_6_r = is_z_mapahY_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet13_1_6QNode_Int,MyDTInt_Bool) > [(lizzieLet13_1_6QNode_Int_1,MyDTInt_Bool),
                                                                    (lizzieLet13_1_6QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet13_1_6QNode_Int_emitted;
  logic [1:0] lizzieLet13_1_6QNode_Int_done;
  assign lizzieLet13_1_6QNode_Int_1_d = (lizzieLet13_1_6QNode_Int_d[0] && (! lizzieLet13_1_6QNode_Int_emitted[0]));
  assign lizzieLet13_1_6QNode_Int_2_d = (lizzieLet13_1_6QNode_Int_d[0] && (! lizzieLet13_1_6QNode_Int_emitted[1]));
  assign lizzieLet13_1_6QNode_Int_done = (lizzieLet13_1_6QNode_Int_emitted | ({lizzieLet13_1_6QNode_Int_2_d[0],
                                                                               lizzieLet13_1_6QNode_Int_1_d[0]} & {lizzieLet13_1_6QNode_Int_2_r,
                                                                                                                   lizzieLet13_1_6QNode_Int_1_r}));
  assign lizzieLet13_1_6QNode_Int_r = (& lizzieLet13_1_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_6QNode_Int_emitted <= (lizzieLet13_1_6QNode_Int_r ? 2'd0 :
                                           lizzieLet13_1_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_1_6QNode_Int_2,MyDTInt_Bool) > (lizzieLet13_1_6QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_2_bufchan_d;
  logic lizzieLet13_1_6QNode_Int_2_bufchan_r;
  assign lizzieLet13_1_6QNode_Int_2_r = ((! lizzieLet13_1_6QNode_Int_2_bufchan_d[0]) || lizzieLet13_1_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_6QNode_Int_2_r)
        lizzieLet13_1_6QNode_Int_2_bufchan_d <= lizzieLet13_1_6QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet13_1_6QNode_Int_2_bufchan_buf;
  assign lizzieLet13_1_6QNode_Int_2_bufchan_r = (! lizzieLet13_1_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_6QNode_Int_2_argbuf_d = (lizzieLet13_1_6QNode_Int_2_bufchan_buf[0] ? lizzieLet13_1_6QNode_Int_2_bufchan_buf :
                                                lizzieLet13_1_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_6QNode_Int_2_argbuf_r && lizzieLet13_1_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_1_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_6QNode_Int_2_argbuf_r) && (! lizzieLet13_1_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_1_6QNode_Int_2_bufchan_buf <= lizzieLet13_1_6QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet13_1_6QVal_Int,MyDTInt_Bool) > (lizzieLet13_1_6QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet13_1_6QVal_Int_bufchan_d;
  logic lizzieLet13_1_6QVal_Int_bufchan_r;
  assign lizzieLet13_1_6QVal_Int_r = ((! lizzieLet13_1_6QVal_Int_bufchan_d[0]) || lizzieLet13_1_6QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_6QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_6QVal_Int_r)
        lizzieLet13_1_6QVal_Int_bufchan_d <= lizzieLet13_1_6QVal_Int_d;
  MyDTInt_Bool_t lizzieLet13_1_6QVal_Int_bufchan_buf;
  assign lizzieLet13_1_6QVal_Int_bufchan_r = (! lizzieLet13_1_6QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_6QVal_Int_1_argbuf_d = (lizzieLet13_1_6QVal_Int_bufchan_buf[0] ? lizzieLet13_1_6QVal_Int_bufchan_buf :
                                               lizzieLet13_1_6QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_6QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_6QVal_Int_1_argbuf_r && lizzieLet13_1_6QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_6QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_6QVal_Int_1_argbuf_r) && (! lizzieLet13_1_6QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_6QVal_Int_bufchan_buf <= lizzieLet13_1_6QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_QTree_Int) : (lizzieLet13_1_7,QTree_Int) (m2ahV_goMux_mux,Pointer_QTree_Int) > [(_24,Pointer_QTree_Int),
                                                                                                  (lizzieLet13_1_7QVal_Int,Pointer_QTree_Int),
                                                                                                  (lizzieLet13_1_7QNode_Int,Pointer_QTree_Int),
                                                                                                  (_23,Pointer_QTree_Int)] */
  logic [3:0] m2ahV_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_7_d[0] && m2ahV_goMux_mux_d[0]))
      unique case (lizzieLet13_1_7_d[2:1])
        2'd0: m2ahV_goMux_mux_onehotd = 4'd1;
        2'd1: m2ahV_goMux_mux_onehotd = 4'd2;
        2'd2: m2ahV_goMux_mux_onehotd = 4'd4;
        2'd3: m2ahV_goMux_mux_onehotd = 4'd8;
        default: m2ahV_goMux_mux_onehotd = 4'd0;
      endcase
    else m2ahV_goMux_mux_onehotd = 4'd0;
  assign _24_d = {m2ahV_goMux_mux_d[16:1],
                  m2ahV_goMux_mux_onehotd[0]};
  assign lizzieLet13_1_7QVal_Int_d = {m2ahV_goMux_mux_d[16:1],
                                      m2ahV_goMux_mux_onehotd[1]};
  assign lizzieLet13_1_7QNode_Int_d = {m2ahV_goMux_mux_d[16:1],
                                       m2ahV_goMux_mux_onehotd[2]};
  assign _23_d = {m2ahV_goMux_mux_d[16:1],
                  m2ahV_goMux_mux_onehotd[3]};
  assign m2ahV_goMux_mux_r = (| (m2ahV_goMux_mux_onehotd & {_23_r,
                                                            lizzieLet13_1_7QNode_Int_r,
                                                            lizzieLet13_1_7QVal_Int_r,
                                                            _24_r}));
  assign lizzieLet13_1_7_r = m2ahV_goMux_mux_r;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet13_1_7QNode_Int,Pointer_QTree_Int) > [(lizzieLet13_1_7QNode_Int_1,Pointer_QTree_Int),
                                                                              (lizzieLet13_1_7QNode_Int_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet13_1_7QNode_Int_emitted;
  logic [1:0] lizzieLet13_1_7QNode_Int_done;
  assign lizzieLet13_1_7QNode_Int_1_d = {lizzieLet13_1_7QNode_Int_d[16:1],
                                         (lizzieLet13_1_7QNode_Int_d[0] && (! lizzieLet13_1_7QNode_Int_emitted[0]))};
  assign lizzieLet13_1_7QNode_Int_2_d = {lizzieLet13_1_7QNode_Int_d[16:1],
                                         (lizzieLet13_1_7QNode_Int_d[0] && (! lizzieLet13_1_7QNode_Int_emitted[1]))};
  assign lizzieLet13_1_7QNode_Int_done = (lizzieLet13_1_7QNode_Int_emitted | ({lizzieLet13_1_7QNode_Int_2_d[0],
                                                                               lizzieLet13_1_7QNode_Int_1_d[0]} & {lizzieLet13_1_7QNode_Int_2_r,
                                                                                                                   lizzieLet13_1_7QNode_Int_1_r}));
  assign lizzieLet13_1_7QNode_Int_r = (& lizzieLet13_1_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_7QNode_Int_emitted <= (lizzieLet13_1_7QNode_Int_r ? 2'd0 :
                                           lizzieLet13_1_7QNode_Int_done);
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_1_7QNode_Int_2,Pointer_QTree_Int) > (lizzieLet13_1_7QNode_Int_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_2_bufchan_d;
  logic lizzieLet13_1_7QNode_Int_2_bufchan_r;
  assign lizzieLet13_1_7QNode_Int_2_r = ((! lizzieLet13_1_7QNode_Int_2_bufchan_d[0]) || lizzieLet13_1_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_7QNode_Int_2_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_1_7QNode_Int_2_r)
        lizzieLet13_1_7QNode_Int_2_bufchan_d <= lizzieLet13_1_7QNode_Int_2_d;
  Pointer_QTree_Int_t lizzieLet13_1_7QNode_Int_2_bufchan_buf;
  assign lizzieLet13_1_7QNode_Int_2_bufchan_r = (! lizzieLet13_1_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_7QNode_Int_2_argbuf_d = (lizzieLet13_1_7QNode_Int_2_bufchan_buf[0] ? lizzieLet13_1_7QNode_Int_2_bufchan_buf :
                                                lizzieLet13_1_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_7QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_7QNode_Int_2_argbuf_r && lizzieLet13_1_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_1_7QNode_Int_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_7QNode_Int_2_argbuf_r) && (! lizzieLet13_1_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_1_7QNode_Int_2_bufchan_buf <= lizzieLet13_1_7QNode_Int_2_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet13_1_7QVal_Int,Pointer_QTree_Int) > (lizzieLet13_1_7QVal_Int_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet13_1_7QVal_Int_bufchan_d;
  logic lizzieLet13_1_7QVal_Int_bufchan_r;
  assign lizzieLet13_1_7QVal_Int_r = ((! lizzieLet13_1_7QVal_Int_bufchan_d[0]) || lizzieLet13_1_7QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_7QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_1_7QVal_Int_r)
        lizzieLet13_1_7QVal_Int_bufchan_d <= lizzieLet13_1_7QVal_Int_d;
  Pointer_QTree_Int_t lizzieLet13_1_7QVal_Int_bufchan_buf;
  assign lizzieLet13_1_7QVal_Int_bufchan_r = (! lizzieLet13_1_7QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_7QVal_Int_1_argbuf_d = (lizzieLet13_1_7QVal_Int_bufchan_buf[0] ? lizzieLet13_1_7QVal_Int_bufchan_buf :
                                               lizzieLet13_1_7QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_7QVal_Int_1_argbuf_r && lizzieLet13_1_7QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_7QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_7QVal_Int_1_argbuf_r) && (! lizzieLet13_1_7QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_7QVal_Int_bufchan_buf <= lizzieLet13_1_7QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet13_1_8,QTree_Int) (op_kronahX_goMux_mux,MyDTInt_Int_Int) > [(_22,MyDTInt_Int_Int),
                                                                                                   (lizzieLet13_1_8QVal_Int,MyDTInt_Int_Int),
                                                                                                   (lizzieLet13_1_8QNode_Int,MyDTInt_Int_Int),
                                                                                                   (_21,MyDTInt_Int_Int)] */
  logic [3:0] op_kronahX_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_8_d[0] && op_kronahX_goMux_mux_d[0]))
      unique case (lizzieLet13_1_8_d[2:1])
        2'd0: op_kronahX_goMux_mux_onehotd = 4'd1;
        2'd1: op_kronahX_goMux_mux_onehotd = 4'd2;
        2'd2: op_kronahX_goMux_mux_onehotd = 4'd4;
        2'd3: op_kronahX_goMux_mux_onehotd = 4'd8;
        default: op_kronahX_goMux_mux_onehotd = 4'd0;
      endcase
    else op_kronahX_goMux_mux_onehotd = 4'd0;
  assign _22_d = op_kronahX_goMux_mux_onehotd[0];
  assign lizzieLet13_1_8QVal_Int_d = op_kronahX_goMux_mux_onehotd[1];
  assign lizzieLet13_1_8QNode_Int_d = op_kronahX_goMux_mux_onehotd[2];
  assign _21_d = op_kronahX_goMux_mux_onehotd[3];
  assign op_kronahX_goMux_mux_r = (| (op_kronahX_goMux_mux_onehotd & {_21_r,
                                                                      lizzieLet13_1_8QNode_Int_r,
                                                                      lizzieLet13_1_8QVal_Int_r,
                                                                      _22_r}));
  assign lizzieLet13_1_8_r = op_kronahX_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet13_1_8QNode_Int,MyDTInt_Int_Int) > [(lizzieLet13_1_8QNode_Int_1,MyDTInt_Int_Int),
                                                                          (lizzieLet13_1_8QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet13_1_8QNode_Int_emitted;
  logic [1:0] lizzieLet13_1_8QNode_Int_done;
  assign lizzieLet13_1_8QNode_Int_1_d = (lizzieLet13_1_8QNode_Int_d[0] && (! lizzieLet13_1_8QNode_Int_emitted[0]));
  assign lizzieLet13_1_8QNode_Int_2_d = (lizzieLet13_1_8QNode_Int_d[0] && (! lizzieLet13_1_8QNode_Int_emitted[1]));
  assign lizzieLet13_1_8QNode_Int_done = (lizzieLet13_1_8QNode_Int_emitted | ({lizzieLet13_1_8QNode_Int_2_d[0],
                                                                               lizzieLet13_1_8QNode_Int_1_d[0]} & {lizzieLet13_1_8QNode_Int_2_r,
                                                                                                                   lizzieLet13_1_8QNode_Int_1_r}));
  assign lizzieLet13_1_8QNode_Int_r = (& lizzieLet13_1_8QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_8QNode_Int_emitted <= 2'd0;
    else
      lizzieLet13_1_8QNode_Int_emitted <= (lizzieLet13_1_8QNode_Int_r ? 2'd0 :
                                           lizzieLet13_1_8QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet13_1_8QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet13_1_8QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_2_bufchan_d;
  logic lizzieLet13_1_8QNode_Int_2_bufchan_r;
  assign lizzieLet13_1_8QNode_Int_2_r = ((! lizzieLet13_1_8QNode_Int_2_bufchan_d[0]) || lizzieLet13_1_8QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_8QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_8QNode_Int_2_r)
        lizzieLet13_1_8QNode_Int_2_bufchan_d <= lizzieLet13_1_8QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet13_1_8QNode_Int_2_bufchan_buf;
  assign lizzieLet13_1_8QNode_Int_2_bufchan_r = (! lizzieLet13_1_8QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet13_1_8QNode_Int_2_argbuf_d = (lizzieLet13_1_8QNode_Int_2_bufchan_buf[0] ? lizzieLet13_1_8QNode_Int_2_bufchan_buf :
                                                lizzieLet13_1_8QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_8QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_8QNode_Int_2_argbuf_r && lizzieLet13_1_8QNode_Int_2_bufchan_buf[0]))
        lizzieLet13_1_8QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_8QNode_Int_2_argbuf_r) && (! lizzieLet13_1_8QNode_Int_2_bufchan_buf[0])))
        lizzieLet13_1_8QNode_Int_2_bufchan_buf <= lizzieLet13_1_8QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet13_1_8QVal_Int,MyDTInt_Int_Int) > (lizzieLet13_1_8QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet13_1_8QVal_Int_bufchan_d;
  logic lizzieLet13_1_8QVal_Int_bufchan_r;
  assign lizzieLet13_1_8QVal_Int_r = ((! lizzieLet13_1_8QVal_Int_bufchan_d[0]) || lizzieLet13_1_8QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_8QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet13_1_8QVal_Int_r)
        lizzieLet13_1_8QVal_Int_bufchan_d <= lizzieLet13_1_8QVal_Int_d;
  MyDTInt_Int_Int_t lizzieLet13_1_8QVal_Int_bufchan_buf;
  assign lizzieLet13_1_8QVal_Int_bufchan_r = (! lizzieLet13_1_8QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_8QVal_Int_1_argbuf_d = (lizzieLet13_1_8QVal_Int_bufchan_buf[0] ? lizzieLet13_1_8QVal_Int_bufchan_buf :
                                               lizzieLet13_1_8QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet13_1_8QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet13_1_8QVal_Int_1_argbuf_r && lizzieLet13_1_8QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_8QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet13_1_8QVal_Int_1_argbuf_r) && (! lizzieLet13_1_8QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_8QVal_Int_bufchan_buf <= lizzieLet13_1_8QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf_f_Int_Int_Int_Int) : (lizzieLet13_1_9,QTree_Int) (sc_0_2_goMux_mux,Pointer_CTf_f_Int_Int_Int_Int) > [(lizzieLet13_1_9QNone_Int,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                           (lizzieLet13_1_9QVal_Int,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                           (lizzieLet13_1_9QNode_Int,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                           (lizzieLet13_1_9QError_Int,Pointer_CTf_f_Int_Int_Int_Int)] */
  logic [3:0] sc_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet13_1_9_d[0] && sc_0_2_goMux_mux_d[0]))
      unique case (lizzieLet13_1_9_d[2:1])
        2'd0: sc_0_2_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_2_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_2_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_2_goMux_mux_onehotd = 4'd8;
        default: sc_0_2_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_2_goMux_mux_onehotd = 4'd0;
  assign lizzieLet13_1_9QNone_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                       sc_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet13_1_9QVal_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                      sc_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet13_1_9QNode_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                       sc_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet13_1_9QError_Int_d = {sc_0_2_goMux_mux_d[16:1],
                                        sc_0_2_goMux_mux_onehotd[3]};
  assign sc_0_2_goMux_mux_r = (| (sc_0_2_goMux_mux_onehotd & {lizzieLet13_1_9QError_Int_r,
                                                              lizzieLet13_1_9QNode_Int_r,
                                                              lizzieLet13_1_9QVal_Int_r,
                                                              lizzieLet13_1_9QNone_Int_r}));
  assign lizzieLet13_1_9_r = sc_0_2_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (lizzieLet13_1_9QError_Int,Pointer_CTf_f_Int_Int_Int_Int) > (lizzieLet13_1_9QError_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QError_Int_bufchan_d;
  logic lizzieLet13_1_9QError_Int_bufchan_r;
  assign lizzieLet13_1_9QError_Int_r = ((! lizzieLet13_1_9QError_Int_bufchan_d[0]) || lizzieLet13_1_9QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_1_9QError_Int_r)
        lizzieLet13_1_9QError_Int_bufchan_d <= lizzieLet13_1_9QError_Int_d;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QError_Int_bufchan_buf;
  assign lizzieLet13_1_9QError_Int_bufchan_r = (! lizzieLet13_1_9QError_Int_bufchan_buf[0]);
  assign lizzieLet13_1_9QError_Int_1_argbuf_d = (lizzieLet13_1_9QError_Int_bufchan_buf[0] ? lizzieLet13_1_9QError_Int_bufchan_buf :
                                                 lizzieLet13_1_9QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_9QError_Int_1_argbuf_r && lizzieLet13_1_9QError_Int_bufchan_buf[0]))
        lizzieLet13_1_9QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_9QError_Int_1_argbuf_r) && (! lizzieLet13_1_9QError_Int_bufchan_buf[0])))
        lizzieLet13_1_9QError_Int_bufchan_buf <= lizzieLet13_1_9QError_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int_Int_Int,
      Dcon Lcall_f_f_Int_Int_Int_Int3) : [(lizzieLet13_1_9QNode_Int,Pointer_CTf_f_Int_Int_Int_Int),
                                          (q1ai1_destruct,Pointer_QTree_Int),
                                          (lizzieLet13_1_7QNode_Int_1,Pointer_QTree_Int),
                                          (lizzieLet13_1_5QNode_Int_1,MyDTInt_Bool),
                                          (lizzieLet13_1_8QNode_Int_1,MyDTInt_Int_Int),
                                          (lizzieLet13_1_6QNode_Int_1,MyDTInt_Bool),
                                          (lizzieLet13_1_3QNode_Int_1,MyDTInt_Int),
                                          (q2ai2_destruct,Pointer_QTree_Int),
                                          (q3ai3_destruct,Pointer_QTree_Int)] > (lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3,CTf_f_Int_Int_Int_Int) */
  assign lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_d = Lcall_f_f_Int_Int_Int_Int3_dc((& {lizzieLet13_1_9QNode_Int_d[0],
                                                                                                                                                                                                                                                           q1ai1_destruct_d[0],
                                                                                                                                                                                                                                                           lizzieLet13_1_7QNode_Int_1_d[0],
                                                                                                                                                                                                                                                           lizzieLet13_1_5QNode_Int_1_d[0],
                                                                                                                                                                                                                                                           lizzieLet13_1_8QNode_Int_1_d[0],
                                                                                                                                                                                                                                                           lizzieLet13_1_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                           lizzieLet13_1_3QNode_Int_1_d[0],
                                                                                                                                                                                                                                                           q2ai2_destruct_d[0],
                                                                                                                                                                                                                                                           q3ai3_destruct_d[0]}), lizzieLet13_1_9QNode_Int_d, q1ai1_destruct_d, lizzieLet13_1_7QNode_Int_1_d, lizzieLet13_1_5QNode_Int_1_d, lizzieLet13_1_8QNode_Int_1_d, lizzieLet13_1_6QNode_Int_1_d, lizzieLet13_1_3QNode_Int_1_d, q2ai2_destruct_d, q3ai3_destruct_d);
  assign {lizzieLet13_1_9QNode_Int_r,
          q1ai1_destruct_r,
          lizzieLet13_1_7QNode_Int_1_r,
          lizzieLet13_1_5QNode_Int_1_r,
          lizzieLet13_1_8QNode_Int_1_r,
          lizzieLet13_1_6QNode_Int_1_r,
          lizzieLet13_1_3QNode_Int_1_r,
          q2ai2_destruct_r,
          q3ai3_destruct_r} = {9 {(lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_r && lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3,CTf_f_Int_Int_Int_Int) > (lizzieLet15_1_argbuf,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d;
  logic lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_r;
  assign lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_r = ((! lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d[0]) || lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d <= {83'd0,
                                                                                                                                                                                                                                1'd0};
    else
      if (lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_r)
        lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d <= lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_d;
  CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf;
  assign lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_r = (! lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet15_1_argbuf_d = (lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0] ? lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf :
                                   lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                                                                                  1'd0};
    else
      if ((lizzieLet15_1_argbuf_r && lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= {83'd0,
                                                                                                                                                                                                                                    1'd0};
      else if (((! lizzieLet15_1_argbuf_r) && (! lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= lizzieLet13_1_9QNode_Int_1q1ai1_1lizzieLet13_1_7QNode_Int_1lizzieLet13_1_5QNode_Int_1lizzieLet13_1_8QNode_Int_1lizzieLet13_1_6QNode_Int_1lizzieLet13_1_3QNode_Int_1q2ai2_1q3ai3_1Lcall_f_f_Int_Int_Int_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (lizzieLet13_1_9QNone_Int,Pointer_CTf_f_Int_Int_Int_Int) > (lizzieLet13_1_9QNone_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNone_Int_bufchan_d;
  logic lizzieLet13_1_9QNone_Int_bufchan_r;
  assign lizzieLet13_1_9QNone_Int_r = ((! lizzieLet13_1_9QNone_Int_bufchan_d[0]) || lizzieLet13_1_9QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_1_9QNone_Int_r)
        lizzieLet13_1_9QNone_Int_bufchan_d <= lizzieLet13_1_9QNone_Int_d;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QNone_Int_bufchan_buf;
  assign lizzieLet13_1_9QNone_Int_bufchan_r = (! lizzieLet13_1_9QNone_Int_bufchan_buf[0]);
  assign lizzieLet13_1_9QNone_Int_1_argbuf_d = (lizzieLet13_1_9QNone_Int_bufchan_buf[0] ? lizzieLet13_1_9QNone_Int_bufchan_buf :
                                                lizzieLet13_1_9QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_9QNone_Int_1_argbuf_r && lizzieLet13_1_9QNone_Int_bufchan_buf[0]))
        lizzieLet13_1_9QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_9QNone_Int_1_argbuf_r) && (! lizzieLet13_1_9QNone_Int_bufchan_buf[0])))
        lizzieLet13_1_9QNone_Int_bufchan_buf <= lizzieLet13_1_9QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (lizzieLet13_1_9QVal_Int,Pointer_CTf_f_Int_Int_Int_Int) > (lizzieLet13_1_9QVal_Int_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QVal_Int_bufchan_d;
  logic lizzieLet13_1_9QVal_Int_bufchan_r;
  assign lizzieLet13_1_9QVal_Int_r = ((! lizzieLet13_1_9QVal_Int_bufchan_d[0]) || lizzieLet13_1_9QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet13_1_9QVal_Int_r)
        lizzieLet13_1_9QVal_Int_bufchan_d <= lizzieLet13_1_9QVal_Int_d;
  Pointer_CTf_f_Int_Int_Int_Int_t lizzieLet13_1_9QVal_Int_bufchan_buf;
  assign lizzieLet13_1_9QVal_Int_bufchan_r = (! lizzieLet13_1_9QVal_Int_bufchan_buf[0]);
  assign lizzieLet13_1_9QVal_Int_1_argbuf_d = (lizzieLet13_1_9QVal_Int_bufchan_buf[0] ? lizzieLet13_1_9QVal_Int_bufchan_buf :
                                               lizzieLet13_1_9QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet13_1_9QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet13_1_9QVal_Int_1_argbuf_r && lizzieLet13_1_9QVal_Int_bufchan_buf[0]))
        lizzieLet13_1_9QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet13_1_9QVal_Int_1_argbuf_r) && (! lizzieLet13_1_9QVal_Int_bufchan_buf[0])))
        lizzieLet13_1_9QVal_Int_bufchan_buf <= lizzieLet13_1_9QVal_Int_bufchan_d;
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int0) : (lizzieLet19_1Lcall_$wnnz_Int0,CT$wnnz_Int) > [(wwstK_4_destruct,Int#),
                                                                                  (ww1XuL_2_destruct,Int#),
                                                                                  (ww2XuO_1_destruct,Int#),
                                                                                  (sc_0_6_destruct,Pointer_CT$wnnz_Int)] */
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int0_emitted;
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int0_done;
  assign wwstK_4_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int0_d[35:4],
                               (lizzieLet19_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int0_emitted[0]))};
  assign ww1XuL_2_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int0_d[67:36],
                                (lizzieLet19_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int0_emitted[1]))};
  assign ww2XuO_1_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int0_d[99:68],
                                (lizzieLet19_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int0_emitted[2]))};
  assign sc_0_6_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int0_d[115:100],
                              (lizzieLet19_1Lcall_$wnnz_Int0_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int0_emitted[3]))};
  assign lizzieLet19_1Lcall_$wnnz_Int0_done = (lizzieLet19_1Lcall_$wnnz_Int0_emitted | ({sc_0_6_destruct_d[0],
                                                                                         ww2XuO_1_destruct_d[0],
                                                                                         ww1XuL_2_destruct_d[0],
                                                                                         wwstK_4_destruct_d[0]} & {sc_0_6_destruct_r,
                                                                                                                   ww2XuO_1_destruct_r,
                                                                                                                   ww1XuL_2_destruct_r,
                                                                                                                   wwstK_4_destruct_r}));
  assign lizzieLet19_1Lcall_$wnnz_Int0_r = (& lizzieLet19_1Lcall_$wnnz_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1Lcall_$wnnz_Int0_emitted <= 4'd0;
    else
      lizzieLet19_1Lcall_$wnnz_Int0_emitted <= (lizzieLet19_1Lcall_$wnnz_Int0_r ? 4'd0 :
                                                lizzieLet19_1Lcall_$wnnz_Int0_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int1) : (lizzieLet19_1Lcall_$wnnz_Int1,CT$wnnz_Int) > [(wwstK_3_destruct,Int#),
                                                                                  (ww1XuL_1_destruct,Int#),
                                                                                  (sc_0_5_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4abZ_3_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int1_emitted;
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int1_done;
  assign wwstK_3_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int1_d[35:4],
                               (lizzieLet19_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int1_emitted[0]))};
  assign ww1XuL_1_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int1_d[67:36],
                                (lizzieLet19_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int1_emitted[1]))};
  assign sc_0_5_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int1_d[83:68],
                              (lizzieLet19_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int1_emitted[2]))};
  assign q4abZ_3_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int1_d[99:84],
                               (lizzieLet19_1Lcall_$wnnz_Int1_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int1_emitted[3]))};
  assign lizzieLet19_1Lcall_$wnnz_Int1_done = (lizzieLet19_1Lcall_$wnnz_Int1_emitted | ({q4abZ_3_destruct_d[0],
                                                                                         sc_0_5_destruct_d[0],
                                                                                         ww1XuL_1_destruct_d[0],
                                                                                         wwstK_3_destruct_d[0]} & {q4abZ_3_destruct_r,
                                                                                                                   sc_0_5_destruct_r,
                                                                                                                   ww1XuL_1_destruct_r,
                                                                                                                   wwstK_3_destruct_r}));
  assign lizzieLet19_1Lcall_$wnnz_Int1_r = (& lizzieLet19_1Lcall_$wnnz_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1Lcall_$wnnz_Int1_emitted <= 4'd0;
    else
      lizzieLet19_1Lcall_$wnnz_Int1_emitted <= (lizzieLet19_1Lcall_$wnnz_Int1_r ? 4'd0 :
                                                lizzieLet19_1Lcall_$wnnz_Int1_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int2) : (lizzieLet19_1Lcall_$wnnz_Int2,CT$wnnz_Int) > [(wwstK_2_destruct,Int#),
                                                                                  (sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4abZ_2_destruct,Pointer_QTree_Int),
                                                                                  (q3abY_2_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int2_emitted;
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int2_done;
  assign wwstK_2_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int2_d[35:4],
                               (lizzieLet19_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int2_emitted[0]))};
  assign sc_0_4_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int2_d[51:36],
                              (lizzieLet19_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int2_emitted[1]))};
  assign q4abZ_2_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int2_d[67:52],
                               (lizzieLet19_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int2_emitted[2]))};
  assign q3abY_2_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int2_d[83:68],
                               (lizzieLet19_1Lcall_$wnnz_Int2_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int2_emitted[3]))};
  assign lizzieLet19_1Lcall_$wnnz_Int2_done = (lizzieLet19_1Lcall_$wnnz_Int2_emitted | ({q3abY_2_destruct_d[0],
                                                                                         q4abZ_2_destruct_d[0],
                                                                                         sc_0_4_destruct_d[0],
                                                                                         wwstK_2_destruct_d[0]} & {q3abY_2_destruct_r,
                                                                                                                   q4abZ_2_destruct_r,
                                                                                                                   sc_0_4_destruct_r,
                                                                                                                   wwstK_2_destruct_r}));
  assign lizzieLet19_1Lcall_$wnnz_Int2_r = (& lizzieLet19_1Lcall_$wnnz_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1Lcall_$wnnz_Int2_emitted <= 4'd0;
    else
      lizzieLet19_1Lcall_$wnnz_Int2_emitted <= (lizzieLet19_1Lcall_$wnnz_Int2_r ? 4'd0 :
                                                lizzieLet19_1Lcall_$wnnz_Int2_done);
  
  /* destruct (Ty CT$wnnz_Int,
          Dcon Lcall_$wnnz_Int3) : (lizzieLet19_1Lcall_$wnnz_Int3,CT$wnnz_Int) > [(sc_0_3_destruct,Pointer_CT$wnnz_Int),
                                                                                  (q4abZ_1_destruct,Pointer_QTree_Int),
                                                                                  (q3abY_1_destruct,Pointer_QTree_Int),
                                                                                  (q2abX_1_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int3_emitted;
  logic [3:0] lizzieLet19_1Lcall_$wnnz_Int3_done;
  assign sc_0_3_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int3_d[19:4],
                              (lizzieLet19_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int3_emitted[0]))};
  assign q4abZ_1_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int3_d[35:20],
                               (lizzieLet19_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int3_emitted[1]))};
  assign q3abY_1_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int3_d[51:36],
                               (lizzieLet19_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int3_emitted[2]))};
  assign q2abX_1_destruct_d = {lizzieLet19_1Lcall_$wnnz_Int3_d[67:52],
                               (lizzieLet19_1Lcall_$wnnz_Int3_d[0] && (! lizzieLet19_1Lcall_$wnnz_Int3_emitted[3]))};
  assign lizzieLet19_1Lcall_$wnnz_Int3_done = (lizzieLet19_1Lcall_$wnnz_Int3_emitted | ({q2abX_1_destruct_d[0],
                                                                                         q3abY_1_destruct_d[0],
                                                                                         q4abZ_1_destruct_d[0],
                                                                                         sc_0_3_destruct_d[0]} & {q2abX_1_destruct_r,
                                                                                                                  q3abY_1_destruct_r,
                                                                                                                  q4abZ_1_destruct_r,
                                                                                                                  sc_0_3_destruct_r}));
  assign lizzieLet19_1Lcall_$wnnz_Int3_r = (& lizzieLet19_1Lcall_$wnnz_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_1Lcall_$wnnz_Int3_emitted <= 4'd0;
    else
      lizzieLet19_1Lcall_$wnnz_Int3_emitted <= (lizzieLet19_1Lcall_$wnnz_Int3_r ? 4'd0 :
                                                lizzieLet19_1Lcall_$wnnz_Int3_done);
  
  /* demux (Ty CT$wnnz_Int,
       Ty CT$wnnz_Int) : (lizzieLet19_2,CT$wnnz_Int) (lizzieLet19_1,CT$wnnz_Int) > [(_20,CT$wnnz_Int),
                                                                                    (lizzieLet19_1Lcall_$wnnz_Int3,CT$wnnz_Int),
                                                                                    (lizzieLet19_1Lcall_$wnnz_Int2,CT$wnnz_Int),
                                                                                    (lizzieLet19_1Lcall_$wnnz_Int1,CT$wnnz_Int),
                                                                                    (lizzieLet19_1Lcall_$wnnz_Int0,CT$wnnz_Int)] */
  logic [4:0] lizzieLet19_1_onehotd;
  always_comb
    if ((lizzieLet19_2_d[0] && lizzieLet19_1_d[0]))
      unique case (lizzieLet19_2_d[3:1])
        3'd0: lizzieLet19_1_onehotd = 5'd1;
        3'd1: lizzieLet19_1_onehotd = 5'd2;
        3'd2: lizzieLet19_1_onehotd = 5'd4;
        3'd3: lizzieLet19_1_onehotd = 5'd8;
        3'd4: lizzieLet19_1_onehotd = 5'd16;
        default: lizzieLet19_1_onehotd = 5'd0;
      endcase
    else lizzieLet19_1_onehotd = 5'd0;
  assign _20_d = {lizzieLet19_1_d[115:1], lizzieLet19_1_onehotd[0]};
  assign lizzieLet19_1Lcall_$wnnz_Int3_d = {lizzieLet19_1_d[115:1],
                                            lizzieLet19_1_onehotd[1]};
  assign lizzieLet19_1Lcall_$wnnz_Int2_d = {lizzieLet19_1_d[115:1],
                                            lizzieLet19_1_onehotd[2]};
  assign lizzieLet19_1Lcall_$wnnz_Int1_d = {lizzieLet19_1_d[115:1],
                                            lizzieLet19_1_onehotd[3]};
  assign lizzieLet19_1Lcall_$wnnz_Int0_d = {lizzieLet19_1_d[115:1],
                                            lizzieLet19_1_onehotd[4]};
  assign lizzieLet19_1_r = (| (lizzieLet19_1_onehotd & {lizzieLet19_1Lcall_$wnnz_Int0_r,
                                                        lizzieLet19_1Lcall_$wnnz_Int1_r,
                                                        lizzieLet19_1Lcall_$wnnz_Int2_r,
                                                        lizzieLet19_1Lcall_$wnnz_Int3_r,
                                                        _20_r}));
  assign lizzieLet19_2_r = lizzieLet19_1_r;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Go) : (lizzieLet19_3,CT$wnnz_Int) (go_15_goMux_data,Go) > [(_19,Go),
                                                                     (lizzieLet19_3Lcall_$wnnz_Int3,Go),
                                                                     (lizzieLet19_3Lcall_$wnnz_Int2,Go),
                                                                     (lizzieLet19_3Lcall_$wnnz_Int1,Go),
                                                                     (lizzieLet19_3Lcall_$wnnz_Int0,Go)] */
  logic [4:0] go_15_goMux_data_onehotd;
  always_comb
    if ((lizzieLet19_3_d[0] && go_15_goMux_data_d[0]))
      unique case (lizzieLet19_3_d[3:1])
        3'd0: go_15_goMux_data_onehotd = 5'd1;
        3'd1: go_15_goMux_data_onehotd = 5'd2;
        3'd2: go_15_goMux_data_onehotd = 5'd4;
        3'd3: go_15_goMux_data_onehotd = 5'd8;
        3'd4: go_15_goMux_data_onehotd = 5'd16;
        default: go_15_goMux_data_onehotd = 5'd0;
      endcase
    else go_15_goMux_data_onehotd = 5'd0;
  assign _19_d = go_15_goMux_data_onehotd[0];
  assign lizzieLet19_3Lcall_$wnnz_Int3_d = go_15_goMux_data_onehotd[1];
  assign lizzieLet19_3Lcall_$wnnz_Int2_d = go_15_goMux_data_onehotd[2];
  assign lizzieLet19_3Lcall_$wnnz_Int1_d = go_15_goMux_data_onehotd[3];
  assign lizzieLet19_3Lcall_$wnnz_Int0_d = go_15_goMux_data_onehotd[4];
  assign go_15_goMux_data_r = (| (go_15_goMux_data_onehotd & {lizzieLet19_3Lcall_$wnnz_Int0_r,
                                                              lizzieLet19_3Lcall_$wnnz_Int1_r,
                                                              lizzieLet19_3Lcall_$wnnz_Int2_r,
                                                              lizzieLet19_3Lcall_$wnnz_Int3_r,
                                                              _19_r}));
  assign lizzieLet19_3_r = go_15_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wnnz_Int0,Go) > (lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d;
  logic lizzieLet19_3Lcall_$wnnz_Int0_bufchan_r;
  assign lizzieLet19_3Lcall_$wnnz_Int0_r = ((! lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d[0]) || lizzieLet19_3Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wnnz_Int0_r)
        lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d <= lizzieLet19_3Lcall_$wnnz_Int0_d;
  Go_t lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf;
  assign lizzieLet19_3Lcall_$wnnz_Int0_bufchan_r = (! lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_d = (lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf[0] ? lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf :
                                                     lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_r && lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_r) && (! lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wnnz_Int0_bufchan_buf <= lizzieLet19_3Lcall_$wnnz_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wnnz_Int1,Go) > (lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d;
  logic lizzieLet19_3Lcall_$wnnz_Int1_bufchan_r;
  assign lizzieLet19_3Lcall_$wnnz_Int1_r = ((! lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d[0]) || lizzieLet19_3Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wnnz_Int1_r)
        lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d <= lizzieLet19_3Lcall_$wnnz_Int1_d;
  Go_t lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf;
  assign lizzieLet19_3Lcall_$wnnz_Int1_bufchan_r = (! lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_d = (lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf[0] ? lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf :
                                                     lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_r && lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wnnz_Int1_1_argbuf_r) && (! lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wnnz_Int1_bufchan_buf <= lizzieLet19_3Lcall_$wnnz_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wnnz_Int2,Go) > (lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet19_3Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet19_3Lcall_$wnnz_Int2_r = ((! lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet19_3Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wnnz_Int2_r)
        lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d <= lizzieLet19_3Lcall_$wnnz_Int2_d;
  Go_t lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet19_3Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_d = (lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf :
                                                     lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_r && lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wnnz_Int2_1_argbuf_r) && (! lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet19_3Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet19_3Lcall_$wnnz_Int3,Go) > (lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf,Go) */
  Go_t lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet19_3Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet19_3Lcall_$wnnz_Int3_r = ((! lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet19_3Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet19_3Lcall_$wnnz_Int3_r)
        lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d <= lizzieLet19_3Lcall_$wnnz_Int3_d;
  Go_t lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet19_3Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_d = (lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf :
                                                     lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_r && lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet19_3Lcall_$wnnz_Int3_1_argbuf_r) && (! lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet19_3Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet19_3Lcall_$wnnz_Int3_bufchan_d;
  
  /* demux (Ty CT$wnnz_Int,
       Ty Int#) : (lizzieLet19_4,CT$wnnz_Int) (srtarg_0_goMux_mux,Int#) > [(lizzieLet19_4L$wnnz_Intsbos,Int#),
                                                                           (lizzieLet19_4Lcall_$wnnz_Int3,Int#),
                                                                           (lizzieLet19_4Lcall_$wnnz_Int2,Int#),
                                                                           (lizzieLet19_4Lcall_$wnnz_Int1,Int#),
                                                                           (lizzieLet19_4Lcall_$wnnz_Int0,Int#)] */
  logic [4:0] srtarg_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet19_4_d[0] && srtarg_0_goMux_mux_d[0]))
      unique case (lizzieLet19_4_d[3:1])
        3'd0: srtarg_0_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_goMux_mux_onehotd = 5'd0;
  assign lizzieLet19_4L$wnnz_Intsbos_d = {srtarg_0_goMux_mux_d[32:1],
                                          srtarg_0_goMux_mux_onehotd[0]};
  assign lizzieLet19_4Lcall_$wnnz_Int3_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[1]};
  assign lizzieLet19_4Lcall_$wnnz_Int2_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[2]};
  assign lizzieLet19_4Lcall_$wnnz_Int1_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[3]};
  assign lizzieLet19_4Lcall_$wnnz_Int0_d = {srtarg_0_goMux_mux_d[32:1],
                                            srtarg_0_goMux_mux_onehotd[4]};
  assign srtarg_0_goMux_mux_r = (| (srtarg_0_goMux_mux_onehotd & {lizzieLet19_4Lcall_$wnnz_Int0_r,
                                                                  lizzieLet19_4Lcall_$wnnz_Int1_r,
                                                                  lizzieLet19_4Lcall_$wnnz_Int2_r,
                                                                  lizzieLet19_4Lcall_$wnnz_Int3_r,
                                                                  lizzieLet19_4L$wnnz_Intsbos_r}));
  assign lizzieLet19_4_r = srtarg_0_goMux_mux_r;
  
  /* fork (Ty Int#) : (lizzieLet19_4L$wnnz_Intsbos,Int#) > [(lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#),
                                                       (lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#)] */
  logic [1:0] lizzieLet19_4L$wnnz_Intsbos_emitted;
  logic [1:0] lizzieLet19_4L$wnnz_Intsbos_done;
  assign lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_d = {lizzieLet19_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet19_4L$wnnz_Intsbos_d[0] && (! lizzieLet19_4L$wnnz_Intsbos_emitted[0]))};
  assign lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_d = {lizzieLet19_4L$wnnz_Intsbos_d[32:1],
                                                               (lizzieLet19_4L$wnnz_Intsbos_d[0] && (! lizzieLet19_4L$wnnz_Intsbos_emitted[1]))};
  assign lizzieLet19_4L$wnnz_Intsbos_done = (lizzieLet19_4L$wnnz_Intsbos_emitted | ({lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                     lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                               lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet19_4L$wnnz_Intsbos_r = (& lizzieLet19_4L$wnnz_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet19_4L$wnnz_Intsbos_emitted <= 2'd0;
    else
      lizzieLet19_4L$wnnz_Intsbos_emitted <= (lizzieLet19_4L$wnnz_Intsbos_r ? 2'd0 :
                                              lizzieLet19_4L$wnnz_Intsbos_done);
  
  /* togo (Ty Int#) : (lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1,Int#) > (call_$wnnz_Int_goConst,Go) */
  assign call_$wnnz_Int_goConst_d = lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_1_r = call_$wnnz_Int_goConst_r;
  
  /* buf (Ty Int#) : (lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2,Int#) > ($wnnz_Int_resbuf,Int#) */
  \Int#_t  lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= {32'd0,
                                                                     1'd0};
    else
      if (lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_d;
  \Int#_t  lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign \$wnnz_Int_resbuf_d  = (lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                 lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                       1'd0};
    else
      if ((\$wnnz_Int_resbuf_r  && lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {32'd0,
                                                                         1'd0};
      else if (((! \$wnnz_Int_resbuf_r ) && (! lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet19_4L$wnnz_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int2) : [(lizzieLet19_4Lcall_$wnnz_Int3,Int#),
                                (sc_0_3_destruct,Pointer_CT$wnnz_Int),
                                (q4abZ_1_destruct,Pointer_QTree_Int),
                                (q3abY_1_destruct,Pointer_QTree_Int)] > (lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) */
  assign lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_d = Lcall_$wnnz_Int2_dc((& {lizzieLet19_4Lcall_$wnnz_Int3_d[0],
                                                                                                               sc_0_3_destruct_d[0],
                                                                                                               q4abZ_1_destruct_d[0],
                                                                                                               q3abY_1_destruct_d[0]}), lizzieLet19_4Lcall_$wnnz_Int3_d, sc_0_3_destruct_d, q4abZ_1_destruct_d, q3abY_1_destruct_d);
  assign {lizzieLet19_4Lcall_$wnnz_Int3_r,
          sc_0_3_destruct_r,
          q4abZ_1_destruct_r,
          q3abY_1_destruct_r} = {4 {(lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_r && lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2,CT$wnnz_Int) > (lizzieLet20_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d;
  logic lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_r;
  assign lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_r = ((! lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d[0]) || lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_r)
        lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d <= lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_d;
  CT$wnnz_Int_t lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf;
  assign lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_r = (! lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf[0]);
  assign lizzieLet20_1_argbuf_d = (lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf[0] ? lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf :
                                   lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet20_1_argbuf_r && lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf[0]))
        lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet20_1_argbuf_r) && (! lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf[0])))
        lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_buf <= lizzieLet19_4Lcall_$wnnz_Int3_1sc_0_3_1q4abZ_1_1q3abY_1_1Lcall_$wnnz_Int2_bufchan_d;
  
  /* buf (Ty Bool) : (lizzieLet1_1wild1X19_1_Eq,Bool) > (lizzieLet2_1_argbuf,Bool) */
  Bool_t lizzieLet1_1wild1X19_1_Eq_bufchan_d;
  logic lizzieLet1_1wild1X19_1_Eq_bufchan_r;
  assign lizzieLet1_1wild1X19_1_Eq_r = ((! lizzieLet1_1wild1X19_1_Eq_bufchan_d[0]) || lizzieLet1_1wild1X19_1_Eq_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X19_1_Eq_bufchan_d <= {1'd0, 1'd0};
    else
      if (lizzieLet1_1wild1X19_1_Eq_r)
        lizzieLet1_1wild1X19_1_Eq_bufchan_d <= lizzieLet1_1wild1X19_1_Eq_d;
  Bool_t lizzieLet1_1wild1X19_1_Eq_bufchan_buf;
  assign lizzieLet1_1wild1X19_1_Eq_bufchan_r = (! lizzieLet1_1wild1X19_1_Eq_bufchan_buf[0]);
  assign lizzieLet2_1_argbuf_d = (lizzieLet1_1wild1X19_1_Eq_bufchan_buf[0] ? lizzieLet1_1wild1X19_1_Eq_bufchan_buf :
                                  lizzieLet1_1wild1X19_1_Eq_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet1_1wild1X19_1_Eq_bufchan_buf <= {1'd0, 1'd0};
    else
      if ((lizzieLet2_1_argbuf_r && lizzieLet1_1wild1X19_1_Eq_bufchan_buf[0]))
        lizzieLet1_1wild1X19_1_Eq_bufchan_buf <= {1'd0, 1'd0};
      else if (((! lizzieLet2_1_argbuf_r) && (! lizzieLet1_1wild1X19_1_Eq_bufchan_buf[0])))
        lizzieLet1_1wild1X19_1_Eq_bufchan_buf <= lizzieLet1_1wild1X19_1_Eq_bufchan_d;
  
  /* destruct (Ty CTf'_f'_Int_Int_Int_Int,
          Dcon Lcall_f'_f'_Int_Int_Int_Int0) : (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0,CTf'_f'_Int_Int_Int_Int) > [(es_12_destruct,Pointer_QTree_Int),
                                                                                                                      (es_13_1_destruct,Pointer_QTree_Int),
                                                                                                                      (es_14_2_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_10_destruct,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [3:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted ;
  logic [3:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_done ;
  assign es_12_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [19:4],
                             (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted [0]))};
  assign es_13_1_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [35:20],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted [1]))};
  assign es_14_2_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [51:36],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted [2]))};
  assign sc_0_10_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [67:52],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted [3]))};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_done  = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted  | ({sc_0_10_destruct_d[0],
                                                                                                                     es_14_2_destruct_d[0],
                                                                                                                     es_13_1_destruct_d[0],
                                                                                                                     es_12_destruct_d[0]} & {sc_0_10_destruct_r,
                                                                                                                                             es_14_2_destruct_r,
                                                                                                                                             es_13_1_destruct_r,
                                                                                                                                             es_12_destruct_r}));
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_r  = (& \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted  <= 4'd0;
    else
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_emitted  <= (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_r  ? 4'd0 :
                                                              \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_done );
  
  /* destruct (Ty CTf'_f'_Int_Int_Int_Int,
          Dcon Lcall_f'_f'_Int_Int_Int_Int1) : (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1,CTf'_f'_Int_Int_Int_Int) > [(es_13_destruct,Pointer_QTree_Int),
                                                                                                                      (es_14_1_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_9_destruct,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                      (q1aic_3_destruct,Pointer_QTree_Int),
                                                                                                                      (is_z_kronai6_4_destruct,MyDTInt_Bool),
                                                                                                                      (op_kronai7_4_destruct,MyDTInt_Int_Int),
                                                                                                                      (vai8_4_destruct,Int),
                                                                                                                      (is_z_mapai9_4_destruct,MyDTInt_Bool),
                                                                                                                      (f_mapaia_4_destruct,MyDTInt_Int)] */
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted ;
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_done ;
  assign es_13_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [19:4],
                             (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [0]))};
  assign es_14_1_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [35:20],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [1]))};
  assign sc_0_9_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [51:36],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [2]))};
  assign q1aic_3_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [67:52],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [3]))};
  assign is_z_kronai6_4_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [4]));
  assign op_kronai7_4_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [5]));
  assign vai8_4_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [99:68],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [6]))};
  assign is_z_mapai9_4_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [7]));
  assign f_mapaia_4_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted [8]));
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_done  = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted  | ({f_mapaia_4_destruct_d[0],
                                                                                                                     is_z_mapai9_4_destruct_d[0],
                                                                                                                     vai8_4_destruct_d[0],
                                                                                                                     op_kronai7_4_destruct_d[0],
                                                                                                                     is_z_kronai6_4_destruct_d[0],
                                                                                                                     q1aic_3_destruct_d[0],
                                                                                                                     sc_0_9_destruct_d[0],
                                                                                                                     es_14_1_destruct_d[0],
                                                                                                                     es_13_destruct_d[0]} & {f_mapaia_4_destruct_r,
                                                                                                                                             is_z_mapai9_4_destruct_r,
                                                                                                                                             vai8_4_destruct_r,
                                                                                                                                             op_kronai7_4_destruct_r,
                                                                                                                                             is_z_kronai6_4_destruct_r,
                                                                                                                                             q1aic_3_destruct_r,
                                                                                                                                             sc_0_9_destruct_r,
                                                                                                                                             es_14_1_destruct_r,
                                                                                                                                             es_13_destruct_r}));
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_r  = (& \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted  <= 9'd0;
    else
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_emitted  <= (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_r  ? 9'd0 :
                                                              \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_done );
  
  /* destruct (Ty CTf'_f'_Int_Int_Int_Int,
          Dcon Lcall_f'_f'_Int_Int_Int_Int2) : (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2,CTf'_f'_Int_Int_Int_Int) > [(es_14_destruct,Pointer_QTree_Int),
                                                                                                                      (sc_0_8_destruct,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                      (q1aic_2_destruct,Pointer_QTree_Int),
                                                                                                                      (is_z_kronai6_3_destruct,MyDTInt_Bool),
                                                                                                                      (op_kronai7_3_destruct,MyDTInt_Int_Int),
                                                                                                                      (vai8_3_destruct,Int),
                                                                                                                      (is_z_mapai9_3_destruct,MyDTInt_Bool),
                                                                                                                      (f_mapaia_3_destruct,MyDTInt_Int),
                                                                                                                      (q2aid_2_destruct,Pointer_QTree_Int)] */
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted ;
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_done ;
  assign es_14_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [19:4],
                             (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [0]))};
  assign sc_0_8_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [35:20],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [1]))};
  assign q1aic_2_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [51:36],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [2]))};
  assign is_z_kronai6_3_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [3]));
  assign op_kronai7_3_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [4]));
  assign vai8_3_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [83:52],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [5]))};
  assign is_z_mapai9_3_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [6]));
  assign f_mapaia_3_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [7]));
  assign q2aid_2_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [99:84],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted [8]))};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_done  = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted  | ({q2aid_2_destruct_d[0],
                                                                                                                     f_mapaia_3_destruct_d[0],
                                                                                                                     is_z_mapai9_3_destruct_d[0],
                                                                                                                     vai8_3_destruct_d[0],
                                                                                                                     op_kronai7_3_destruct_d[0],
                                                                                                                     is_z_kronai6_3_destruct_d[0],
                                                                                                                     q1aic_2_destruct_d[0],
                                                                                                                     sc_0_8_destruct_d[0],
                                                                                                                     es_14_destruct_d[0]} & {q2aid_2_destruct_r,
                                                                                                                                             f_mapaia_3_destruct_r,
                                                                                                                                             is_z_mapai9_3_destruct_r,
                                                                                                                                             vai8_3_destruct_r,
                                                                                                                                             op_kronai7_3_destruct_r,
                                                                                                                                             is_z_kronai6_3_destruct_r,
                                                                                                                                             q1aic_2_destruct_r,
                                                                                                                                             sc_0_8_destruct_r,
                                                                                                                                             es_14_destruct_r}));
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_r  = (& \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted  <= 9'd0;
    else
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_emitted  <= (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_r  ? 9'd0 :
                                                              \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_done );
  
  /* destruct (Ty CTf'_f'_Int_Int_Int_Int,
          Dcon Lcall_f'_f'_Int_Int_Int_Int3) : (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3,CTf'_f'_Int_Int_Int_Int) > [(sc_0_7_destruct,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                      (q1aic_1_destruct,Pointer_QTree_Int),
                                                                                                                      (is_z_kronai6_2_destruct,MyDTInt_Bool),
                                                                                                                      (op_kronai7_2_destruct,MyDTInt_Int_Int),
                                                                                                                      (vai8_2_destruct,Int),
                                                                                                                      (is_z_mapai9_2_destruct,MyDTInt_Bool),
                                                                                                                      (f_mapaia_2_destruct,MyDTInt_Int),
                                                                                                                      (q2aid_1_destruct,Pointer_QTree_Int),
                                                                                                                      (q3aie_1_destruct,Pointer_QTree_Int)] */
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted ;
  logic [8:0] \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_done ;
  assign sc_0_7_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [19:4],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [0]))};
  assign q1aic_1_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [35:20],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [1]))};
  assign is_z_kronai6_2_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [2]));
  assign op_kronai7_2_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [3]));
  assign vai8_2_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [67:36],
                              (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [4]))};
  assign is_z_mapai9_2_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [5]));
  assign f_mapaia_2_destruct_d = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [6]));
  assign q2aid_1_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [83:68],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [7]))};
  assign q3aie_1_destruct_d = {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [99:84],
                               (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d [0] && (! \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted [8]))};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_done  = (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted  | ({q3aie_1_destruct_d[0],
                                                                                                                     q2aid_1_destruct_d[0],
                                                                                                                     f_mapaia_2_destruct_d[0],
                                                                                                                     is_z_mapai9_2_destruct_d[0],
                                                                                                                     vai8_2_destruct_d[0],
                                                                                                                     op_kronai7_2_destruct_d[0],
                                                                                                                     is_z_kronai6_2_destruct_d[0],
                                                                                                                     q1aic_1_destruct_d[0],
                                                                                                                     sc_0_7_destruct_d[0]} & {q3aie_1_destruct_r,
                                                                                                                                              q2aid_1_destruct_r,
                                                                                                                                              f_mapaia_2_destruct_r,
                                                                                                                                              is_z_mapai9_2_destruct_r,
                                                                                                                                              vai8_2_destruct_r,
                                                                                                                                              op_kronai7_2_destruct_r,
                                                                                                                                              is_z_kronai6_2_destruct_r,
                                                                                                                                              q1aic_1_destruct_r,
                                                                                                                                              sc_0_7_destruct_r}));
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_r  = (& \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted  <= 9'd0;
    else
      \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_emitted  <= (\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_r  ? 9'd0 :
                                                              \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_done );
  
  /* demux (Ty CTf'_f'_Int_Int_Int_Int,
       Ty CTf'_f'_Int_Int_Int_Int) : (lizzieLet23_2,CTf'_f'_Int_Int_Int_Int) (lizzieLet23_1,CTf'_f'_Int_Int_Int_Int) > [(_18,CTf'_f'_Int_Int_Int_Int),
                                                                                                                        (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3,CTf'_f'_Int_Int_Int_Int),
                                                                                                                        (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2,CTf'_f'_Int_Int_Int_Int),
                                                                                                                        (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1,CTf'_f'_Int_Int_Int_Int),
                                                                                                                        (lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0,CTf'_f'_Int_Int_Int_Int)] */
  logic [4:0] lizzieLet23_1_onehotd;
  always_comb
    if ((lizzieLet23_2_d[0] && lizzieLet23_1_d[0]))
      unique case (lizzieLet23_2_d[3:1])
        3'd0: lizzieLet23_1_onehotd = 5'd1;
        3'd1: lizzieLet23_1_onehotd = 5'd2;
        3'd2: lizzieLet23_1_onehotd = 5'd4;
        3'd3: lizzieLet23_1_onehotd = 5'd8;
        3'd4: lizzieLet23_1_onehotd = 5'd16;
        default: lizzieLet23_1_onehotd = 5'd0;
      endcase
    else lizzieLet23_1_onehotd = 5'd0;
  assign _18_d = {lizzieLet23_1_d[99:1], lizzieLet23_1_onehotd[0]};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_d  = {lizzieLet23_1_d[99:1],
                                                          lizzieLet23_1_onehotd[1]};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_d  = {lizzieLet23_1_d[99:1],
                                                          lizzieLet23_1_onehotd[2]};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_d  = {lizzieLet23_1_d[99:1],
                                                          lizzieLet23_1_onehotd[3]};
  assign \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_d  = {lizzieLet23_1_d[99:1],
                                                          lizzieLet23_1_onehotd[4]};
  assign lizzieLet23_1_r = (| (lizzieLet23_1_onehotd & {\lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int0_r ,
                                                        \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int1_r ,
                                                        \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int2_r ,
                                                        \lizzieLet23_1Lcall_f'_f'_Int_Int_Int_Int3_r ,
                                                        _18_r}));
  assign lizzieLet23_2_r = lizzieLet23_1_r;
  
  /* demux (Ty CTf'_f'_Int_Int_Int_Int,
       Ty Go) : (lizzieLet23_3,CTf'_f'_Int_Int_Int_Int) (go_16_goMux_data,Go) > [(_17,Go),
                                                                                 (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3,Go),
                                                                                 (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2,Go),
                                                                                 (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1,Go),
                                                                                 (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0,Go)] */
  logic [4:0] go_16_goMux_data_onehotd;
  always_comb
    if ((lizzieLet23_3_d[0] && go_16_goMux_data_d[0]))
      unique case (lizzieLet23_3_d[3:1])
        3'd0: go_16_goMux_data_onehotd = 5'd1;
        3'd1: go_16_goMux_data_onehotd = 5'd2;
        3'd2: go_16_goMux_data_onehotd = 5'd4;
        3'd3: go_16_goMux_data_onehotd = 5'd8;
        3'd4: go_16_goMux_data_onehotd = 5'd16;
        default: go_16_goMux_data_onehotd = 5'd0;
      endcase
    else go_16_goMux_data_onehotd = 5'd0;
  assign _17_d = go_16_goMux_data_onehotd[0];
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_d  = go_16_goMux_data_onehotd[1];
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_d  = go_16_goMux_data_onehotd[2];
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_d  = go_16_goMux_data_onehotd[3];
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_d  = go_16_goMux_data_onehotd[4];
  assign go_16_goMux_data_r = (| (go_16_goMux_data_onehotd & {\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_r ,
                                                              \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_r ,
                                                              \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_r ,
                                                              \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_r ,
                                                              _17_r}));
  assign lizzieLet23_3_r = go_16_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0,Go) > (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf,Go) */
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_r  = ((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d [0]) || \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_r )
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_d ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r  = (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0]);
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_d  = (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  :
                                                                   \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_r  && \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_r ) && (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1,Go) > (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf,Go) */
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_r  = ((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d [0]) || \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_r )
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_d ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r  = (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0]);
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_d  = (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  :
                                                                   \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_r  && \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_1_argbuf_r ) && (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2,Go) > (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf,Go) */
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_r  = ((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d [0]) || \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_r )
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_d ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r  = (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0]);
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_d  = (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  :
                                                                   \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_r  && \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_1_argbuf_r ) && (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d ;
  
  /* buf (Ty Go) : (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3,Go) > (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf,Go) */
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_r  = ((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d [0]) || \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d  <= 1'd0;
    else
      if (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_r )
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_d ;
  Go_t \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r  = (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0]);
  assign \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_d  = (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  :
                                                                   \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= 1'd0;
    else
      if ((\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_r  && \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= 1'd0;
      else if (((! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_1_argbuf_r ) && (! \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d ;
  
  /* demux (Ty CTf'_f'_Int_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet23_4,CTf'_f'_Int_Int_Int_Int) (srtarg_0_1_goMux_mux,Pointer_QTree_Int) > [(lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                   (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                   (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                   (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                   (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet23_4_d[0] && srtarg_0_1_goMux_mux_d[0]))
      unique case (lizzieLet23_4_d[3:1])
        3'd0: srtarg_0_1_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_1_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_1_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_1_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_1_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_1_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_1_goMux_mux_onehotd = 5'd0;
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                        srtarg_0_1_goMux_mux_onehotd[0]};
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                          srtarg_0_1_goMux_mux_onehotd[1]};
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                          srtarg_0_1_goMux_mux_onehotd[2]};
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                          srtarg_0_1_goMux_mux_onehotd[3]};
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_d  = {srtarg_0_1_goMux_mux_d[16:1],
                                                          srtarg_0_1_goMux_mux_onehotd[4]};
  assign srtarg_0_1_goMux_mux_r = (| (srtarg_0_1_goMux_mux_onehotd & {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_r ,
                                                                      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_r ,
                                                                      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_r ,
                                                                      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_r ,
                                                                      \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_r }));
  assign lizzieLet23_4_r = srtarg_0_1_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0,Pointer_QTree_Int),
                         (es_12_destruct,Pointer_QTree_Int),
                         (es_13_1_destruct,Pointer_QTree_Int),
                         (es_14_2_destruct,Pointer_QTree_Int)] > (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int,QTree_Int) */
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d  = QNode_Int_dc((& {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_d [0],
                                                                                                              es_12_destruct_d[0],
                                                                                                              es_13_1_destruct_d[0],
                                                                                                              es_14_2_destruct_d[0]}), \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_d , es_12_destruct_d, es_13_1_destruct_d, es_14_2_destruct_d);
  assign {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_r ,
          es_12_destruct_r,
          es_13_1_destruct_r,
          es_14_2_destruct_r} = {4 {(\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r  && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d [0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int,QTree_Int) > (lizzieLet27_1_argbuf,QTree_Int) */
  QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r  = ((! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d [0]) || \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d  <= {66'd0,
                                                                                                    1'd0};
    else
      if (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_r )
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_d ;
  QTree_Int_t \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_r  = (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf [0]);
  assign lizzieLet27_1_argbuf_d = (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf [0] ? \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf  :
                                   \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                      1'd0};
    else
      if ((lizzieLet27_1_argbuf_r && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf [0]))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf  <= {66'd0,
                                                                                                        1'd0};
      else if (((! lizzieLet27_1_argbuf_r) && (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf [0])))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_buf  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int0_1es_12_1es_13_1_1es_14_2_1QNode_Int_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int_Int_Int_Int,
      Dcon Lcall_f'_f'_Int_Int_Int_Int0) : [(lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1,Pointer_QTree_Int),
                                            (es_13_destruct,Pointer_QTree_Int),
                                            (es_14_1_destruct,Pointer_QTree_Int),
                                            (sc_0_9_destruct,Pointer_CTf'_f'_Int_Int_Int_Int)] > (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0,CTf'_f'_Int_Int_Int_Int) */
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_d  = \Lcall_f'_f'_Int_Int_Int_Int0_dc ((& {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_d [0],
                                                                                                                                                     es_13_destruct_d[0],
                                                                                                                                                     es_14_1_destruct_d[0],
                                                                                                                                                     sc_0_9_destruct_d[0]}), \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_d , es_13_destruct_d, es_14_1_destruct_d, sc_0_9_destruct_d);
  assign {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_r ,
          es_13_destruct_r,
          es_14_1_destruct_r,
          sc_0_9_destruct_r} = {4 {(\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_r  && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_d [0])}};
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0,CTf'_f'_Int_Int_Int_Int) > (lizzieLet26_1_argbuf,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_r  = ((! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d [0]) || \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d  <= {99'd0,
                                                                                                                      1'd0};
    else
      if (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_r )
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_r  = (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0]);
  assign lizzieLet26_1_argbuf_d = (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0] ? \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  :
                                   \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                        1'd0};
    else
      if ((lizzieLet26_1_argbuf_r && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0]))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= {99'd0,
                                                                                                                          1'd0};
      else if (((! lizzieLet26_1_argbuf_r) && (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf [0])))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_buf  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int1_1es_13_1es_14_1_1sc_0_9_1Lcall_f'_f'_Int_Int_Int_Int0_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int_Int_Int_Int,
      Dcon Lcall_f'_f'_Int_Int_Int_Int1) : [(lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2,Pointer_QTree_Int),
                                            (es_14_destruct,Pointer_QTree_Int),
                                            (sc_0_8_destruct,Pointer_CTf'_f'_Int_Int_Int_Int),
                                            (q1aic_2_destruct,Pointer_QTree_Int),
                                            (is_z_kronai6_3_1,MyDTInt_Bool),
                                            (op_kronai7_3_1,MyDTInt_Int_Int),
                                            (vai8_3_1,Int),
                                            (is_z_mapai9_3_1,MyDTInt_Bool),
                                            (f_mapaia_3_1,MyDTInt_Int)] > (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1,CTf'_f'_Int_Int_Int_Int) */
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_d  = \Lcall_f'_f'_Int_Int_Int_Int1_dc ((& {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_d [0],
                                                                                                                                                                                                                      es_14_destruct_d[0],
                                                                                                                                                                                                                      sc_0_8_destruct_d[0],
                                                                                                                                                                                                                      q1aic_2_destruct_d[0],
                                                                                                                                                                                                                      is_z_kronai6_3_1_d[0],
                                                                                                                                                                                                                      op_kronai7_3_1_d[0],
                                                                                                                                                                                                                      vai8_3_1_d[0],
                                                                                                                                                                                                                      is_z_mapai9_3_1_d[0],
                                                                                                                                                                                                                      f_mapaia_3_1_d[0]}), \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_d , es_14_destruct_d, sc_0_8_destruct_d, q1aic_2_destruct_d, is_z_kronai6_3_1_d, op_kronai7_3_1_d, vai8_3_1_d, is_z_mapai9_3_1_d, f_mapaia_3_1_d);
  assign {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_r ,
          es_14_destruct_r,
          sc_0_8_destruct_r,
          q1aic_2_destruct_r,
          is_z_kronai6_3_1_r,
          op_kronai7_3_1_r,
          vai8_3_1_r,
          is_z_mapai9_3_1_r,
          f_mapaia_3_1_r} = {9 {(\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_r  && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_d [0])}};
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1,CTf'_f'_Int_Int_Int_Int) > (lizzieLet25_1_argbuf,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_r  = ((! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d [0]) || \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d  <= {99'd0,
                                                                                                                                                                                       1'd0};
    else
      if (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_r )
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_r  = (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0]);
  assign lizzieLet25_1_argbuf_d = (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0] ? \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  :
                                   \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                                                         1'd0};
    else
      if ((lizzieLet25_1_argbuf_r && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0]))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= {99'd0,
                                                                                                                                                                                           1'd0};
      else if (((! lizzieLet25_1_argbuf_r) && (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf [0])))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_buf  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int2_1es_14_1sc_0_8_1q1aic_2_1is_z_kronai6_3_1op_kronai7_3_1vai8_3_1is_z_mapai9_3_1f_mapaia_3_1Lcall_f'_f'_Int_Int_Int_Int1_bufchan_d ;
  
  /* dcon (Ty CTf'_f'_Int_Int_Int_Int,
      Dcon Lcall_f'_f'_Int_Int_Int_Int2) : [(lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3,Pointer_QTree_Int),
                                            (sc_0_7_destruct,Pointer_CTf'_f'_Int_Int_Int_Int),
                                            (q1aic_1_destruct,Pointer_QTree_Int),
                                            (is_z_kronai6_2_1,MyDTInt_Bool),
                                            (op_kronai7_2_1,MyDTInt_Int_Int),
                                            (vai8_2_1,Int),
                                            (is_z_mapai9_2_1,MyDTInt_Bool),
                                            (f_mapaia_2_1,MyDTInt_Int),
                                            (q2aid_1_destruct,Pointer_QTree_Int)] > (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2,CTf'_f'_Int_Int_Int_Int) */
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_d  = \Lcall_f'_f'_Int_Int_Int_Int2_dc ((& {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_d [0],
                                                                                                                                                                                                                        sc_0_7_destruct_d[0],
                                                                                                                                                                                                                        q1aic_1_destruct_d[0],
                                                                                                                                                                                                                        is_z_kronai6_2_1_d[0],
                                                                                                                                                                                                                        op_kronai7_2_1_d[0],
                                                                                                                                                                                                                        vai8_2_1_d[0],
                                                                                                                                                                                                                        is_z_mapai9_2_1_d[0],
                                                                                                                                                                                                                        f_mapaia_2_1_d[0],
                                                                                                                                                                                                                        q2aid_1_destruct_d[0]}), \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_d , sc_0_7_destruct_d, q1aic_1_destruct_d, is_z_kronai6_2_1_d, op_kronai7_2_1_d, vai8_2_1_d, is_z_mapai9_2_1_d, f_mapaia_2_1_d, q2aid_1_destruct_d);
  assign {\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_r ,
          sc_0_7_destruct_r,
          q1aic_1_destruct_r,
          is_z_kronai6_2_1_r,
          op_kronai7_2_1_r,
          vai8_2_1_r,
          is_z_mapai9_2_1_r,
          f_mapaia_2_1_r,
          q2aid_1_destruct_r} = {9 {(\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_r  && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_d [0])}};
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2,CTf'_f'_Int_Int_Int_Int) > (lizzieLet24_1_argbuf,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d ;
  logic \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_r  = ((! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d [0]) || \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d  <= {99'd0,
                                                                                                                                                                                         1'd0};
    else
      if (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_r )
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf ;
  assign \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_r  = (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0]);
  assign lizzieLet24_1_argbuf_d = (\lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0] ? \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  :
                                   \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                                                           1'd0};
    else
      if ((lizzieLet24_1_argbuf_r && \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0]))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= {99'd0,
                                                                                                                                                                                             1'd0};
      else if (((! lizzieLet24_1_argbuf_r) && (! \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf [0])))
        \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_buf  <= \lizzieLet23_4Lcall_f'_f'_Int_Int_Int_Int3_1sc_0_7_1q1aic_1_1is_z_kronai6_2_1op_kronai7_2_1vai8_2_1is_z_mapai9_2_1f_mapaia_2_1q2aid_1_1Lcall_f'_f'_Int_Int_Int_Int2_bufchan_d ;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                             (lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted ;
  logic [1:0] \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_done ;
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d  = {\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d [16:1],
                                                                             (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d [0] && (! \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted [0]))};
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d  = {\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d [16:1],
                                                                             (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_d [0] && (! \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted [1]))};
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_done  = (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted  | ({\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d [0],
                                                                                                                 \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d [0]} & {\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r ,
                                                                                                                                                                                         \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r }));
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_r  = (& \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted  <= 2'd0;
    else
      \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_emitted  <= (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_r  ? 2'd0 :
                                                            \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_done );
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f'_f'_Int_Int_Int_Int_goConst,Go) */
  assign \call_f'_f'_Int_Int_Int_Int_goConst_d  = \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d [0];
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r  = \call_f'_f'_Int_Int_Int_Int_goConst_r ;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (f'_f'_Int_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  logic \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r ;
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r  = ((! \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d [0]) || \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= {16'd0,
                                                                                   1'd0};
    else
      if (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r )
        \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d  <= \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d ;
  Pointer_QTree_Int_t \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf ;
  assign \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r  = (! \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]);
  assign \f'_f'_Int_Int_Int_Int_resbuf_d  = (\lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0] ? \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  :
                                             \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                     1'd0};
    else
      if ((\f'_f'_Int_Int_Int_Int_resbuf_r  && \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0]))
        \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= {16'd0,
                                                                                       1'd0};
      else if (((! \f'_f'_Int_Int_Int_Int_resbuf_r ) && (! \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf [0])))
        \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf  <= \lizzieLet23_4Lf'_f'_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d ;
  
  /* destruct (Ty CTf_f_Int_Int_Int_Int,
          Dcon Lcall_f_f_Int_Int_Int_Int0) : (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0,CTf_f_Int_Int_Int_Int) > [(es_1_1_destruct,Pointer_QTree_Int),
                                                                                                                (es_2_2_destruct,Pointer_QTree_Int),
                                                                                                                (es_3_3_destruct,Pointer_QTree_Int),
                                                                                                                (sc_0_14_destruct,Pointer_CTf_f_Int_Int_Int_Int)] */
  logic [3:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted;
  logic [3:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_done;
  assign es_1_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[19:4],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted[0]))};
  assign es_2_2_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[35:20],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted[1]))};
  assign es_3_3_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[51:36],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted[2]))};
  assign sc_0_14_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[67:52],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted[3]))};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_done = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted | ({sc_0_14_destruct_d[0],
                                                                                                             es_3_3_destruct_d[0],
                                                                                                             es_2_2_destruct_d[0],
                                                                                                             es_1_1_destruct_d[0]} & {sc_0_14_destruct_r,
                                                                                                                                      es_3_3_destruct_r,
                                                                                                                                      es_2_2_destruct_r,
                                                                                                                                      es_1_1_destruct_r}));
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_r = (& lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted <= 4'd0;
    else
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_emitted <= (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_r ? 4'd0 :
                                                          lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_done);
  
  /* destruct (Ty CTf_f_Int_Int_Int_Int,
          Dcon Lcall_f_f_Int_Int_Int_Int1) : (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1,CTf_f_Int_Int_Int_Int) > [(es_2_1_destruct,Pointer_QTree_Int),
                                                                                                                (es_3_2_destruct,Pointer_QTree_Int),
                                                                                                                (sc_0_13_destruct,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                (q1ai1_3_destruct,Pointer_QTree_Int),
                                                                                                                (m2ahV_4_destruct,Pointer_QTree_Int),
                                                                                                                (is_z_kronahW_4_destruct,MyDTInt_Bool),
                                                                                                                (op_kronahX_4_destruct,MyDTInt_Int_Int),
                                                                                                                (is_z_mapahY_4_destruct,MyDTInt_Bool),
                                                                                                                (f_mapahZ_4_destruct,MyDTInt_Int)] */
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted;
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_done;
  assign es_2_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[19:4],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[0]))};
  assign es_3_2_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[35:20],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[1]))};
  assign sc_0_13_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[51:36],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[2]))};
  assign q1ai1_3_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[67:52],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[3]))};
  assign m2ahV_4_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[83:68],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[4]))};
  assign is_z_kronahW_4_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[5]));
  assign op_kronahX_4_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[6]));
  assign is_z_mapahY_4_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[7]));
  assign f_mapahZ_4_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted[8]));
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_done = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted | ({f_mapahZ_4_destruct_d[0],
                                                                                                             is_z_mapahY_4_destruct_d[0],
                                                                                                             op_kronahX_4_destruct_d[0],
                                                                                                             is_z_kronahW_4_destruct_d[0],
                                                                                                             m2ahV_4_destruct_d[0],
                                                                                                             q1ai1_3_destruct_d[0],
                                                                                                             sc_0_13_destruct_d[0],
                                                                                                             es_3_2_destruct_d[0],
                                                                                                             es_2_1_destruct_d[0]} & {f_mapahZ_4_destruct_r,
                                                                                                                                      is_z_mapahY_4_destruct_r,
                                                                                                                                      op_kronahX_4_destruct_r,
                                                                                                                                      is_z_kronahW_4_destruct_r,
                                                                                                                                      m2ahV_4_destruct_r,
                                                                                                                                      q1ai1_3_destruct_r,
                                                                                                                                      sc_0_13_destruct_r,
                                                                                                                                      es_3_2_destruct_r,
                                                                                                                                      es_2_1_destruct_r}));
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_r = (& lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted <= 9'd0;
    else
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_emitted <= (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_r ? 9'd0 :
                                                          lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_done);
  
  /* destruct (Ty CTf_f_Int_Int_Int_Int,
          Dcon Lcall_f_f_Int_Int_Int_Int2) : (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2,CTf_f_Int_Int_Int_Int) > [(es_3_1_destruct,Pointer_QTree_Int),
                                                                                                                (sc_0_12_destruct,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                (q1ai1_2_destruct,Pointer_QTree_Int),
                                                                                                                (m2ahV_3_destruct,Pointer_QTree_Int),
                                                                                                                (is_z_kronahW_3_destruct,MyDTInt_Bool),
                                                                                                                (op_kronahX_3_destruct,MyDTInt_Int_Int),
                                                                                                                (is_z_mapahY_3_destruct,MyDTInt_Bool),
                                                                                                                (f_mapahZ_3_destruct,MyDTInt_Int),
                                                                                                                (q2ai2_2_destruct,Pointer_QTree_Int)] */
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted;
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_done;
  assign es_3_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[19:4],
                              (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[0]))};
  assign sc_0_12_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[35:20],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[1]))};
  assign q1ai1_2_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[51:36],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[2]))};
  assign m2ahV_3_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[67:52],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[3]))};
  assign is_z_kronahW_3_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[4]));
  assign op_kronahX_3_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[5]));
  assign is_z_mapahY_3_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[6]));
  assign f_mapahZ_3_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[7]));
  assign q2ai2_2_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[83:68],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted[8]))};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_done = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted | ({q2ai2_2_destruct_d[0],
                                                                                                             f_mapahZ_3_destruct_d[0],
                                                                                                             is_z_mapahY_3_destruct_d[0],
                                                                                                             op_kronahX_3_destruct_d[0],
                                                                                                             is_z_kronahW_3_destruct_d[0],
                                                                                                             m2ahV_3_destruct_d[0],
                                                                                                             q1ai1_2_destruct_d[0],
                                                                                                             sc_0_12_destruct_d[0],
                                                                                                             es_3_1_destruct_d[0]} & {q2ai2_2_destruct_r,
                                                                                                                                      f_mapahZ_3_destruct_r,
                                                                                                                                      is_z_mapahY_3_destruct_r,
                                                                                                                                      op_kronahX_3_destruct_r,
                                                                                                                                      is_z_kronahW_3_destruct_r,
                                                                                                                                      m2ahV_3_destruct_r,
                                                                                                                                      q1ai1_2_destruct_r,
                                                                                                                                      sc_0_12_destruct_r,
                                                                                                                                      es_3_1_destruct_r}));
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_r = (& lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted <= 9'd0;
    else
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_emitted <= (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_r ? 9'd0 :
                                                          lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_done);
  
  /* destruct (Ty CTf_f_Int_Int_Int_Int,
          Dcon Lcall_f_f_Int_Int_Int_Int3) : (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3,CTf_f_Int_Int_Int_Int) > [(sc_0_11_destruct,Pointer_CTf_f_Int_Int_Int_Int),
                                                                                                                (q1ai1_1_destruct,Pointer_QTree_Int),
                                                                                                                (m2ahV_2_destruct,Pointer_QTree_Int),
                                                                                                                (is_z_kronahW_2_destruct,MyDTInt_Bool),
                                                                                                                (op_kronahX_2_destruct,MyDTInt_Int_Int),
                                                                                                                (is_z_mapahY_2_destruct,MyDTInt_Bool),
                                                                                                                (f_mapahZ_2_destruct,MyDTInt_Int),
                                                                                                                (q2ai2_1_destruct,Pointer_QTree_Int),
                                                                                                                (q3ai3_1_destruct,Pointer_QTree_Int)] */
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted;
  logic [8:0] lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_done;
  assign sc_0_11_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[19:4],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[0]))};
  assign q1ai1_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[35:20],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[1]))};
  assign m2ahV_2_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[51:36],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[2]))};
  assign is_z_kronahW_2_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[3]));
  assign op_kronahX_2_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[4]));
  assign is_z_mapahY_2_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[5]));
  assign f_mapahZ_2_destruct_d = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[6]));
  assign q2ai2_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[67:52],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[7]))};
  assign q3ai3_1_destruct_d = {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[83:68],
                               (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d[0] && (! lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted[8]))};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_done = (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted | ({q3ai3_1_destruct_d[0],
                                                                                                             q2ai2_1_destruct_d[0],
                                                                                                             f_mapahZ_2_destruct_d[0],
                                                                                                             is_z_mapahY_2_destruct_d[0],
                                                                                                             op_kronahX_2_destruct_d[0],
                                                                                                             is_z_kronahW_2_destruct_d[0],
                                                                                                             m2ahV_2_destruct_d[0],
                                                                                                             q1ai1_1_destruct_d[0],
                                                                                                             sc_0_11_destruct_d[0]} & {q3ai3_1_destruct_r,
                                                                                                                                       q2ai2_1_destruct_r,
                                                                                                                                       f_mapahZ_2_destruct_r,
                                                                                                                                       is_z_mapahY_2_destruct_r,
                                                                                                                                       op_kronahX_2_destruct_r,
                                                                                                                                       is_z_kronahW_2_destruct_r,
                                                                                                                                       m2ahV_2_destruct_r,
                                                                                                                                       q1ai1_1_destruct_r,
                                                                                                                                       sc_0_11_destruct_r}));
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_r = (& lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted <= 9'd0;
    else
      lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_emitted <= (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_r ? 9'd0 :
                                                          lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_done);
  
  /* demux (Ty CTf_f_Int_Int_Int_Int,
       Ty CTf_f_Int_Int_Int_Int) : (lizzieLet28_2,CTf_f_Int_Int_Int_Int) (lizzieLet28_1,CTf_f_Int_Int_Int_Int) > [(_16,CTf_f_Int_Int_Int_Int),
                                                                                                                  (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3,CTf_f_Int_Int_Int_Int),
                                                                                                                  (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2,CTf_f_Int_Int_Int_Int),
                                                                                                                  (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1,CTf_f_Int_Int_Int_Int),
                                                                                                                  (lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0,CTf_f_Int_Int_Int_Int)] */
  logic [4:0] lizzieLet28_1_onehotd;
  always_comb
    if ((lizzieLet28_2_d[0] && lizzieLet28_1_d[0]))
      unique case (lizzieLet28_2_d[3:1])
        3'd0: lizzieLet28_1_onehotd = 5'd1;
        3'd1: lizzieLet28_1_onehotd = 5'd2;
        3'd2: lizzieLet28_1_onehotd = 5'd4;
        3'd3: lizzieLet28_1_onehotd = 5'd8;
        3'd4: lizzieLet28_1_onehotd = 5'd16;
        default: lizzieLet28_1_onehotd = 5'd0;
      endcase
    else lizzieLet28_1_onehotd = 5'd0;
  assign _16_d = {lizzieLet28_1_d[83:1], lizzieLet28_1_onehotd[0]};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_d = {lizzieLet28_1_d[83:1],
                                                      lizzieLet28_1_onehotd[1]};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_d = {lizzieLet28_1_d[83:1],
                                                      lizzieLet28_1_onehotd[2]};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_d = {lizzieLet28_1_d[83:1],
                                                      lizzieLet28_1_onehotd[3]};
  assign lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_d = {lizzieLet28_1_d[83:1],
                                                      lizzieLet28_1_onehotd[4]};
  assign lizzieLet28_1_r = (| (lizzieLet28_1_onehotd & {lizzieLet28_1Lcall_f_f_Int_Int_Int_Int0_r,
                                                        lizzieLet28_1Lcall_f_f_Int_Int_Int_Int1_r,
                                                        lizzieLet28_1Lcall_f_f_Int_Int_Int_Int2_r,
                                                        lizzieLet28_1Lcall_f_f_Int_Int_Int_Int3_r,
                                                        _16_r}));
  assign lizzieLet28_2_r = lizzieLet28_1_r;
  
  /* demux (Ty CTf_f_Int_Int_Int_Int,
       Ty Go) : (lizzieLet28_3,CTf_f_Int_Int_Int_Int) (go_17_goMux_data,Go) > [(_15,Go),
                                                                               (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3,Go),
                                                                               (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2,Go),
                                                                               (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1,Go),
                                                                               (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0,Go)] */
  logic [4:0] go_17_goMux_data_onehotd;
  always_comb
    if ((lizzieLet28_3_d[0] && go_17_goMux_data_d[0]))
      unique case (lizzieLet28_3_d[3:1])
        3'd0: go_17_goMux_data_onehotd = 5'd1;
        3'd1: go_17_goMux_data_onehotd = 5'd2;
        3'd2: go_17_goMux_data_onehotd = 5'd4;
        3'd3: go_17_goMux_data_onehotd = 5'd8;
        3'd4: go_17_goMux_data_onehotd = 5'd16;
        default: go_17_goMux_data_onehotd = 5'd0;
      endcase
    else go_17_goMux_data_onehotd = 5'd0;
  assign _15_d = go_17_goMux_data_onehotd[0];
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_d = go_17_goMux_data_onehotd[1];
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_d = go_17_goMux_data_onehotd[2];
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_d = go_17_goMux_data_onehotd[3];
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_d = go_17_goMux_data_onehotd[4];
  assign go_17_goMux_data_r = (| (go_17_goMux_data_onehotd & {lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_r,
                                                              lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_r,
                                                              lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_r,
                                                              lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_r,
                                                              _15_r}));
  assign lizzieLet28_3_r = go_17_goMux_data_r;
  
  /* buf (Ty Go) : (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0,Go) > (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf,Go) */
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_r;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_r = ((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d[0]) || lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d <= 1'd0;
    else
      if (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_r)
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_d;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_r = (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_d = (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0] ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf :
                                                               lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_r && lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= 1'd0;
      else if (((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_1_argbuf_r) && (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1,Go) > (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf,Go) */
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_r;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_r = ((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d[0]) || lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d <= 1'd0;
    else
      if (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_r)
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_d;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_r = (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_d = (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0] ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf :
                                                               lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_r && lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_1_argbuf_r) && (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2,Go) > (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf,Go) */
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_r;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_r = ((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d[0]) || lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d <= 1'd0;
    else
      if (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_r)
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_d;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_r = (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_d = (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0] ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf :
                                                               lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_r && lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_1_argbuf_r) && (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3,Go) > (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf,Go) */
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d;
  logic lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_r;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_r = ((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d[0]) || lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d <= 1'd0;
    else
      if (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_r)
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_d;
  Go_t lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf;
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_r = (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0]);
  assign lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_d = (lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0] ? lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf :
                                                               lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_r && lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0]))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= 1'd0;
      else if (((! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_1_argbuf_r) && (! lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf[0])))
        lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_buf <= lizzieLet28_3Lcall_f_f_Int_Int_Int_Int3_bufchan_d;
  
  /* demux (Ty CTf_f_Int_Int_Int_Int,
       Ty Pointer_QTree_Int) : (lizzieLet28_4,CTf_f_Int_Int_Int_Int) (srtarg_0_2_goMux_mux,Pointer_QTree_Int) > [(lizzieLet28_4Lf_f_Int_Int_Int_Intsbos,Pointer_QTree_Int),
                                                                                                                 (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3,Pointer_QTree_Int),
                                                                                                                 (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2,Pointer_QTree_Int),
                                                                                                                 (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1,Pointer_QTree_Int),
                                                                                                                 (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0,Pointer_QTree_Int)] */
  logic [4:0] srtarg_0_2_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet28_4_d[0] && srtarg_0_2_goMux_mux_d[0]))
      unique case (lizzieLet28_4_d[3:1])
        3'd0: srtarg_0_2_goMux_mux_onehotd = 5'd1;
        3'd1: srtarg_0_2_goMux_mux_onehotd = 5'd2;
        3'd2: srtarg_0_2_goMux_mux_onehotd = 5'd4;
        3'd3: srtarg_0_2_goMux_mux_onehotd = 5'd8;
        3'd4: srtarg_0_2_goMux_mux_onehotd = 5'd16;
        default: srtarg_0_2_goMux_mux_onehotd = 5'd0;
      endcase
    else srtarg_0_2_goMux_mux_onehotd = 5'd0;
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                    srtarg_0_2_goMux_mux_onehotd[0]};
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[1]};
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[2]};
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[3]};
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_d = {srtarg_0_2_goMux_mux_d[16:1],
                                                      srtarg_0_2_goMux_mux_onehotd[4]};
  assign srtarg_0_2_goMux_mux_r = (| (srtarg_0_2_goMux_mux_onehotd & {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_r,
                                                                      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_r,
                                                                      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_r,
                                                                      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_r,
                                                                      lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_r}));
  assign lizzieLet28_4_r = srtarg_0_2_goMux_mux_r;
  
  /* dcon (Ty QTree_Int,
      Dcon QNode_Int) : [(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0,Pointer_QTree_Int),
                         (es_1_1_destruct,Pointer_QTree_Int),
                         (es_2_2_destruct,Pointer_QTree_Int),
                         (es_3_3_destruct,Pointer_QTree_Int)] > (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int,QTree_Int) */
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d = QNode_Int_dc((& {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_d[0],
                                                                                                         es_1_1_destruct_d[0],
                                                                                                         es_2_2_destruct_d[0],
                                                                                                         es_3_3_destruct_d[0]}), lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_d, es_1_1_destruct_d, es_2_2_destruct_d, es_3_3_destruct_d);
  assign {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_r,
          es_1_1_destruct_r,
          es_2_2_destruct_r,
          es_3_3_destruct_r} = {4 {(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int,QTree_Int) > (lizzieLet32_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r = ((! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d[0]) || lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d <= {66'd0,
                                                                                               1'd0};
    else
      if (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_r)
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_d;
  QTree_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_r = (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0]);
  assign lizzieLet32_1_argbuf_d = (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0] ? lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf :
                                   lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet32_1_argbuf_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0]))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= {66'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet32_1_argbuf_r) && (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf[0])))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_buf <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int0_1es_1_1_1es_2_2_1es_3_3_1QNode_Int_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int_Int_Int,
      Dcon Lcall_f_f_Int_Int_Int_Int0) : [(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1,Pointer_QTree_Int),
                                          (es_2_1_destruct,Pointer_QTree_Int),
                                          (es_3_2_destruct,Pointer_QTree_Int),
                                          (sc_0_13_destruct,Pointer_CTf_f_Int_Int_Int_Int)] > (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0,CTf_f_Int_Int_Int_Int) */
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_d = Lcall_f_f_Int_Int_Int_Int0_dc((& {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_d[0],
                                                                                                                                            es_2_1_destruct_d[0],
                                                                                                                                            es_3_2_destruct_d[0],
                                                                                                                                            sc_0_13_destruct_d[0]}), lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_d, es_2_1_destruct_d, es_3_2_destruct_d, sc_0_13_destruct_d);
  assign {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_r,
          es_2_1_destruct_r,
          es_3_2_destruct_r,
          sc_0_13_destruct_r} = {4 {(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0,CTf_f_Int_Int_Int_Int) > (lizzieLet31_1_argbuf,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_r;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_r = ((! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d[0]) || lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d <= {83'd0,
                                                                                                                 1'd0};
    else
      if (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_r)
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_d;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_r = (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0]);
  assign lizzieLet31_1_argbuf_d = (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0] ? lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf :
                                   lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                   1'd0};
    else
      if ((lizzieLet31_1_argbuf_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0]))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= {83'd0,
                                                                                                                     1'd0};
      else if (((! lizzieLet31_1_argbuf_r) && (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf[0])))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_buf <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int1_1es_2_1_1es_3_2_1sc_0_13_1Lcall_f_f_Int_Int_Int_Int0_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int_Int_Int,
      Dcon Lcall_f_f_Int_Int_Int_Int1) : [(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2,Pointer_QTree_Int),
                                          (es_3_1_destruct,Pointer_QTree_Int),
                                          (sc_0_12_destruct,Pointer_CTf_f_Int_Int_Int_Int),
                                          (q1ai1_2_destruct,Pointer_QTree_Int),
                                          (m2ahV_3_1,Pointer_QTree_Int),
                                          (is_z_kronahW_3_1,MyDTInt_Bool),
                                          (op_kronahX_3_1,MyDTInt_Int_Int),
                                          (is_z_mapahY_3_1,MyDTInt_Bool),
                                          (f_mapahZ_3_1,MyDTInt_Int)] > (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1,CTf_f_Int_Int_Int_Int) */
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_d = Lcall_f_f_Int_Int_Int_Int1_dc((& {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_d[0],
                                                                                                                                                                                                               es_3_1_destruct_d[0],
                                                                                                                                                                                                               sc_0_12_destruct_d[0],
                                                                                                                                                                                                               q1ai1_2_destruct_d[0],
                                                                                                                                                                                                               m2ahV_3_1_d[0],
                                                                                                                                                                                                               is_z_kronahW_3_1_d[0],
                                                                                                                                                                                                               op_kronahX_3_1_d[0],
                                                                                                                                                                                                               is_z_mapahY_3_1_d[0],
                                                                                                                                                                                                               f_mapahZ_3_1_d[0]}), lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_d, es_3_1_destruct_d, sc_0_12_destruct_d, q1ai1_2_destruct_d, m2ahV_3_1_d, is_z_kronahW_3_1_d, op_kronahX_3_1_d, is_z_mapahY_3_1_d, f_mapahZ_3_1_d);
  assign {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_r,
          es_3_1_destruct_r,
          sc_0_12_destruct_r,
          q1ai1_2_destruct_r,
          m2ahV_3_1_r,
          is_z_kronahW_3_1_r,
          op_kronahX_3_1_r,
          is_z_mapahY_3_1_r,
          f_mapahZ_3_1_r} = {9 {(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1,CTf_f_Int_Int_Int_Int) > (lizzieLet30_1_argbuf,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_r;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_r = ((! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d[0]) || lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d <= {83'd0,
                                                                                                                                                                                    1'd0};
    else
      if (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_r)
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_d;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_r = (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0]);
  assign lizzieLet30_1_argbuf_d = (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0] ? lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf :
                                   lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                                                      1'd0};
    else
      if ((lizzieLet30_1_argbuf_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0]))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= {83'd0,
                                                                                                                                                                                        1'd0};
      else if (((! lizzieLet30_1_argbuf_r) && (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf[0])))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_buf <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int2_1es_3_1_1sc_0_12_1q1ai1_2_1m2ahV_3_1is_z_kronahW_3_1op_kronahX_3_1is_z_mapahY_3_1f_mapahZ_3_1Lcall_f_f_Int_Int_Int_Int1_bufchan_d;
  
  /* dcon (Ty CTf_f_Int_Int_Int_Int,
      Dcon Lcall_f_f_Int_Int_Int_Int2) : [(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3,Pointer_QTree_Int),
                                          (sc_0_11_destruct,Pointer_CTf_f_Int_Int_Int_Int),
                                          (q1ai1_1_destruct,Pointer_QTree_Int),
                                          (m2ahV_2_1,Pointer_QTree_Int),
                                          (is_z_kronahW_2_1,MyDTInt_Bool),
                                          (op_kronahX_2_1,MyDTInt_Int_Int),
                                          (is_z_mapahY_2_1,MyDTInt_Bool),
                                          (f_mapahZ_2_1,MyDTInt_Int),
                                          (q2ai2_1_destruct,Pointer_QTree_Int)] > (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2,CTf_f_Int_Int_Int_Int) */
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_d = Lcall_f_f_Int_Int_Int_Int2_dc((& {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_d[0],
                                                                                                                                                                                                                sc_0_11_destruct_d[0],
                                                                                                                                                                                                                q1ai1_1_destruct_d[0],
                                                                                                                                                                                                                m2ahV_2_1_d[0],
                                                                                                                                                                                                                is_z_kronahW_2_1_d[0],
                                                                                                                                                                                                                op_kronahX_2_1_d[0],
                                                                                                                                                                                                                is_z_mapahY_2_1_d[0],
                                                                                                                                                                                                                f_mapahZ_2_1_d[0],
                                                                                                                                                                                                                q2ai2_1_destruct_d[0]}), lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_d, sc_0_11_destruct_d, q1ai1_1_destruct_d, m2ahV_2_1_d, is_z_kronahW_2_1_d, op_kronahX_2_1_d, is_z_mapahY_2_1_d, f_mapahZ_2_1_d, q2ai2_1_destruct_d);
  assign {lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_r,
          sc_0_11_destruct_r,
          q1ai1_1_destruct_r,
          m2ahV_2_1_r,
          is_z_kronahW_2_1_r,
          op_kronahX_2_1_r,
          is_z_mapahY_2_1_r,
          f_mapahZ_2_1_r,
          q2ai2_1_destruct_r} = {9 {(lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_d[0])}};
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2,CTf_f_Int_Int_Int_Int) > (lizzieLet29_1_argbuf,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d;
  logic lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_r;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_r = ((! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d[0]) || lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d <= {83'd0,
                                                                                                                                                                                     1'd0};
    else
      if (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_r)
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_d;
  CTf_f_Int_Int_Int_Int_t lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf;
  assign lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_r = (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0]);
  assign lizzieLet29_1_argbuf_d = (lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0] ? lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf :
                                   lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                                                       1'd0};
    else
      if ((lizzieLet29_1_argbuf_r && lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0]))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= {83'd0,
                                                                                                                                                                                         1'd0};
      else if (((! lizzieLet29_1_argbuf_r) && (! lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf[0])))
        lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_buf <= lizzieLet28_4Lcall_f_f_Int_Int_Int_Int3_1sc_0_11_1q1ai1_1_1m2ahV_2_1is_z_kronahW_2_1op_kronahX_2_1is_z_mapahY_2_1f_mapahZ_2_1q2ai2_1_1Lcall_f_f_Int_Int_Int_Int2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos,Pointer_QTree_Int) > [(lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int),
                                                                                           (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int)] */
  logic [1:0] lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted;
  logic [1:0] lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_done;
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d = {lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d[16:1],
                                                                         (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d[0] && (! lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted[0]))};
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d = {lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d[16:1],
                                                                         (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_d[0] && (! lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted[1]))};
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_done = (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted | ({lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d[0],
                                                                                                         lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d[0]} & {lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r,
                                                                                                                                                                             lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r}));
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_r = (& lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted <= 2'd0;
    else
      lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_emitted <= (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_r ? 2'd0 :
                                                        lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_done);
  
  /* togo (Ty Pointer_QTree_Int) : (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1,Pointer_QTree_Int) > (call_f_f_Int_Int_Int_Int_goConst,Go) */
  assign call_f_f_Int_Int_Int_Int_goConst_d = lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_d[0];
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_1_r = call_f_f_Int_Int_Int_Int_goConst_r;
  
  /* buf (Ty Pointer_QTree_Int) : (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2,Pointer_QTree_Int) > (f_f_Int_Int_Int_Int_resbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  logic lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r;
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r = ((! lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d[0]) || lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= {16'd0,
                                                                               1'd0};
    else
      if (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_r)
        lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d <= lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_d;
  Pointer_QTree_Int_t lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf;
  assign lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_r = (! lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]);
  assign f_f_Int_Int_Int_Int_resbuf_d = (lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0] ? lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf :
                                         lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                 1'd0};
    else
      if ((f_f_Int_Int_Int_Int_resbuf_r && lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0]))
        lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= {16'd0,
                                                                                   1'd0};
      else if (((! f_f_Int_Int_Int_Int_resbuf_r) && (! lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf[0])))
        lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_buf <= lizzieLet28_4Lf_f_Int_Int_Int_Intsbos_1_merge_merge_fork_2_bufchan_d;
  
  /* demux (Ty MyBool,
       Ty Go) : (lizzieLet3_1,MyBool) (arg0_1Dcon_eqZero_3I#_3,Go) > [(lizzieLet3_1MyFalse,Go),
                                                                      (lizzieLet3_1MyTrue,Go)] */
  logic [1:0] \arg0_1Dcon_eqZero_3I#_3_onehotd ;
  always_comb
    if ((lizzieLet3_1_d[0] && \arg0_1Dcon_eqZero_3I#_3_d [0]))
      unique case (lizzieLet3_1_d[1:1])
        1'd0: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd1;
        1'd1: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd2;
        default: \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd0;
      endcase
    else \arg0_1Dcon_eqZero_3I#_3_onehotd  = 2'd0;
  assign lizzieLet3_1MyFalse_d = \arg0_1Dcon_eqZero_3I#_3_onehotd [0];
  assign lizzieLet3_1MyTrue_d = \arg0_1Dcon_eqZero_3I#_3_onehotd [1];
  assign \arg0_1Dcon_eqZero_3I#_3_r  = (| (\arg0_1Dcon_eqZero_3I#_3_onehotd  & {lizzieLet3_1MyTrue_r,
                                                                                lizzieLet3_1MyFalse_r}));
  assign lizzieLet3_1_r = \arg0_1Dcon_eqZero_3I#_3_r ;
  
  /* dcon (Ty MyBool,
      Dcon MyFalse) : [(lizzieLet3_1MyFalse,Go)] > (lizzieLet3_1MyFalse_1MyFalse,MyBool) */
  assign lizzieLet3_1MyFalse_1MyFalse_d = MyFalse_dc((& {lizzieLet3_1MyFalse_d[0]}), lizzieLet3_1MyFalse_d);
  assign {lizzieLet3_1MyFalse_r} = {1 {(lizzieLet3_1MyFalse_1MyFalse_r && lizzieLet3_1MyFalse_1MyFalse_d[0])}};
  
  /* dcon (Ty MyBool,
      Dcon MyTrue) : [(lizzieLet3_1MyTrue,Go)] > (lizzieLet3_1MyTrue_1MyTrue,MyBool) */
  assign lizzieLet3_1MyTrue_1MyTrue_d = MyTrue_dc((& {lizzieLet3_1MyTrue_d[0]}), lizzieLet3_1MyTrue_d);
  assign {lizzieLet3_1MyTrue_r} = {1 {(lizzieLet3_1MyTrue_1MyTrue_r && lizzieLet3_1MyTrue_1MyTrue_d[0])}};
  
  /* mux (Ty MyBool,
     Ty MyBool) : (lizzieLet3_2,MyBool) [(lizzieLet3_1MyFalse_1MyFalse,MyBool),
                                         (lizzieLet3_1MyTrue_1MyTrue,MyBool)] > (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux,MyBool) */
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux;
  logic [1:0] lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot;
  always_comb
    unique case (lizzieLet3_2_d[1:1])
      1'd0:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd1,
                                                                            lizzieLet3_1MyFalse_1MyFalse_d};
      1'd1:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd2,
                                                                            lizzieLet3_1MyTrue_1MyTrue_d};
      default:
        {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot,
         lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux} = {2'd0,
                                                                            {1'd0, 1'd0}};
    endcase
  assign lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d = {lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[1:1],
                                                                         (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_mux[0] && lizzieLet3_2_d[0])};
  assign lizzieLet3_2_r = (lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_d[0] && lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_r);
  assign {lizzieLet3_1MyTrue_1MyTrue_r,
          lizzieLet3_1MyFalse_1MyFalse_r} = (lizzieLet3_2_r ? lizzieLet3_1MyFalse_1MyFalselizzieLet3_1MyTrue_1MyTrue_mux_onehot :
                                             2'd0);
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet4_1QNode_Int,QTree_Int) > [(q1abW_destruct,Pointer_QTree_Int),
                                                                 (q2abX_destruct,Pointer_QTree_Int),
                                                                 (q3abY_destruct,Pointer_QTree_Int),
                                                                 (q4abZ_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet4_1QNode_Int_emitted;
  logic [3:0] lizzieLet4_1QNode_Int_done;
  assign q1abW_destruct_d = {lizzieLet4_1QNode_Int_d[18:3],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[0]))};
  assign q2abX_destruct_d = {lizzieLet4_1QNode_Int_d[34:19],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[1]))};
  assign q3abY_destruct_d = {lizzieLet4_1QNode_Int_d[50:35],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[2]))};
  assign q4abZ_destruct_d = {lizzieLet4_1QNode_Int_d[66:51],
                             (lizzieLet4_1QNode_Int_d[0] && (! lizzieLet4_1QNode_Int_emitted[3]))};
  assign lizzieLet4_1QNode_Int_done = (lizzieLet4_1QNode_Int_emitted | ({q4abZ_destruct_d[0],
                                                                         q3abY_destruct_d[0],
                                                                         q2abX_destruct_d[0],
                                                                         q1abW_destruct_d[0]} & {q4abZ_destruct_r,
                                                                                                 q3abY_destruct_r,
                                                                                                 q2abX_destruct_r,
                                                                                                 q1abW_destruct_r}));
  assign lizzieLet4_1QNode_Int_r = (& lizzieLet4_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet4_1QNode_Int_emitted <= (lizzieLet4_1QNode_Int_r ? 4'd0 :
                                        lizzieLet4_1QNode_Int_done);
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet4_2,QTree_Int) (lizzieLet4_1,QTree_Int) > [(_14,QTree_Int),
                                                                            (_13,QTree_Int),
                                                                            (lizzieLet4_1QNode_Int,QTree_Int),
                                                                            (_12,QTree_Int)] */
  logic [3:0] lizzieLet4_1_onehotd;
  always_comb
    if ((lizzieLet4_2_d[0] && lizzieLet4_1_d[0]))
      unique case (lizzieLet4_2_d[2:1])
        2'd0: lizzieLet4_1_onehotd = 4'd1;
        2'd1: lizzieLet4_1_onehotd = 4'd2;
        2'd2: lizzieLet4_1_onehotd = 4'd4;
        2'd3: lizzieLet4_1_onehotd = 4'd8;
        default: lizzieLet4_1_onehotd = 4'd0;
      endcase
    else lizzieLet4_1_onehotd = 4'd0;
  assign _14_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[0]};
  assign _13_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[1]};
  assign lizzieLet4_1QNode_Int_d = {lizzieLet4_1_d[66:1],
                                    lizzieLet4_1_onehotd[2]};
  assign _12_d = {lizzieLet4_1_d[66:1], lizzieLet4_1_onehotd[3]};
  assign lizzieLet4_1_r = (| (lizzieLet4_1_onehotd & {_12_r,
                                                      lizzieLet4_1QNode_Int_r,
                                                      _13_r,
                                                      _14_r}));
  assign lizzieLet4_2_r = lizzieLet4_1_r;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet4_3,QTree_Int) (go_10_goMux_data,Go) > [(lizzieLet4_3QNone_Int,Go),
                                                                  (lizzieLet4_3QVal_Int,Go),
                                                                  (lizzieLet4_3QNode_Int,Go),
                                                                  (lizzieLet4_3QError_Int,Go)] */
  logic [3:0] go_10_goMux_data_onehotd;
  always_comb
    if ((lizzieLet4_3_d[0] && go_10_goMux_data_d[0]))
      unique case (lizzieLet4_3_d[2:1])
        2'd0: go_10_goMux_data_onehotd = 4'd1;
        2'd1: go_10_goMux_data_onehotd = 4'd2;
        2'd2: go_10_goMux_data_onehotd = 4'd4;
        2'd3: go_10_goMux_data_onehotd = 4'd8;
        default: go_10_goMux_data_onehotd = 4'd0;
      endcase
    else go_10_goMux_data_onehotd = 4'd0;
  assign lizzieLet4_3QNone_Int_d = go_10_goMux_data_onehotd[0];
  assign lizzieLet4_3QVal_Int_d = go_10_goMux_data_onehotd[1];
  assign lizzieLet4_3QNode_Int_d = go_10_goMux_data_onehotd[2];
  assign lizzieLet4_3QError_Int_d = go_10_goMux_data_onehotd[3];
  assign go_10_goMux_data_r = (| (go_10_goMux_data_onehotd & {lizzieLet4_3QError_Int_r,
                                                              lizzieLet4_3QNode_Int_r,
                                                              lizzieLet4_3QVal_Int_r,
                                                              lizzieLet4_3QNone_Int_r}));
  assign lizzieLet4_3_r = go_10_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet4_3QError_Int,Go) > [(lizzieLet4_3QError_Int_1,Go),
                                              (lizzieLet4_3QError_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QError_Int_emitted;
  logic [1:0] lizzieLet4_3QError_Int_done;
  assign lizzieLet4_3QError_Int_1_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[0]));
  assign lizzieLet4_3QError_Int_2_d = (lizzieLet4_3QError_Int_d[0] && (! lizzieLet4_3QError_Int_emitted[1]));
  assign lizzieLet4_3QError_Int_done = (lizzieLet4_3QError_Int_emitted | ({lizzieLet4_3QError_Int_2_d[0],
                                                                           lizzieLet4_3QError_Int_1_d[0]} & {lizzieLet4_3QError_Int_2_r,
                                                                                                             lizzieLet4_3QError_Int_1_r}));
  assign lizzieLet4_3QError_Int_r = (& lizzieLet4_3QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QError_Int_emitted <= (lizzieLet4_3QError_Int_r ? 2'd0 :
                                         lizzieLet4_3QError_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_1,Go) > (lizzieLet4_3QError_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_1_bufchan_d;
  logic lizzieLet4_3QError_Int_1_bufchan_r;
  assign lizzieLet4_3QError_Int_1_r = ((! lizzieLet4_3QError_Int_1_bufchan_d[0]) || lizzieLet4_3QError_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_1_r)
        lizzieLet4_3QError_Int_1_bufchan_d <= lizzieLet4_3QError_Int_1_d;
  Go_t lizzieLet4_3QError_Int_1_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_bufchan_r = (! lizzieLet4_3QError_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_1_argbuf_d = (lizzieLet4_3QError_Int_1_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_bufchan_buf :
                                              lizzieLet4_3QError_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_1_argbuf_r && lizzieLet4_3QError_Int_1_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_bufchan_buf <= lizzieLet4_3QError_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QError_Int_1_argbuf,Go) > (lizzieLet4_3QError_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QError_Int_1_argbuf_0_d = {32'd0,
                                                lizzieLet4_3QError_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QError_Int_1_argbuf_r = lizzieLet4_3QError_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QError_Int_1_argbuf_0,Int#) > (lizzieLet11_1_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QError_Int_1_argbuf_0_r = ((! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QError_Int_1_argbuf_0_r)
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QError_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QError_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet11_1_1_argbuf_d = (lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf :
                                     lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet11_1_1_argbuf_r && lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet11_1_1_argbuf_r) && (! lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QError_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QError_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QError_Int_2,Go) > (lizzieLet4_3QError_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QError_Int_2_bufchan_d;
  logic lizzieLet4_3QError_Int_2_bufchan_r;
  assign lizzieLet4_3QError_Int_2_r = ((! lizzieLet4_3QError_Int_2_bufchan_d[0]) || lizzieLet4_3QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QError_Int_2_r)
        lizzieLet4_3QError_Int_2_bufchan_d <= lizzieLet4_3QError_Int_2_d;
  Go_t lizzieLet4_3QError_Int_2_bufchan_buf;
  assign lizzieLet4_3QError_Int_2_bufchan_r = (! lizzieLet4_3QError_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QError_Int_2_argbuf_d = (lizzieLet4_3QError_Int_2_bufchan_buf[0] ? lizzieLet4_3QError_Int_2_bufchan_buf :
                                              lizzieLet4_3QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QError_Int_2_argbuf_r && lizzieLet4_3QError_Int_2_bufchan_buf[0]))
        lizzieLet4_3QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QError_Int_2_argbuf_r) && (! lizzieLet4_3QError_Int_2_bufchan_buf[0])))
        lizzieLet4_3QError_Int_2_bufchan_buf <= lizzieLet4_3QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNode_Int,Go) > (lizzieLet4_3QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNode_Int_bufchan_d;
  logic lizzieLet4_3QNode_Int_bufchan_r;
  assign lizzieLet4_3QNode_Int_r = ((! lizzieLet4_3QNode_Int_bufchan_d[0]) || lizzieLet4_3QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNode_Int_r)
        lizzieLet4_3QNode_Int_bufchan_d <= lizzieLet4_3QNode_Int_d;
  Go_t lizzieLet4_3QNode_Int_bufchan_buf;
  assign lizzieLet4_3QNode_Int_bufchan_r = (! lizzieLet4_3QNode_Int_bufchan_buf[0]);
  assign lizzieLet4_3QNode_Int_1_argbuf_d = (lizzieLet4_3QNode_Int_bufchan_buf[0] ? lizzieLet4_3QNode_Int_bufchan_buf :
                                             lizzieLet4_3QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNode_Int_1_argbuf_r && lizzieLet4_3QNode_Int_bufchan_buf[0]))
        lizzieLet4_3QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNode_Int_1_argbuf_r) && (! lizzieLet4_3QNode_Int_bufchan_buf[0])))
        lizzieLet4_3QNode_Int_bufchan_buf <= lizzieLet4_3QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet4_3QNone_Int,Go) > [(lizzieLet4_3QNone_Int_1,Go),
                                             (lizzieLet4_3QNone_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QNone_Int_emitted;
  logic [1:0] lizzieLet4_3QNone_Int_done;
  assign lizzieLet4_3QNone_Int_1_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[0]));
  assign lizzieLet4_3QNone_Int_2_d = (lizzieLet4_3QNone_Int_d[0] && (! lizzieLet4_3QNone_Int_emitted[1]));
  assign lizzieLet4_3QNone_Int_done = (lizzieLet4_3QNone_Int_emitted | ({lizzieLet4_3QNone_Int_2_d[0],
                                                                         lizzieLet4_3QNone_Int_1_d[0]} & {lizzieLet4_3QNone_Int_2_r,
                                                                                                          lizzieLet4_3QNone_Int_1_r}));
  assign lizzieLet4_3QNone_Int_r = (& lizzieLet4_3QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QNone_Int_emitted <= (lizzieLet4_3QNone_Int_r ? 2'd0 :
                                        lizzieLet4_3QNone_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_1,Go) > (lizzieLet4_3QNone_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_1_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_r = ((! lizzieLet4_3QNone_Int_1_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_1_r)
        lizzieLet4_3QNone_Int_1_bufchan_d <= lizzieLet4_3QNone_Int_1_d;
  Go_t lizzieLet4_3QNone_Int_1_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_bufchan_r = (! lizzieLet4_3QNone_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_1_argbuf_d = (lizzieLet4_3QNone_Int_1_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_bufchan_buf :
                                             lizzieLet4_3QNone_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_1_argbuf_r && lizzieLet4_3QNone_Int_1_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_bufchan_buf <= lizzieLet4_3QNone_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 0) : (lizzieLet4_3QNone_Int_1_argbuf,Go) > (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) */
  assign lizzieLet4_3QNone_Int_1_argbuf_0_d = {32'd0,
                                               lizzieLet4_3QNone_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QNone_Int_1_argbuf_r = lizzieLet4_3QNone_Int_1_argbuf_0_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QNone_Int_1_argbuf_0,Int#) > (lizzieLet11_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  logic lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_r = ((! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d[0]) || lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QNone_Int_1_argbuf_0_r)
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d <= lizzieLet4_3QNone_Int_1_argbuf_0_d;
  \Int#_t  lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf;
  assign lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_r = (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]);
  assign lizzieLet11_1_argbuf_d = (lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0] ? lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf :
                                   lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet11_1_argbuf_r && lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet11_1_argbuf_r) && (! lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_buf <= lizzieLet4_3QNone_Int_1_argbuf_0_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QNone_Int_2,Go) > (lizzieLet4_3QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QNone_Int_2_bufchan_d;
  logic lizzieLet4_3QNone_Int_2_bufchan_r;
  assign lizzieLet4_3QNone_Int_2_r = ((! lizzieLet4_3QNone_Int_2_bufchan_d[0]) || lizzieLet4_3QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QNone_Int_2_r)
        lizzieLet4_3QNone_Int_2_bufchan_d <= lizzieLet4_3QNone_Int_2_d;
  Go_t lizzieLet4_3QNone_Int_2_bufchan_buf;
  assign lizzieLet4_3QNone_Int_2_bufchan_r = (! lizzieLet4_3QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QNone_Int_2_argbuf_d = (lizzieLet4_3QNone_Int_2_bufchan_buf[0] ? lizzieLet4_3QNone_Int_2_bufchan_buf :
                                             lizzieLet4_3QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QNone_Int_2_argbuf_r && lizzieLet4_3QNone_Int_2_bufchan_buf[0]))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QNone_Int_2_argbuf_r) && (! lizzieLet4_3QNone_Int_2_bufchan_buf[0])))
        lizzieLet4_3QNone_Int_2_bufchan_buf <= lizzieLet4_3QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C4,Ty Go) : [(lizzieLet4_3QNone_Int_2_argbuf,Go),
                           (lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf,Go),
                           (lizzieLet4_3QVal_Int_2_argbuf,Go),
                           (lizzieLet4_3QError_Int_2_argbuf,Go)] > (go_15_goMux_choice,C4) (go_15_goMux_data,Go) */
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_select_d = ((| lizzieLet4_3QNone_Int_2_argbuf_select_q) ? lizzieLet4_3QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet4_3QNone_Int_2_argbuf_d[0] ? 4'd1 :
                                                     (lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_d[0] ? 4'd2 :
                                                      (lizzieLet4_3QVal_Int_2_argbuf_d[0] ? 4'd4 :
                                                       (lizzieLet4_3QError_Int_2_argbuf_d[0] ? 4'd8 :
                                                        4'd0)))));
  logic [3:0] lizzieLet4_3QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= 4'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_select_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 4'd0 :
                                                  lizzieLet4_3QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet4_3QNone_Int_2_argbuf_emit_q <= (lizzieLet4_3QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet4_3QNone_Int_2_argbuf_emit_d;
  assign lizzieLet4_3QNone_Int_2_argbuf_emit_d = (lizzieLet4_3QNone_Int_2_argbuf_emit_q | ({go_15_goMux_choice_d[0],
                                                                                            go_15_goMux_data_d[0]} & {go_15_goMux_choice_r,
                                                                                                                      go_15_goMux_data_r}));
  logic lizzieLet4_3QNone_Int_2_argbuf_done;
  assign lizzieLet4_3QNone_Int_2_argbuf_done = (& lizzieLet4_3QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet4_3QError_Int_2_argbuf_r,
          lizzieLet4_3QVal_Int_2_argbuf_r,
          lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_r,
          lizzieLet4_3QNone_Int_2_argbuf_r} = (lizzieLet4_3QNone_Int_2_argbuf_done ? lizzieLet4_3QNone_Int_2_argbuf_select_d :
                                               4'd0);
  assign go_15_goMux_data_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QNone_Int_2_argbuf_d :
                               ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet19_3Lcall_$wnnz_Int0_1_argbuf_d :
                                ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QVal_Int_2_argbuf_d :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet4_3QError_Int_2_argbuf_d :
                                  1'd0))));
  assign go_15_goMux_choice_d = ((lizzieLet4_3QNone_Int_2_argbuf_select_d[0] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C1_4_dc(1'd1) :
                                 ((lizzieLet4_3QNone_Int_2_argbuf_select_d[1] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C2_4_dc(1'd1) :
                                  ((lizzieLet4_3QNone_Int_2_argbuf_select_d[2] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C3_4_dc(1'd1) :
                                   ((lizzieLet4_3QNone_Int_2_argbuf_select_d[3] && (! lizzieLet4_3QNone_Int_2_argbuf_emit_q[1])) ? C4_4_dc(1'd1) :
                                    {2'd0, 1'd0}))));
  
  /* fork (Ty Go) : (lizzieLet4_3QVal_Int,Go) > [(lizzieLet4_3QVal_Int_1,Go),
                                            (lizzieLet4_3QVal_Int_2,Go)] */
  logic [1:0] lizzieLet4_3QVal_Int_emitted;
  logic [1:0] lizzieLet4_3QVal_Int_done;
  assign lizzieLet4_3QVal_Int_1_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[0]));
  assign lizzieLet4_3QVal_Int_2_d = (lizzieLet4_3QVal_Int_d[0] && (! lizzieLet4_3QVal_Int_emitted[1]));
  assign lizzieLet4_3QVal_Int_done = (lizzieLet4_3QVal_Int_emitted | ({lizzieLet4_3QVal_Int_2_d[0],
                                                                       lizzieLet4_3QVal_Int_1_d[0]} & {lizzieLet4_3QVal_Int_2_r,
                                                                                                       lizzieLet4_3QVal_Int_1_r}));
  assign lizzieLet4_3QVal_Int_r = (& lizzieLet4_3QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_emitted <= 2'd0;
    else
      lizzieLet4_3QVal_Int_emitted <= (lizzieLet4_3QVal_Int_r ? 2'd0 :
                                       lizzieLet4_3QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_1,Go) > (lizzieLet4_3QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_r = ((! lizzieLet4_3QVal_Int_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_1_r)
        lizzieLet4_3QVal_Int_1_bufchan_d <= lizzieLet4_3QVal_Int_1_d;
  Go_t lizzieLet4_3QVal_Int_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_1_argbuf_d = (lizzieLet4_3QVal_Int_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_bufchan_buf :
                                            lizzieLet4_3QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_1_argbuf_r && lizzieLet4_3QVal_Int_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_bufchan_d;
  
  /* const (Ty Int#,
       Lit 1) : (lizzieLet4_3QVal_Int_1_argbuf,Go) > (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) */
  assign lizzieLet4_3QVal_Int_1_argbuf_1_d = {32'd1,
                                              lizzieLet4_3QVal_Int_1_argbuf_d[0]};
  assign lizzieLet4_3QVal_Int_1_argbuf_r = lizzieLet4_3QVal_Int_1_argbuf_1_r;
  
  /* buf (Ty Int#) : (lizzieLet4_3QVal_Int_1_argbuf_1,Int#) > (lizzieLet12_1_argbuf,Int#) */
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  logic lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_r = ((! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d[0]) || lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet4_3QVal_Int_1_argbuf_1_r)
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d <= lizzieLet4_3QVal_Int_1_argbuf_1_d;
  \Int#_t  lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf;
  assign lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_r = (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]);
  assign lizzieLet12_1_argbuf_d = (lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0] ? lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf :
                                   lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet12_1_argbuf_r && lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet12_1_argbuf_r) && (! lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_buf <= lizzieLet4_3QVal_Int_1_argbuf_1_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet4_3QVal_Int_2,Go) > (lizzieLet4_3QVal_Int_2_argbuf,Go) */
  Go_t lizzieLet4_3QVal_Int_2_bufchan_d;
  logic lizzieLet4_3QVal_Int_2_bufchan_r;
  assign lizzieLet4_3QVal_Int_2_r = ((! lizzieLet4_3QVal_Int_2_bufchan_d[0]) || lizzieLet4_3QVal_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet4_3QVal_Int_2_r)
        lizzieLet4_3QVal_Int_2_bufchan_d <= lizzieLet4_3QVal_Int_2_d;
  Go_t lizzieLet4_3QVal_Int_2_bufchan_buf;
  assign lizzieLet4_3QVal_Int_2_bufchan_r = (! lizzieLet4_3QVal_Int_2_bufchan_buf[0]);
  assign lizzieLet4_3QVal_Int_2_argbuf_d = (lizzieLet4_3QVal_Int_2_bufchan_buf[0] ? lizzieLet4_3QVal_Int_2_bufchan_buf :
                                            lizzieLet4_3QVal_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet4_3QVal_Int_2_argbuf_r && lizzieLet4_3QVal_Int_2_bufchan_buf[0]))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet4_3QVal_Int_2_argbuf_r) && (! lizzieLet4_3QVal_Int_2_bufchan_buf[0])))
        lizzieLet4_3QVal_Int_2_bufchan_buf <= lizzieLet4_3QVal_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4,QTree_Int) (sc_0_goMux_mux,Pointer_CT$wnnz_Int) > [(lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                                                                                  (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int)] */
  logic [3:0] sc_0_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet4_4_d[0] && sc_0_goMux_mux_d[0]))
      unique case (lizzieLet4_4_d[2:1])
        2'd0: sc_0_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_goMux_mux_onehotd = 4'd8;
        default: sc_0_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_goMux_mux_onehotd = 4'd0;
  assign lizzieLet4_4QNone_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[0]};
  assign lizzieLet4_4QVal_Int_d = {sc_0_goMux_mux_d[16:1],
                                   sc_0_goMux_mux_onehotd[1]};
  assign lizzieLet4_4QNode_Int_d = {sc_0_goMux_mux_d[16:1],
                                    sc_0_goMux_mux_onehotd[2]};
  assign lizzieLet4_4QError_Int_d = {sc_0_goMux_mux_d[16:1],
                                     sc_0_goMux_mux_onehotd[3]};
  assign sc_0_goMux_mux_r = (| (sc_0_goMux_mux_onehotd & {lizzieLet4_4QError_Int_r,
                                                          lizzieLet4_4QNode_Int_r,
                                                          lizzieLet4_4QVal_Int_r,
                                                          lizzieLet4_4QNone_Int_r}));
  assign lizzieLet4_4_r = sc_0_goMux_mux_r;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QError_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QError_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_d;
  logic lizzieLet4_4QError_Int_bufchan_r;
  assign lizzieLet4_4QError_Int_r = ((! lizzieLet4_4QError_Int_bufchan_d[0]) || lizzieLet4_4QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QError_Int_r)
        lizzieLet4_4QError_Int_bufchan_d <= lizzieLet4_4QError_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QError_Int_bufchan_buf;
  assign lizzieLet4_4QError_Int_bufchan_r = (! lizzieLet4_4QError_Int_bufchan_buf[0]);
  assign lizzieLet4_4QError_Int_1_argbuf_d = (lizzieLet4_4QError_Int_bufchan_buf[0] ? lizzieLet4_4QError_Int_bufchan_buf :
                                              lizzieLet4_4QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QError_Int_1_argbuf_r && lizzieLet4_4QError_Int_bufchan_buf[0]))
        lizzieLet4_4QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QError_Int_1_argbuf_r) && (! lizzieLet4_4QError_Int_bufchan_buf[0])))
        lizzieLet4_4QError_Int_bufchan_buf <= lizzieLet4_4QError_Int_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int3) : [(lizzieLet4_4QNode_Int,Pointer_CT$wnnz_Int),
                                (q4abZ_destruct,Pointer_QTree_Int),
                                (q3abY_destruct,Pointer_QTree_Int),
                                (q2abX_destruct,Pointer_QTree_Int)] > (lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3,CT$wnnz_Int) */
  assign lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_d = Lcall_$wnnz_Int3_dc((& {lizzieLet4_4QNode_Int_d[0],
                                                                                                  q4abZ_destruct_d[0],
                                                                                                  q3abY_destruct_d[0],
                                                                                                  q2abX_destruct_d[0]}), lizzieLet4_4QNode_Int_d, q4abZ_destruct_d, q3abY_destruct_d, q2abX_destruct_d);
  assign {lizzieLet4_4QNode_Int_r,
          q4abZ_destruct_r,
          q3abY_destruct_r,
          q2abX_destruct_r} = {4 {(lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_r && lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3,CT$wnnz_Int) > (lizzieLet5_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d;
  logic lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_r;
  assign lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_r = ((! lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d[0]) || lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d <= {115'd0,
                                                                                 1'd0};
    else
      if (lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_r)
        lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d <= lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_d;
  CT$wnnz_Int_t lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf;
  assign lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_r = (! lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf[0]);
  assign lizzieLet5_1_argbuf_d = (lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf[0] ? lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf :
                                  lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                   1'd0};
    else
      if ((lizzieLet5_1_argbuf_r && lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf[0]))
        lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf <= {115'd0,
                                                                                     1'd0};
      else if (((! lizzieLet5_1_argbuf_r) && (! lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf[0])))
        lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_buf <= lizzieLet4_4QNode_Int_1q4abZ_1q3abY_1q2abX_1Lcall_$wnnz_Int3_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QNone_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QNone_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_d;
  logic lizzieLet4_4QNone_Int_bufchan_r;
  assign lizzieLet4_4QNone_Int_r = ((! lizzieLet4_4QNone_Int_bufchan_d[0]) || lizzieLet4_4QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QNone_Int_r)
        lizzieLet4_4QNone_Int_bufchan_d <= lizzieLet4_4QNone_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QNone_Int_bufchan_buf;
  assign lizzieLet4_4QNone_Int_bufchan_r = (! lizzieLet4_4QNone_Int_bufchan_buf[0]);
  assign lizzieLet4_4QNone_Int_1_argbuf_d = (lizzieLet4_4QNone_Int_bufchan_buf[0] ? lizzieLet4_4QNone_Int_bufchan_buf :
                                             lizzieLet4_4QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QNone_Int_1_argbuf_r && lizzieLet4_4QNone_Int_bufchan_buf[0]))
        lizzieLet4_4QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QNone_Int_1_argbuf_r) && (! lizzieLet4_4QNone_Int_bufchan_buf[0])))
        lizzieLet4_4QNone_Int_bufchan_buf <= lizzieLet4_4QNone_Int_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (lizzieLet4_4QVal_Int,Pointer_CT$wnnz_Int) > (lizzieLet4_4QVal_Int_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_d;
  logic lizzieLet4_4QVal_Int_bufchan_r;
  assign lizzieLet4_4QVal_Int_r = ((! lizzieLet4_4QVal_Int_bufchan_d[0]) || lizzieLet4_4QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet4_4QVal_Int_r)
        lizzieLet4_4QVal_Int_bufchan_d <= lizzieLet4_4QVal_Int_d;
  Pointer_CT$wnnz_Int_t lizzieLet4_4QVal_Int_bufchan_buf;
  assign lizzieLet4_4QVal_Int_bufchan_r = (! lizzieLet4_4QVal_Int_bufchan_buf[0]);
  assign lizzieLet4_4QVal_Int_1_argbuf_d = (lizzieLet4_4QVal_Int_bufchan_buf[0] ? lizzieLet4_4QVal_Int_bufchan_buf :
                                            lizzieLet4_4QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet4_4QVal_Int_1_argbuf_r && lizzieLet4_4QVal_Int_bufchan_buf[0]))
        lizzieLet4_4QVal_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet4_4QVal_Int_1_argbuf_r) && (! lizzieLet4_4QVal_Int_bufchan_buf[0])))
        lizzieLet4_4QVal_Int_bufchan_buf <= lizzieLet4_4QVal_Int_bufchan_d;
  
  /* destruct (Ty QTree_Int,
          Dcon QNode_Int) : (lizzieLet6_1QNode_Int,QTree_Int) > [(q1aic_destruct,Pointer_QTree_Int),
                                                                 (q2aid_destruct,Pointer_QTree_Int),
                                                                 (q3aie_destruct,Pointer_QTree_Int),
                                                                 (q4aif_destruct,Pointer_QTree_Int)] */
  logic [3:0] lizzieLet6_1QNode_Int_emitted;
  logic [3:0] lizzieLet6_1QNode_Int_done;
  assign q1aic_destruct_d = {lizzieLet6_1QNode_Int_d[18:3],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[0]))};
  assign q2aid_destruct_d = {lizzieLet6_1QNode_Int_d[34:19],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[1]))};
  assign q3aie_destruct_d = {lizzieLet6_1QNode_Int_d[50:35],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[2]))};
  assign q4aif_destruct_d = {lizzieLet6_1QNode_Int_d[66:51],
                             (lizzieLet6_1QNode_Int_d[0] && (! lizzieLet6_1QNode_Int_emitted[3]))};
  assign lizzieLet6_1QNode_Int_done = (lizzieLet6_1QNode_Int_emitted | ({q4aif_destruct_d[0],
                                                                         q3aie_destruct_d[0],
                                                                         q2aid_destruct_d[0],
                                                                         q1aic_destruct_d[0]} & {q4aif_destruct_r,
                                                                                                 q3aie_destruct_r,
                                                                                                 q2aid_destruct_r,
                                                                                                 q1aic_destruct_r}));
  assign lizzieLet6_1QNode_Int_r = (& lizzieLet6_1QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_1QNode_Int_emitted <= 4'd0;
    else
      lizzieLet6_1QNode_Int_emitted <= (lizzieLet6_1QNode_Int_r ? 4'd0 :
                                        lizzieLet6_1QNode_Int_done);
  
  /* destruct (Ty QTree_Int,
          Dcon QVal_Int) : (lizzieLet6_1QVal_Int,QTree_Int) > [(v'aib_destruct,Int)] */
  assign \v'aib_destruct_d  = {lizzieLet6_1QVal_Int_d[34:3],
                               lizzieLet6_1QVal_Int_d[0]};
  assign lizzieLet6_1QVal_Int_r = \v'aib_destruct_r ;
  
  /* demux (Ty QTree_Int,
       Ty QTree_Int) : (lizzieLet6_2,QTree_Int) (lizzieLet6_1,QTree_Int) > [(_11,QTree_Int),
                                                                            (lizzieLet6_1QVal_Int,QTree_Int),
                                                                            (lizzieLet6_1QNode_Int,QTree_Int),
                                                                            (_10,QTree_Int)] */
  logic [3:0] lizzieLet6_1_onehotd;
  always_comb
    if ((lizzieLet6_2_d[0] && lizzieLet6_1_d[0]))
      unique case (lizzieLet6_2_d[2:1])
        2'd0: lizzieLet6_1_onehotd = 4'd1;
        2'd1: lizzieLet6_1_onehotd = 4'd2;
        2'd2: lizzieLet6_1_onehotd = 4'd4;
        2'd3: lizzieLet6_1_onehotd = 4'd8;
        default: lizzieLet6_1_onehotd = 4'd0;
      endcase
    else lizzieLet6_1_onehotd = 4'd0;
  assign _11_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[0]};
  assign lizzieLet6_1QVal_Int_d = {lizzieLet6_1_d[66:1],
                                   lizzieLet6_1_onehotd[1]};
  assign lizzieLet6_1QNode_Int_d = {lizzieLet6_1_d[66:1],
                                    lizzieLet6_1_onehotd[2]};
  assign _10_d = {lizzieLet6_1_d[66:1], lizzieLet6_1_onehotd[3]};
  assign lizzieLet6_1_r = (| (lizzieLet6_1_onehotd & {_10_r,
                                                      lizzieLet6_1QNode_Int_r,
                                                      lizzieLet6_1QVal_Int_r,
                                                      _11_r}));
  assign lizzieLet6_2_r = lizzieLet6_1_r;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int) : (lizzieLet6_3,QTree_Int) (f_mapaia_goMux_mux,MyDTInt_Int) > [(_9,MyDTInt_Int),
                                                                                      (lizzieLet6_3QVal_Int,MyDTInt_Int),
                                                                                      (lizzieLet6_3QNode_Int,MyDTInt_Int),
                                                                                      (_8,MyDTInt_Int)] */
  logic [3:0] f_mapaia_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_3_d[0] && f_mapaia_goMux_mux_d[0]))
      unique case (lizzieLet6_3_d[2:1])
        2'd0: f_mapaia_goMux_mux_onehotd = 4'd1;
        2'd1: f_mapaia_goMux_mux_onehotd = 4'd2;
        2'd2: f_mapaia_goMux_mux_onehotd = 4'd4;
        2'd3: f_mapaia_goMux_mux_onehotd = 4'd8;
        default: f_mapaia_goMux_mux_onehotd = 4'd0;
      endcase
    else f_mapaia_goMux_mux_onehotd = 4'd0;
  assign _9_d = f_mapaia_goMux_mux_onehotd[0];
  assign lizzieLet6_3QVal_Int_d = f_mapaia_goMux_mux_onehotd[1];
  assign lizzieLet6_3QNode_Int_d = f_mapaia_goMux_mux_onehotd[2];
  assign _8_d = f_mapaia_goMux_mux_onehotd[3];
  assign f_mapaia_goMux_mux_r = (| (f_mapaia_goMux_mux_onehotd & {_8_r,
                                                                  lizzieLet6_3QNode_Int_r,
                                                                  lizzieLet6_3QVal_Int_r,
                                                                  _9_r}));
  assign lizzieLet6_3_r = f_mapaia_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int) : (lizzieLet6_3QNode_Int,MyDTInt_Int) > [(lizzieLet6_3QNode_Int_1,MyDTInt_Int),
                                                               (lizzieLet6_3QNode_Int_2,MyDTInt_Int)] */
  logic [1:0] lizzieLet6_3QNode_Int_emitted;
  logic [1:0] lizzieLet6_3QNode_Int_done;
  assign lizzieLet6_3QNode_Int_1_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[0]));
  assign lizzieLet6_3QNode_Int_2_d = (lizzieLet6_3QNode_Int_d[0] && (! lizzieLet6_3QNode_Int_emitted[1]));
  assign lizzieLet6_3QNode_Int_done = (lizzieLet6_3QNode_Int_emitted | ({lizzieLet6_3QNode_Int_2_d[0],
                                                                         lizzieLet6_3QNode_Int_1_d[0]} & {lizzieLet6_3QNode_Int_2_r,
                                                                                                          lizzieLet6_3QNode_Int_1_r}));
  assign lizzieLet6_3QNode_Int_r = (& lizzieLet6_3QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_3QNode_Int_emitted <= (lizzieLet6_3QNode_Int_r ? 2'd0 :
                                        lizzieLet6_3QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int) : (lizzieLet6_3QNode_Int_2,MyDTInt_Int) > (lizzieLet6_3QNode_Int_2_argbuf,MyDTInt_Int) */
  MyDTInt_Int_t lizzieLet6_3QNode_Int_2_bufchan_d;
  logic lizzieLet6_3QNode_Int_2_bufchan_r;
  assign lizzieLet6_3QNode_Int_2_r = ((! lizzieLet6_3QNode_Int_2_bufchan_d[0]) || lizzieLet6_3QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_3QNode_Int_2_r)
        lizzieLet6_3QNode_Int_2_bufchan_d <= lizzieLet6_3QNode_Int_2_d;
  MyDTInt_Int_t lizzieLet6_3QNode_Int_2_bufchan_buf;
  assign lizzieLet6_3QNode_Int_2_bufchan_r = (! lizzieLet6_3QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_3QNode_Int_2_argbuf_d = (lizzieLet6_3QNode_Int_2_bufchan_buf[0] ? lizzieLet6_3QNode_Int_2_bufchan_buf :
                                             lizzieLet6_3QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_3QNode_Int_2_argbuf_r && lizzieLet6_3QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_3QNode_Int_2_argbuf_r) && (! lizzieLet6_3QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_3QNode_Int_2_bufchan_buf <= lizzieLet6_3QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Go) : (lizzieLet6_4,QTree_Int) (go_11_goMux_data,Go) > [(lizzieLet6_4QNone_Int,Go),
                                                                  (lizzieLet6_4QVal_Int,Go),
                                                                  (lizzieLet6_4QNode_Int,Go),
                                                                  (lizzieLet6_4QError_Int,Go)] */
  logic [3:0] go_11_goMux_data_onehotd;
  always_comb
    if ((lizzieLet6_4_d[0] && go_11_goMux_data_d[0]))
      unique case (lizzieLet6_4_d[2:1])
        2'd0: go_11_goMux_data_onehotd = 4'd1;
        2'd1: go_11_goMux_data_onehotd = 4'd2;
        2'd2: go_11_goMux_data_onehotd = 4'd4;
        2'd3: go_11_goMux_data_onehotd = 4'd8;
        default: go_11_goMux_data_onehotd = 4'd0;
      endcase
    else go_11_goMux_data_onehotd = 4'd0;
  assign lizzieLet6_4QNone_Int_d = go_11_goMux_data_onehotd[0];
  assign lizzieLet6_4QVal_Int_d = go_11_goMux_data_onehotd[1];
  assign lizzieLet6_4QNode_Int_d = go_11_goMux_data_onehotd[2];
  assign lizzieLet6_4QError_Int_d = go_11_goMux_data_onehotd[3];
  assign go_11_goMux_data_r = (| (go_11_goMux_data_onehotd & {lizzieLet6_4QError_Int_r,
                                                              lizzieLet6_4QNode_Int_r,
                                                              lizzieLet6_4QVal_Int_r,
                                                              lizzieLet6_4QNone_Int_r}));
  assign lizzieLet6_4_r = go_11_goMux_data_r;
  
  /* fork (Ty Go) : (lizzieLet6_4QError_Int,Go) > [(lizzieLet6_4QError_Int_1,Go),
                                              (lizzieLet6_4QError_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QError_Int_emitted;
  logic [1:0] lizzieLet6_4QError_Int_done;
  assign lizzieLet6_4QError_Int_1_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[0]));
  assign lizzieLet6_4QError_Int_2_d = (lizzieLet6_4QError_Int_d[0] && (! lizzieLet6_4QError_Int_emitted[1]));
  assign lizzieLet6_4QError_Int_done = (lizzieLet6_4QError_Int_emitted | ({lizzieLet6_4QError_Int_2_d[0],
                                                                           lizzieLet6_4QError_Int_1_d[0]} & {lizzieLet6_4QError_Int_2_r,
                                                                                                             lizzieLet6_4QError_Int_1_r}));
  assign lizzieLet6_4QError_Int_r = (& lizzieLet6_4QError_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QError_Int_emitted <= (lizzieLet6_4QError_Int_r ? 2'd0 :
                                         lizzieLet6_4QError_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QError_Int) : [(lizzieLet6_4QError_Int_1,Go)] > (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) */
  assign lizzieLet6_4QError_Int_1QError_Int_d = QError_Int_dc((& {lizzieLet6_4QError_Int_1_d[0]}), lizzieLet6_4QError_Int_1_d);
  assign {lizzieLet6_4QError_Int_1_r} = {1 {(lizzieLet6_4QError_Int_1QError_Int_r && lizzieLet6_4QError_Int_1QError_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QError_Int_1QError_Int,QTree_Int) > (lizzieLet12_1_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  logic lizzieLet6_4QError_Int_1QError_Int_bufchan_r;
  assign lizzieLet6_4QError_Int_1QError_Int_r = ((! lizzieLet6_4QError_Int_1QError_Int_bufchan_d[0]) || lizzieLet6_4QError_Int_1QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QError_Int_1QError_Int_r)
        lizzieLet6_4QError_Int_1QError_Int_bufchan_d <= lizzieLet6_4QError_Int_1QError_Int_d;
  QTree_Int_t lizzieLet6_4QError_Int_1QError_Int_bufchan_buf;
  assign lizzieLet6_4QError_Int_1QError_Int_bufchan_r = (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]);
  assign lizzieLet12_1_1_argbuf_d = (lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0] ? lizzieLet6_4QError_Int_1QError_Int_bufchan_buf :
                                     lizzieLet6_4QError_Int_1QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet12_1_1_argbuf_r && lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0]))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet12_1_1_argbuf_r) && (! lizzieLet6_4QError_Int_1QError_Int_bufchan_buf[0])))
        lizzieLet6_4QError_Int_1QError_Int_bufchan_buf <= lizzieLet6_4QError_Int_1QError_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QError_Int_2,Go) > (lizzieLet6_4QError_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QError_Int_2_bufchan_d;
  logic lizzieLet6_4QError_Int_2_bufchan_r;
  assign lizzieLet6_4QError_Int_2_r = ((! lizzieLet6_4QError_Int_2_bufchan_d[0]) || lizzieLet6_4QError_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QError_Int_2_r)
        lizzieLet6_4QError_Int_2_bufchan_d <= lizzieLet6_4QError_Int_2_d;
  Go_t lizzieLet6_4QError_Int_2_bufchan_buf;
  assign lizzieLet6_4QError_Int_2_bufchan_r = (! lizzieLet6_4QError_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QError_Int_2_argbuf_d = (lizzieLet6_4QError_Int_2_bufchan_buf[0] ? lizzieLet6_4QError_Int_2_bufchan_buf :
                                              lizzieLet6_4QError_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QError_Int_2_argbuf_r && lizzieLet6_4QError_Int_2_bufchan_buf[0]))
        lizzieLet6_4QError_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QError_Int_2_argbuf_r) && (! lizzieLet6_4QError_Int_2_bufchan_buf[0])))
        lizzieLet6_4QError_Int_2_bufchan_buf <= lizzieLet6_4QError_Int_2_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNode_Int,Go) > (lizzieLet6_4QNode_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QNode_Int_bufchan_d;
  logic lizzieLet6_4QNode_Int_bufchan_r;
  assign lizzieLet6_4QNode_Int_r = ((! lizzieLet6_4QNode_Int_bufchan_d[0]) || lizzieLet6_4QNode_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNode_Int_r)
        lizzieLet6_4QNode_Int_bufchan_d <= lizzieLet6_4QNode_Int_d;
  Go_t lizzieLet6_4QNode_Int_bufchan_buf;
  assign lizzieLet6_4QNode_Int_bufchan_r = (! lizzieLet6_4QNode_Int_bufchan_buf[0]);
  assign lizzieLet6_4QNode_Int_1_argbuf_d = (lizzieLet6_4QNode_Int_bufchan_buf[0] ? lizzieLet6_4QNode_Int_bufchan_buf :
                                             lizzieLet6_4QNode_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNode_Int_1_argbuf_r && lizzieLet6_4QNode_Int_bufchan_buf[0]))
        lizzieLet6_4QNode_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNode_Int_1_argbuf_r) && (! lizzieLet6_4QNode_Int_bufchan_buf[0])))
        lizzieLet6_4QNode_Int_bufchan_buf <= lizzieLet6_4QNode_Int_bufchan_d;
  
  /* fork (Ty Go) : (lizzieLet6_4QNone_Int,Go) > [(lizzieLet6_4QNone_Int_1,Go),
                                             (lizzieLet6_4QNone_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QNone_Int_emitted;
  logic [1:0] lizzieLet6_4QNone_Int_done;
  assign lizzieLet6_4QNone_Int_1_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[0]));
  assign lizzieLet6_4QNone_Int_2_d = (lizzieLet6_4QNone_Int_d[0] && (! lizzieLet6_4QNone_Int_emitted[1]));
  assign lizzieLet6_4QNone_Int_done = (lizzieLet6_4QNone_Int_emitted | ({lizzieLet6_4QNone_Int_2_d[0],
                                                                         lizzieLet6_4QNone_Int_1_d[0]} & {lizzieLet6_4QNone_Int_2_r,
                                                                                                          lizzieLet6_4QNone_Int_1_r}));
  assign lizzieLet6_4QNone_Int_r = (& lizzieLet6_4QNone_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QNone_Int_emitted <= (lizzieLet6_4QNone_Int_r ? 2'd0 :
                                        lizzieLet6_4QNone_Int_done);
  
  /* dcon (Ty QTree_Int,
      Dcon QNone_Int) : [(lizzieLet6_4QNone_Int_1,Go)] > (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) */
  assign lizzieLet6_4QNone_Int_1QNone_Int_d = QNone_Int_dc((& {lizzieLet6_4QNone_Int_1_d[0]}), lizzieLet6_4QNone_Int_1_d);
  assign {lizzieLet6_4QNone_Int_1_r} = {1 {(lizzieLet6_4QNone_Int_1QNone_Int_r && lizzieLet6_4QNone_Int_1QNone_Int_d[0])}};
  
  /* buf (Ty QTree_Int) : (lizzieLet6_4QNone_Int_1QNone_Int,QTree_Int) > (lizzieLet7_1_argbuf,QTree_Int) */
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  logic lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r;
  assign lizzieLet6_4QNone_Int_1QNone_Int_r = ((! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d[0]) || lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= {66'd0, 1'd0};
    else
      if (lizzieLet6_4QNone_Int_1QNone_Int_r)
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d <= lizzieLet6_4QNone_Int_1QNone_Int_d;
  QTree_Int_t lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf;
  assign lizzieLet6_4QNone_Int_1QNone_Int_bufchan_r = (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]);
  assign lizzieLet7_1_argbuf_d = (lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0] ? lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf :
                                  lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((lizzieLet7_1_argbuf_r && lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= {66'd0, 1'd0};
      else if (((! lizzieLet7_1_argbuf_r) && (! lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_1QNone_Int_bufchan_buf <= lizzieLet6_4QNone_Int_1QNone_Int_bufchan_d;
  
  /* buf (Ty Go) : (lizzieLet6_4QNone_Int_2,Go) > (lizzieLet6_4QNone_Int_2_argbuf,Go) */
  Go_t lizzieLet6_4QNone_Int_2_bufchan_d;
  logic lizzieLet6_4QNone_Int_2_bufchan_r;
  assign lizzieLet6_4QNone_Int_2_r = ((! lizzieLet6_4QNone_Int_2_bufchan_d[0]) || lizzieLet6_4QNone_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QNone_Int_2_r)
        lizzieLet6_4QNone_Int_2_bufchan_d <= lizzieLet6_4QNone_Int_2_d;
  Go_t lizzieLet6_4QNone_Int_2_bufchan_buf;
  assign lizzieLet6_4QNone_Int_2_bufchan_r = (! lizzieLet6_4QNone_Int_2_bufchan_buf[0]);
  assign lizzieLet6_4QNone_Int_2_argbuf_d = (lizzieLet6_4QNone_Int_2_bufchan_buf[0] ? lizzieLet6_4QNone_Int_2_bufchan_buf :
                                             lizzieLet6_4QNone_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QNone_Int_2_argbuf_r && lizzieLet6_4QNone_Int_2_bufchan_buf[0]))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QNone_Int_2_argbuf_r) && (! lizzieLet6_4QNone_Int_2_bufchan_buf[0])))
        lizzieLet6_4QNone_Int_2_bufchan_buf <= lizzieLet6_4QNone_Int_2_bufchan_d;
  
  /* mergectrl (Ty C6,Ty Go) : [(lizzieLet6_4QNone_Int_2_argbuf,Go),
                           (lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf,Go),
                           (es_7_1_2MyFalse_2_argbuf,Go),
                           (es_7_1_2MyTrue_2_argbuf,Go),
                           (es_2_2MyTrue_2_argbuf,Go),
                           (lizzieLet6_4QError_Int_2_argbuf,Go)] > (go_16_goMux_choice,C6) (go_16_goMux_data,Go) */
  logic [5:0] lizzieLet6_4QNone_Int_2_argbuf_select_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_select_d = ((| lizzieLet6_4QNone_Int_2_argbuf_select_q) ? lizzieLet6_4QNone_Int_2_argbuf_select_q :
                                                    (lizzieLet6_4QNone_Int_2_argbuf_d[0] ? 6'd1 :
                                                     (\lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_d [0] ? 6'd2 :
                                                      (es_7_1_2MyFalse_2_argbuf_d[0] ? 6'd4 :
                                                       (es_7_1_2MyTrue_2_argbuf_d[0] ? 6'd8 :
                                                        (es_2_2MyTrue_2_argbuf_d[0] ? 6'd16 :
                                                         (lizzieLet6_4QError_Int_2_argbuf_d[0] ? 6'd32 :
                                                          6'd0)))))));
  logic [5:0] lizzieLet6_4QNone_Int_2_argbuf_select_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= 6'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_select_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 6'd0 :
                                                  lizzieLet6_4QNone_Int_2_argbuf_select_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_q;
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QNone_Int_2_argbuf_emit_q <= 2'd0;
    else
      lizzieLet6_4QNone_Int_2_argbuf_emit_q <= (lizzieLet6_4QNone_Int_2_argbuf_done ? 2'd0 :
                                                lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  logic [1:0] lizzieLet6_4QNone_Int_2_argbuf_emit_d;
  assign lizzieLet6_4QNone_Int_2_argbuf_emit_d = (lizzieLet6_4QNone_Int_2_argbuf_emit_q | ({go_16_goMux_choice_d[0],
                                                                                            go_16_goMux_data_d[0]} & {go_16_goMux_choice_r,
                                                                                                                      go_16_goMux_data_r}));
  logic lizzieLet6_4QNone_Int_2_argbuf_done;
  assign lizzieLet6_4QNone_Int_2_argbuf_done = (& lizzieLet6_4QNone_Int_2_argbuf_emit_d);
  assign {lizzieLet6_4QError_Int_2_argbuf_r,
          es_2_2MyTrue_2_argbuf_r,
          es_7_1_2MyTrue_2_argbuf_r,
          es_7_1_2MyFalse_2_argbuf_r,
          \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_r ,
          lizzieLet6_4QNone_Int_2_argbuf_r} = (lizzieLet6_4QNone_Int_2_argbuf_done ? lizzieLet6_4QNone_Int_2_argbuf_select_d :
                                               6'd0);
  assign go_16_goMux_data_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QNone_Int_2_argbuf_d :
                               ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? \lizzieLet23_3Lcall_f'_f'_Int_Int_Int_Int0_1_argbuf_d  :
                                ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? es_7_1_2MyFalse_2_argbuf_d :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? es_7_1_2MyTrue_2_argbuf_d :
                                  ((lizzieLet6_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? es_2_2MyTrue_2_argbuf_d :
                                   ((lizzieLet6_4QNone_Int_2_argbuf_select_d[5] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[0])) ? lizzieLet6_4QError_Int_2_argbuf_d :
                                    1'd0))))));
  assign go_16_goMux_choice_d = ((lizzieLet6_4QNone_Int_2_argbuf_select_d[0] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C1_6_dc(1'd1) :
                                 ((lizzieLet6_4QNone_Int_2_argbuf_select_d[1] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C2_6_dc(1'd1) :
                                  ((lizzieLet6_4QNone_Int_2_argbuf_select_d[2] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C3_6_dc(1'd1) :
                                   ((lizzieLet6_4QNone_Int_2_argbuf_select_d[3] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C4_6_dc(1'd1) :
                                    ((lizzieLet6_4QNone_Int_2_argbuf_select_d[4] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C5_6_dc(1'd1) :
                                     ((lizzieLet6_4QNone_Int_2_argbuf_select_d[5] && (! lizzieLet6_4QNone_Int_2_argbuf_emit_q[1])) ? C6_6_dc(1'd1) :
                                      {3'd0, 1'd0}))))));
  
  /* fork (Ty Go) : (lizzieLet6_4QVal_Int,Go) > [(lizzieLet6_4QVal_Int_1,Go),
                                            (lizzieLet6_4QVal_Int_2,Go)] */
  logic [1:0] lizzieLet6_4QVal_Int_emitted;
  logic [1:0] lizzieLet6_4QVal_Int_done;
  assign lizzieLet6_4QVal_Int_1_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[0]));
  assign lizzieLet6_4QVal_Int_2_d = (lizzieLet6_4QVal_Int_d[0] && (! lizzieLet6_4QVal_Int_emitted[1]));
  assign lizzieLet6_4QVal_Int_done = (lizzieLet6_4QVal_Int_emitted | ({lizzieLet6_4QVal_Int_2_d[0],
                                                                       lizzieLet6_4QVal_Int_1_d[0]} & {lizzieLet6_4QVal_Int_2_r,
                                                                                                       lizzieLet6_4QVal_Int_1_r}));
  assign lizzieLet6_4QVal_Int_r = (& lizzieLet6_4QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_4QVal_Int_emitted <= (lizzieLet6_4QVal_Int_r ? 2'd0 :
                                       lizzieLet6_4QVal_Int_done);
  
  /* buf (Ty Go) : (lizzieLet6_4QVal_Int_1,Go) > (lizzieLet6_4QVal_Int_1_argbuf,Go) */
  Go_t lizzieLet6_4QVal_Int_1_bufchan_d;
  logic lizzieLet6_4QVal_Int_1_bufchan_r;
  assign lizzieLet6_4QVal_Int_1_r = ((! lizzieLet6_4QVal_Int_1_bufchan_d[0]) || lizzieLet6_4QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_4QVal_Int_1_r)
        lizzieLet6_4QVal_Int_1_bufchan_d <= lizzieLet6_4QVal_Int_1_d;
  Go_t lizzieLet6_4QVal_Int_1_bufchan_buf;
  assign lizzieLet6_4QVal_Int_1_bufchan_r = (! lizzieLet6_4QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_4QVal_Int_1_argbuf_d = (lizzieLet6_4QVal_Int_1_bufchan_buf[0] ? lizzieLet6_4QVal_Int_1_bufchan_buf :
                                            lizzieLet6_4QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_4QVal_Int_1_argbuf_r && lizzieLet6_4QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_4QVal_Int_1_argbuf_r) && (! lizzieLet6_4QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_4QVal_Int_1_bufchan_buf <= lizzieLet6_4QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupGo___MyDTInt_Bool___Int,
      Dcon TupGo___MyDTInt_Bool___Int) : [(lizzieLet6_4QVal_Int_1_argbuf,Go),
                                          (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool),
                                          (es_1_1_argbuf,Int)] > (applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1,TupGo___MyDTInt_Bool___Int) */
  assign applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d = TupGo___MyDTInt_Bool___Int_dc((& {lizzieLet6_4QVal_Int_1_argbuf_d[0],
                                                                                             lizzieLet6_5QVal_Int_1_argbuf_d[0],
                                                                                             es_1_1_argbuf_d[0]}), lizzieLet6_4QVal_Int_1_argbuf_d, lizzieLet6_5QVal_Int_1_argbuf_d, es_1_1_argbuf_d);
  assign {lizzieLet6_4QVal_Int_1_argbuf_r,
          lizzieLet6_5QVal_Int_1_argbuf_r,
          es_1_1_argbuf_r} = {3 {(applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_r && applyfnInt_Bool_5TupGo___MyDTInt_Bool___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_5,QTree_Int) (is_z_kronai6_goMux_mux,MyDTInt_Bool) > [(_7,MyDTInt_Bool),
                                                                                            (lizzieLet6_5QVal_Int,MyDTInt_Bool),
                                                                                            (lizzieLet6_5QNode_Int,MyDTInt_Bool),
                                                                                            (_6,MyDTInt_Bool)] */
  logic [3:0] is_z_kronai6_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_5_d[0] && is_z_kronai6_goMux_mux_d[0]))
      unique case (lizzieLet6_5_d[2:1])
        2'd0: is_z_kronai6_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_kronai6_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_kronai6_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_kronai6_goMux_mux_onehotd = 4'd8;
        default: is_z_kronai6_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_kronai6_goMux_mux_onehotd = 4'd0;
  assign _7_d = is_z_kronai6_goMux_mux_onehotd[0];
  assign lizzieLet6_5QVal_Int_d = is_z_kronai6_goMux_mux_onehotd[1];
  assign lizzieLet6_5QNode_Int_d = is_z_kronai6_goMux_mux_onehotd[2];
  assign _6_d = is_z_kronai6_goMux_mux_onehotd[3];
  assign is_z_kronai6_goMux_mux_r = (| (is_z_kronai6_goMux_mux_onehotd & {_6_r,
                                                                          lizzieLet6_5QNode_Int_r,
                                                                          lizzieLet6_5QVal_Int_r,
                                                                          _7_r}));
  assign lizzieLet6_5_r = is_z_kronai6_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int,MyDTInt_Bool) > [(lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                                                 (lizzieLet6_5QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_5QNode_Int_emitted;
  logic [1:0] lizzieLet6_5QNode_Int_done;
  assign lizzieLet6_5QNode_Int_1_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[0]));
  assign lizzieLet6_5QNode_Int_2_d = (lizzieLet6_5QNode_Int_d[0] && (! lizzieLet6_5QNode_Int_emitted[1]));
  assign lizzieLet6_5QNode_Int_done = (lizzieLet6_5QNode_Int_emitted | ({lizzieLet6_5QNode_Int_2_d[0],
                                                                         lizzieLet6_5QNode_Int_1_d[0]} & {lizzieLet6_5QNode_Int_2_r,
                                                                                                          lizzieLet6_5QNode_Int_1_r}));
  assign lizzieLet6_5QNode_Int_r = (& lizzieLet6_5QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_5QNode_Int_emitted <= (lizzieLet6_5QNode_Int_r ? 2'd0 :
                                        lizzieLet6_5QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_5QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_d;
  logic lizzieLet6_5QNode_Int_2_bufchan_r;
  assign lizzieLet6_5QNode_Int_2_r = ((! lizzieLet6_5QNode_Int_2_bufchan_d[0]) || lizzieLet6_5QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QNode_Int_2_r)
        lizzieLet6_5QNode_Int_2_bufchan_d <= lizzieLet6_5QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_5QNode_Int_2_bufchan_buf;
  assign lizzieLet6_5QNode_Int_2_bufchan_r = (! lizzieLet6_5QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_5QNode_Int_2_argbuf_d = (lizzieLet6_5QNode_Int_2_bufchan_buf[0] ? lizzieLet6_5QNode_Int_2_bufchan_buf :
                                             lizzieLet6_5QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QNode_Int_2_argbuf_r && lizzieLet6_5QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QNode_Int_2_argbuf_r) && (! lizzieLet6_5QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_5QNode_Int_2_bufchan_buf <= lizzieLet6_5QNode_Int_2_bufchan_d;
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_5QVal_Int,MyDTInt_Bool) > (lizzieLet6_5QVal_Int_1_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_d;
  logic lizzieLet6_5QVal_Int_bufchan_r;
  assign lizzieLet6_5QVal_Int_r = ((! lizzieLet6_5QVal_Int_bufchan_d[0]) || lizzieLet6_5QVal_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_5QVal_Int_r)
        lizzieLet6_5QVal_Int_bufchan_d <= lizzieLet6_5QVal_Int_d;
  MyDTInt_Bool_t lizzieLet6_5QVal_Int_bufchan_buf;
  assign lizzieLet6_5QVal_Int_bufchan_r = (! lizzieLet6_5QVal_Int_bufchan_buf[0]);
  assign lizzieLet6_5QVal_Int_1_argbuf_d = (lizzieLet6_5QVal_Int_bufchan_buf[0] ? lizzieLet6_5QVal_Int_bufchan_buf :
                                            lizzieLet6_5QVal_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_5QVal_Int_1_argbuf_r && lizzieLet6_5QVal_Int_bufchan_buf[0]))
        lizzieLet6_5QVal_Int_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_5QVal_Int_1_argbuf_r) && (! lizzieLet6_5QVal_Int_bufchan_buf[0])))
        lizzieLet6_5QVal_Int_bufchan_buf <= lizzieLet6_5QVal_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Bool) : (lizzieLet6_6,QTree_Int) (is_z_mapai9_goMux_mux,MyDTInt_Bool) > [(_5,MyDTInt_Bool),
                                                                                           (lizzieLet6_6QVal_Int,MyDTInt_Bool),
                                                                                           (lizzieLet6_6QNode_Int,MyDTInt_Bool),
                                                                                           (_4,MyDTInt_Bool)] */
  logic [3:0] is_z_mapai9_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_6_d[0] && is_z_mapai9_goMux_mux_d[0]))
      unique case (lizzieLet6_6_d[2:1])
        2'd0: is_z_mapai9_goMux_mux_onehotd = 4'd1;
        2'd1: is_z_mapai9_goMux_mux_onehotd = 4'd2;
        2'd2: is_z_mapai9_goMux_mux_onehotd = 4'd4;
        2'd3: is_z_mapai9_goMux_mux_onehotd = 4'd8;
        default: is_z_mapai9_goMux_mux_onehotd = 4'd0;
      endcase
    else is_z_mapai9_goMux_mux_onehotd = 4'd0;
  assign _5_d = is_z_mapai9_goMux_mux_onehotd[0];
  assign lizzieLet6_6QVal_Int_d = is_z_mapai9_goMux_mux_onehotd[1];
  assign lizzieLet6_6QNode_Int_d = is_z_mapai9_goMux_mux_onehotd[2];
  assign _4_d = is_z_mapai9_goMux_mux_onehotd[3];
  assign is_z_mapai9_goMux_mux_r = (| (is_z_mapai9_goMux_mux_onehotd & {_4_r,
                                                                        lizzieLet6_6QNode_Int_r,
                                                                        lizzieLet6_6QVal_Int_r,
                                                                        _5_r}));
  assign lizzieLet6_6_r = is_z_mapai9_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Bool) : (lizzieLet6_6QNode_Int,MyDTInt_Bool) > [(lizzieLet6_6QNode_Int_1,MyDTInt_Bool),
                                                                 (lizzieLet6_6QNode_Int_2,MyDTInt_Bool)] */
  logic [1:0] lizzieLet6_6QNode_Int_emitted;
  logic [1:0] lizzieLet6_6QNode_Int_done;
  assign lizzieLet6_6QNode_Int_1_d = (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[0]));
  assign lizzieLet6_6QNode_Int_2_d = (lizzieLet6_6QNode_Int_d[0] && (! lizzieLet6_6QNode_Int_emitted[1]));
  assign lizzieLet6_6QNode_Int_done = (lizzieLet6_6QNode_Int_emitted | ({lizzieLet6_6QNode_Int_2_d[0],
                                                                         lizzieLet6_6QNode_Int_1_d[0]} & {lizzieLet6_6QNode_Int_2_r,
                                                                                                          lizzieLet6_6QNode_Int_1_r}));
  assign lizzieLet6_6QNode_Int_r = (& lizzieLet6_6QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_6QNode_Int_emitted <= (lizzieLet6_6QNode_Int_r ? 2'd0 :
                                        lizzieLet6_6QNode_Int_done);
  
  /* buf (Ty MyDTInt_Bool) : (lizzieLet6_6QNode_Int_2,MyDTInt_Bool) > (lizzieLet6_6QNode_Int_2_argbuf,MyDTInt_Bool) */
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_2_bufchan_d;
  logic lizzieLet6_6QNode_Int_2_bufchan_r;
  assign lizzieLet6_6QNode_Int_2_r = ((! lizzieLet6_6QNode_Int_2_bufchan_d[0]) || lizzieLet6_6QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_6QNode_Int_2_r)
        lizzieLet6_6QNode_Int_2_bufchan_d <= lizzieLet6_6QNode_Int_2_d;
  MyDTInt_Bool_t lizzieLet6_6QNode_Int_2_bufchan_buf;
  assign lizzieLet6_6QNode_Int_2_bufchan_r = (! lizzieLet6_6QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_6QNode_Int_2_argbuf_d = (lizzieLet6_6QNode_Int_2_bufchan_buf[0] ? lizzieLet6_6QNode_Int_2_bufchan_buf :
                                             lizzieLet6_6QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_6QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_6QNode_Int_2_argbuf_r && lizzieLet6_6QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_6QNode_Int_2_argbuf_r) && (! lizzieLet6_6QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_6QNode_Int_2_bufchan_buf <= lizzieLet6_6QNode_Int_2_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty MyDTInt_Int_Int) : (lizzieLet6_7,QTree_Int) (op_kronai7_goMux_mux,MyDTInt_Int_Int) > [(_3,MyDTInt_Int_Int),
                                                                                                (lizzieLet6_7QVal_Int,MyDTInt_Int_Int),
                                                                                                (lizzieLet6_7QNode_Int,MyDTInt_Int_Int),
                                                                                                (_2,MyDTInt_Int_Int)] */
  logic [3:0] op_kronai7_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_7_d[0] && op_kronai7_goMux_mux_d[0]))
      unique case (lizzieLet6_7_d[2:1])
        2'd0: op_kronai7_goMux_mux_onehotd = 4'd1;
        2'd1: op_kronai7_goMux_mux_onehotd = 4'd2;
        2'd2: op_kronai7_goMux_mux_onehotd = 4'd4;
        2'd3: op_kronai7_goMux_mux_onehotd = 4'd8;
        default: op_kronai7_goMux_mux_onehotd = 4'd0;
      endcase
    else op_kronai7_goMux_mux_onehotd = 4'd0;
  assign _3_d = op_kronai7_goMux_mux_onehotd[0];
  assign lizzieLet6_7QVal_Int_d = op_kronai7_goMux_mux_onehotd[1];
  assign lizzieLet6_7QNode_Int_d = op_kronai7_goMux_mux_onehotd[2];
  assign _2_d = op_kronai7_goMux_mux_onehotd[3];
  assign op_kronai7_goMux_mux_r = (| (op_kronai7_goMux_mux_onehotd & {_2_r,
                                                                      lizzieLet6_7QNode_Int_r,
                                                                      lizzieLet6_7QVal_Int_r,
                                                                      _3_r}));
  assign lizzieLet6_7_r = op_kronai7_goMux_mux_r;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_7QNode_Int,MyDTInt_Int_Int) > [(lizzieLet6_7QNode_Int_1,MyDTInt_Int_Int),
                                                                       (lizzieLet6_7QNode_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_7QNode_Int_emitted;
  logic [1:0] lizzieLet6_7QNode_Int_done;
  assign lizzieLet6_7QNode_Int_1_d = (lizzieLet6_7QNode_Int_d[0] && (! lizzieLet6_7QNode_Int_emitted[0]));
  assign lizzieLet6_7QNode_Int_2_d = (lizzieLet6_7QNode_Int_d[0] && (! lizzieLet6_7QNode_Int_emitted[1]));
  assign lizzieLet6_7QNode_Int_done = (lizzieLet6_7QNode_Int_emitted | ({lizzieLet6_7QNode_Int_2_d[0],
                                                                         lizzieLet6_7QNode_Int_1_d[0]} & {lizzieLet6_7QNode_Int_2_r,
                                                                                                          lizzieLet6_7QNode_Int_1_r}));
  assign lizzieLet6_7QNode_Int_r = (& lizzieLet6_7QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_7QNode_Int_emitted <= (lizzieLet6_7QNode_Int_r ? 2'd0 :
                                        lizzieLet6_7QNode_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_7QNode_Int_2,MyDTInt_Int_Int) > (lizzieLet6_7QNode_Int_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_2_bufchan_d;
  logic lizzieLet6_7QNode_Int_2_bufchan_r;
  assign lizzieLet6_7QNode_Int_2_r = ((! lizzieLet6_7QNode_Int_2_bufchan_d[0]) || lizzieLet6_7QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QNode_Int_2_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_7QNode_Int_2_r)
        lizzieLet6_7QNode_Int_2_bufchan_d <= lizzieLet6_7QNode_Int_2_d;
  MyDTInt_Int_Int_t lizzieLet6_7QNode_Int_2_bufchan_buf;
  assign lizzieLet6_7QNode_Int_2_bufchan_r = (! lizzieLet6_7QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_7QNode_Int_2_argbuf_d = (lizzieLet6_7QNode_Int_2_bufchan_buf[0] ? lizzieLet6_7QNode_Int_2_bufchan_buf :
                                             lizzieLet6_7QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QNode_Int_2_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_7QNode_Int_2_argbuf_r && lizzieLet6_7QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_7QNode_Int_2_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_7QNode_Int_2_argbuf_r) && (! lizzieLet6_7QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_7QNode_Int_2_bufchan_buf <= lizzieLet6_7QNode_Int_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (lizzieLet6_7QVal_Int,MyDTInt_Int_Int) > [(lizzieLet6_7QVal_Int_1,MyDTInt_Int_Int),
                                                                      (lizzieLet6_7QVal_Int_2,MyDTInt_Int_Int)] */
  logic [1:0] lizzieLet6_7QVal_Int_emitted;
  logic [1:0] lizzieLet6_7QVal_Int_done;
  assign lizzieLet6_7QVal_Int_1_d = (lizzieLet6_7QVal_Int_d[0] && (! lizzieLet6_7QVal_Int_emitted[0]));
  assign lizzieLet6_7QVal_Int_2_d = (lizzieLet6_7QVal_Int_d[0] && (! lizzieLet6_7QVal_Int_emitted[1]));
  assign lizzieLet6_7QVal_Int_done = (lizzieLet6_7QVal_Int_emitted | ({lizzieLet6_7QVal_Int_2_d[0],
                                                                       lizzieLet6_7QVal_Int_1_d[0]} & {lizzieLet6_7QVal_Int_2_r,
                                                                                                       lizzieLet6_7QVal_Int_1_r}));
  assign lizzieLet6_7QVal_Int_r = (& lizzieLet6_7QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_7QVal_Int_emitted <= (lizzieLet6_7QVal_Int_r ? 2'd0 :
                                       lizzieLet6_7QVal_Int_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (lizzieLet6_7QVal_Int_1,MyDTInt_Int_Int) > (lizzieLet6_7QVal_Int_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_1_bufchan_d;
  logic lizzieLet6_7QVal_Int_1_bufchan_r;
  assign lizzieLet6_7QVal_Int_1_r = ((! lizzieLet6_7QVal_Int_1_bufchan_d[0]) || lizzieLet6_7QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QVal_Int_1_bufchan_d <= 1'd0;
    else
      if (lizzieLet6_7QVal_Int_1_r)
        lizzieLet6_7QVal_Int_1_bufchan_d <= lizzieLet6_7QVal_Int_1_d;
  MyDTInt_Int_Int_t lizzieLet6_7QVal_Int_1_bufchan_buf;
  assign lizzieLet6_7QVal_Int_1_bufchan_r = (! lizzieLet6_7QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_7QVal_Int_1_argbuf_d = (lizzieLet6_7QVal_Int_1_bufchan_buf[0] ? lizzieLet6_7QVal_Int_1_bufchan_buf :
                                            lizzieLet6_7QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_7QVal_Int_1_bufchan_buf <= 1'd0;
    else
      if ((lizzieLet6_7QVal_Int_1_argbuf_r && lizzieLet6_7QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_7QVal_Int_1_bufchan_buf <= 1'd0;
      else if (((! lizzieLet6_7QVal_Int_1_argbuf_r) && (! lizzieLet6_7QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_7QVal_Int_1_bufchan_buf <= lizzieLet6_7QVal_Int_1_bufchan_d;
  
  /* dcon (Ty TupMyDTInt_Int_Int___Int___Int,
      Dcon TupMyDTInt_Int_Int___Int___Int) : [(lizzieLet6_7QVal_Int_1_argbuf,MyDTInt_Int_Int),
                                              (lizzieLet6_9QVal_Int_1_argbuf,Int),
                                              (v'aib_1_argbuf,Int)] > (applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1,TupMyDTInt_Int_Int___Int___Int) */
  assign applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d = TupMyDTInt_Int_Int___Int___Int_dc((& {lizzieLet6_7QVal_Int_1_argbuf_d[0],
                                                                                                        lizzieLet6_9QVal_Int_1_argbuf_d[0],
                                                                                                        \v'aib_1_argbuf_d [0]}), lizzieLet6_7QVal_Int_1_argbuf_d, lizzieLet6_9QVal_Int_1_argbuf_d, \v'aib_1_argbuf_d );
  assign {lizzieLet6_7QVal_Int_1_argbuf_r,
          lizzieLet6_9QVal_Int_1_argbuf_r,
          \v'aib_1_argbuf_r } = {3 {(applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_r && applyfnInt_Int_Int_5TupMyDTInt_Int_Int___Int___Int_1_d[0])}};
  
  /* demux (Ty QTree_Int,
       Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (lizzieLet6_8,QTree_Int) (sc_0_1_goMux_mux,Pointer_CTf'_f'_Int_Int_Int_Int) > [(lizzieLet6_8QNone_Int,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet6_8QVal_Int,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet6_8QNode_Int,Pointer_CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet6_8QError_Int,Pointer_CTf'_f'_Int_Int_Int_Int)] */
  logic [3:0] sc_0_1_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_8_d[0] && sc_0_1_goMux_mux_d[0]))
      unique case (lizzieLet6_8_d[2:1])
        2'd0: sc_0_1_goMux_mux_onehotd = 4'd1;
        2'd1: sc_0_1_goMux_mux_onehotd = 4'd2;
        2'd2: sc_0_1_goMux_mux_onehotd = 4'd4;
        2'd3: sc_0_1_goMux_mux_onehotd = 4'd8;
        default: sc_0_1_goMux_mux_onehotd = 4'd0;
      endcase
    else sc_0_1_goMux_mux_onehotd = 4'd0;
  assign lizzieLet6_8QNone_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[0]};
  assign lizzieLet6_8QVal_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                   sc_0_1_goMux_mux_onehotd[1]};
  assign lizzieLet6_8QNode_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                    sc_0_1_goMux_mux_onehotd[2]};
  assign lizzieLet6_8QError_Int_d = {sc_0_1_goMux_mux_d[16:1],
                                     sc_0_1_goMux_mux_onehotd[3]};
  assign sc_0_1_goMux_mux_r = (| (sc_0_1_goMux_mux_onehotd & {lizzieLet6_8QError_Int_r,
                                                              lizzieLet6_8QNode_Int_r,
                                                              lizzieLet6_8QVal_Int_r,
                                                              lizzieLet6_8QNone_Int_r}));
  assign lizzieLet6_8_r = sc_0_1_goMux_mux_r;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (lizzieLet6_8QError_Int,Pointer_CTf'_f'_Int_Int_Int_Int) > (lizzieLet6_8QError_Int_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QError_Int_bufchan_d;
  logic lizzieLet6_8QError_Int_bufchan_r;
  assign lizzieLet6_8QError_Int_r = ((! lizzieLet6_8QError_Int_bufchan_d[0]) || lizzieLet6_8QError_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QError_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_8QError_Int_r)
        lizzieLet6_8QError_Int_bufchan_d <= lizzieLet6_8QError_Int_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QError_Int_bufchan_buf;
  assign lizzieLet6_8QError_Int_bufchan_r = (! lizzieLet6_8QError_Int_bufchan_buf[0]);
  assign lizzieLet6_8QError_Int_1_argbuf_d = (lizzieLet6_8QError_Int_bufchan_buf[0] ? lizzieLet6_8QError_Int_bufchan_buf :
                                              lizzieLet6_8QError_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_8QError_Int_1_argbuf_r && lizzieLet6_8QError_Int_bufchan_buf[0]))
        lizzieLet6_8QError_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_8QError_Int_1_argbuf_r) && (! lizzieLet6_8QError_Int_bufchan_buf[0])))
        lizzieLet6_8QError_Int_bufchan_buf <= lizzieLet6_8QError_Int_bufchan_d;
  
  /* dcon (Ty CTf'_f'_Int_Int_Int_Int,
      Dcon Lcall_f'_f'_Int_Int_Int_Int3) : [(lizzieLet6_8QNode_Int,Pointer_CTf'_f'_Int_Int_Int_Int),
                                            (q1aic_destruct,Pointer_QTree_Int),
                                            (lizzieLet6_5QNode_Int_1,MyDTInt_Bool),
                                            (lizzieLet6_7QNode_Int_1,MyDTInt_Int_Int),
                                            (lizzieLet6_9QNode_Int_1,Int),
                                            (lizzieLet6_6QNode_Int_1,MyDTInt_Bool),
                                            (lizzieLet6_3QNode_Int_1,MyDTInt_Int),
                                            (q2aid_destruct,Pointer_QTree_Int),
                                            (q3aie_destruct,Pointer_QTree_Int)] > (lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3,CTf'_f'_Int_Int_Int_Int) */
  assign \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_d  = \Lcall_f'_f'_Int_Int_Int_Int3_dc ((& {lizzieLet6_8QNode_Int_d[0],
                                                                                                                                                                                                                                                 q1aic_destruct_d[0],
                                                                                                                                                                                                                                                 lizzieLet6_5QNode_Int_1_d[0],
                                                                                                                                                                                                                                                 lizzieLet6_7QNode_Int_1_d[0],
                                                                                                                                                                                                                                                 lizzieLet6_9QNode_Int_1_d[0],
                                                                                                                                                                                                                                                 lizzieLet6_6QNode_Int_1_d[0],
                                                                                                                                                                                                                                                 lizzieLet6_3QNode_Int_1_d[0],
                                                                                                                                                                                                                                                 q2aid_destruct_d[0],
                                                                                                                                                                                                                                                 q3aie_destruct_d[0]}), lizzieLet6_8QNode_Int_d, q1aic_destruct_d, lizzieLet6_5QNode_Int_1_d, lizzieLet6_7QNode_Int_1_d, lizzieLet6_9QNode_Int_1_d, lizzieLet6_6QNode_Int_1_d, lizzieLet6_3QNode_Int_1_d, q2aid_destruct_d, q3aie_destruct_d);
  assign {lizzieLet6_8QNode_Int_r,
          q1aic_destruct_r,
          lizzieLet6_5QNode_Int_1_r,
          lizzieLet6_7QNode_Int_1_r,
          lizzieLet6_9QNode_Int_1_r,
          lizzieLet6_6QNode_Int_1_r,
          lizzieLet6_3QNode_Int_1_r,
          q2aid_destruct_r,
          q3aie_destruct_r} = {9 {(\lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_r  && \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_d [0])}};
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3,CTf'_f'_Int_Int_Int_Int) > (lizzieLet11_2_1_argbuf,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d ;
  logic \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r ;
  assign \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_r  = ((! \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d [0]) || \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d  <= {99'd0,
                                                                                                                                                                                                                  1'd0};
    else
      if (\lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_r )
        \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d  <= \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf ;
  assign \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_r  = (! \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0]);
  assign lizzieLet11_2_1_argbuf_d = (\lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0] ? \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  :
                                     \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                                                                    1'd0};
    else
      if ((lizzieLet11_2_1_argbuf_r && \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0]))
        \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= {99'd0,
                                                                                                                                                                                                                      1'd0};
      else if (((! lizzieLet11_2_1_argbuf_r) && (! \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf [0])))
        \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_buf  <= \lizzieLet6_8QNode_Int_1q1aic_1lizzieLet6_5QNode_Int_1lizzieLet6_7QNode_Int_1lizzieLet6_9QNode_Int_1lizzieLet6_6QNode_Int_1lizzieLet6_3QNode_Int_1q2aid_1q3aie_1Lcall_f'_f'_Int_Int_Int_Int3_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (lizzieLet6_8QNone_Int,Pointer_CTf'_f'_Int_Int_Int_Int) > (lizzieLet6_8QNone_Int_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QNone_Int_bufchan_d;
  logic lizzieLet6_8QNone_Int_bufchan_r;
  assign lizzieLet6_8QNone_Int_r = ((! lizzieLet6_8QNone_Int_bufchan_d[0]) || lizzieLet6_8QNone_Int_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QNone_Int_bufchan_d <= {16'd0, 1'd0};
    else
      if (lizzieLet6_8QNone_Int_r)
        lizzieLet6_8QNone_Int_bufchan_d <= lizzieLet6_8QNone_Int_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  lizzieLet6_8QNone_Int_bufchan_buf;
  assign lizzieLet6_8QNone_Int_bufchan_r = (! lizzieLet6_8QNone_Int_bufchan_buf[0]);
  assign lizzieLet6_8QNone_Int_1_argbuf_d = (lizzieLet6_8QNone_Int_bufchan_buf[0] ? lizzieLet6_8QNone_Int_bufchan_buf :
                                             lizzieLet6_8QNone_Int_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet6_8QNone_Int_1_argbuf_r && lizzieLet6_8QNone_Int_bufchan_buf[0]))
        lizzieLet6_8QNone_Int_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet6_8QNone_Int_1_argbuf_r) && (! lizzieLet6_8QNone_Int_bufchan_buf[0])))
        lizzieLet6_8QNone_Int_bufchan_buf <= lizzieLet6_8QNone_Int_bufchan_d;
  
  /* demux (Ty QTree_Int,
       Ty Int) : (lizzieLet6_9,QTree_Int) (vai8_goMux_mux,Int) > [(_1,Int),
                                                                  (lizzieLet6_9QVal_Int,Int),
                                                                  (lizzieLet6_9QNode_Int,Int),
                                                                  (_0,Int)] */
  logic [3:0] vai8_goMux_mux_onehotd;
  always_comb
    if ((lizzieLet6_9_d[0] && vai8_goMux_mux_d[0]))
      unique case (lizzieLet6_9_d[2:1])
        2'd0: vai8_goMux_mux_onehotd = 4'd1;
        2'd1: vai8_goMux_mux_onehotd = 4'd2;
        2'd2: vai8_goMux_mux_onehotd = 4'd4;
        2'd3: vai8_goMux_mux_onehotd = 4'd8;
        default: vai8_goMux_mux_onehotd = 4'd0;
      endcase
    else vai8_goMux_mux_onehotd = 4'd0;
  assign _1_d = {vai8_goMux_mux_d[32:1], vai8_goMux_mux_onehotd[0]};
  assign lizzieLet6_9QVal_Int_d = {vai8_goMux_mux_d[32:1],
                                   vai8_goMux_mux_onehotd[1]};
  assign lizzieLet6_9QNode_Int_d = {vai8_goMux_mux_d[32:1],
                                    vai8_goMux_mux_onehotd[2]};
  assign _0_d = {vai8_goMux_mux_d[32:1], vai8_goMux_mux_onehotd[3]};
  assign vai8_goMux_mux_r = (| (vai8_goMux_mux_onehotd & {_0_r,
                                                          lizzieLet6_9QNode_Int_r,
                                                          lizzieLet6_9QVal_Int_r,
                                                          _1_r}));
  assign lizzieLet6_9_r = vai8_goMux_mux_r;
  
  /* fork (Ty Int) : (lizzieLet6_9QNode_Int,Int) > [(lizzieLet6_9QNode_Int_1,Int),
                                               (lizzieLet6_9QNode_Int_2,Int)] */
  logic [1:0] lizzieLet6_9QNode_Int_emitted;
  logic [1:0] lizzieLet6_9QNode_Int_done;
  assign lizzieLet6_9QNode_Int_1_d = {lizzieLet6_9QNode_Int_d[32:1],
                                      (lizzieLet6_9QNode_Int_d[0] && (! lizzieLet6_9QNode_Int_emitted[0]))};
  assign lizzieLet6_9QNode_Int_2_d = {lizzieLet6_9QNode_Int_d[32:1],
                                      (lizzieLet6_9QNode_Int_d[0] && (! lizzieLet6_9QNode_Int_emitted[1]))};
  assign lizzieLet6_9QNode_Int_done = (lizzieLet6_9QNode_Int_emitted | ({lizzieLet6_9QNode_Int_2_d[0],
                                                                         lizzieLet6_9QNode_Int_1_d[0]} & {lizzieLet6_9QNode_Int_2_r,
                                                                                                          lizzieLet6_9QNode_Int_1_r}));
  assign lizzieLet6_9QNode_Int_r = (& lizzieLet6_9QNode_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_9QNode_Int_emitted <= 2'd0;
    else
      lizzieLet6_9QNode_Int_emitted <= (lizzieLet6_9QNode_Int_r ? 2'd0 :
                                        lizzieLet6_9QNode_Int_done);
  
  /* buf (Ty Int) : (lizzieLet6_9QNode_Int_2,Int) > (lizzieLet6_9QNode_Int_2_argbuf,Int) */
  Int_t lizzieLet6_9QNode_Int_2_bufchan_d;
  logic lizzieLet6_9QNode_Int_2_bufchan_r;
  assign lizzieLet6_9QNode_Int_2_r = ((! lizzieLet6_9QNode_Int_2_bufchan_d[0]) || lizzieLet6_9QNode_Int_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QNode_Int_2_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet6_9QNode_Int_2_r)
        lizzieLet6_9QNode_Int_2_bufchan_d <= lizzieLet6_9QNode_Int_2_d;
  Int_t lizzieLet6_9QNode_Int_2_bufchan_buf;
  assign lizzieLet6_9QNode_Int_2_bufchan_r = (! lizzieLet6_9QNode_Int_2_bufchan_buf[0]);
  assign lizzieLet6_9QNode_Int_2_argbuf_d = (lizzieLet6_9QNode_Int_2_bufchan_buf[0] ? lizzieLet6_9QNode_Int_2_bufchan_buf :
                                             lizzieLet6_9QNode_Int_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet6_9QNode_Int_2_argbuf_r && lizzieLet6_9QNode_Int_2_bufchan_buf[0]))
        lizzieLet6_9QNode_Int_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet6_9QNode_Int_2_argbuf_r) && (! lizzieLet6_9QNode_Int_2_bufchan_buf[0])))
        lizzieLet6_9QNode_Int_2_bufchan_buf <= lizzieLet6_9QNode_Int_2_bufchan_d;
  
  /* fork (Ty Int) : (lizzieLet6_9QVal_Int,Int) > [(lizzieLet6_9QVal_Int_1,Int),
                                              (lizzieLet6_9QVal_Int_2,Int)] */
  logic [1:0] lizzieLet6_9QVal_Int_emitted;
  logic [1:0] lizzieLet6_9QVal_Int_done;
  assign lizzieLet6_9QVal_Int_1_d = {lizzieLet6_9QVal_Int_d[32:1],
                                     (lizzieLet6_9QVal_Int_d[0] && (! lizzieLet6_9QVal_Int_emitted[0]))};
  assign lizzieLet6_9QVal_Int_2_d = {lizzieLet6_9QVal_Int_d[32:1],
                                     (lizzieLet6_9QVal_Int_d[0] && (! lizzieLet6_9QVal_Int_emitted[1]))};
  assign lizzieLet6_9QVal_Int_done = (lizzieLet6_9QVal_Int_emitted | ({lizzieLet6_9QVal_Int_2_d[0],
                                                                       lizzieLet6_9QVal_Int_1_d[0]} & {lizzieLet6_9QVal_Int_2_r,
                                                                                                       lizzieLet6_9QVal_Int_1_r}));
  assign lizzieLet6_9QVal_Int_r = (& lizzieLet6_9QVal_Int_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) lizzieLet6_9QVal_Int_emitted <= 2'd0;
    else
      lizzieLet6_9QVal_Int_emitted <= (lizzieLet6_9QVal_Int_r ? 2'd0 :
                                       lizzieLet6_9QVal_Int_done);
  
  /* buf (Ty Int) : (lizzieLet6_9QVal_Int_1,Int) > (lizzieLet6_9QVal_Int_1_argbuf,Int) */
  Int_t lizzieLet6_9QVal_Int_1_bufchan_d;
  logic lizzieLet6_9QVal_Int_1_bufchan_r;
  assign lizzieLet6_9QVal_Int_1_r = ((! lizzieLet6_9QVal_Int_1_bufchan_d[0]) || lizzieLet6_9QVal_Int_1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QVal_Int_1_bufchan_d <= {32'd0, 1'd0};
    else
      if (lizzieLet6_9QVal_Int_1_r)
        lizzieLet6_9QVal_Int_1_bufchan_d <= lizzieLet6_9QVal_Int_1_d;
  Int_t lizzieLet6_9QVal_Int_1_bufchan_buf;
  assign lizzieLet6_9QVal_Int_1_bufchan_r = (! lizzieLet6_9QVal_Int_1_bufchan_buf[0]);
  assign lizzieLet6_9QVal_Int_1_argbuf_d = (lizzieLet6_9QVal_Int_1_bufchan_buf[0] ? lizzieLet6_9QVal_Int_1_bufchan_buf :
                                            lizzieLet6_9QVal_Int_1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      lizzieLet6_9QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((lizzieLet6_9QVal_Int_1_argbuf_r && lizzieLet6_9QVal_Int_1_bufchan_buf[0]))
        lizzieLet6_9QVal_Int_1_bufchan_buf <= {32'd0, 1'd0};
      else if (((! lizzieLet6_9QVal_Int_1_argbuf_r) && (! lizzieLet6_9QVal_Int_1_bufchan_buf[0])))
        lizzieLet6_9QVal_Int_1_bufchan_buf <= lizzieLet6_9QVal_Int_1_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m1ahU_goMux_mux,Pointer_QTree_Int) > (m1ahU_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m1ahU_goMux_mux_bufchan_d;
  logic m1ahU_goMux_mux_bufchan_r;
  assign m1ahU_goMux_mux_r = ((! m1ahU_goMux_mux_bufchan_d[0]) || m1ahU_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ahU_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m1ahU_goMux_mux_r)
        m1ahU_goMux_mux_bufchan_d <= m1ahU_goMux_mux_d;
  Pointer_QTree_Int_t m1ahU_goMux_mux_bufchan_buf;
  assign m1ahU_goMux_mux_bufchan_r = (! m1ahU_goMux_mux_bufchan_buf[0]);
  assign m1ahU_1_argbuf_d = (m1ahU_goMux_mux_bufchan_buf[0] ? m1ahU_goMux_mux_bufchan_buf :
                             m1ahU_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m1ahU_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m1ahU_1_argbuf_r && m1ahU_goMux_mux_bufchan_buf[0]))
        m1ahU_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m1ahU_1_argbuf_r) && (! m1ahU_goMux_mux_bufchan_buf[0])))
        m1ahU_goMux_mux_bufchan_buf <= m1ahU_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2ahV_2_2,Pointer_QTree_Int) > (m2ahV_2_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ahV_2_2_bufchan_d;
  logic m2ahV_2_2_bufchan_r;
  assign m2ahV_2_2_r = ((! m2ahV_2_2_bufchan_d[0]) || m2ahV_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_2_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ahV_2_2_r) m2ahV_2_2_bufchan_d <= m2ahV_2_2_d;
  Pointer_QTree_Int_t m2ahV_2_2_bufchan_buf;
  assign m2ahV_2_2_bufchan_r = (! m2ahV_2_2_bufchan_buf[0]);
  assign m2ahV_2_2_argbuf_d = (m2ahV_2_2_bufchan_buf[0] ? m2ahV_2_2_bufchan_buf :
                               m2ahV_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_2_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ahV_2_2_argbuf_r && m2ahV_2_2_bufchan_buf[0]))
        m2ahV_2_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ahV_2_2_argbuf_r) && (! m2ahV_2_2_bufchan_buf[0])))
        m2ahV_2_2_bufchan_buf <= m2ahV_2_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2ahV_2_destruct,Pointer_QTree_Int) > [(m2ahV_2_1,Pointer_QTree_Int),
                                                                      (m2ahV_2_2,Pointer_QTree_Int)] */
  logic [1:0] m2ahV_2_destruct_emitted;
  logic [1:0] m2ahV_2_destruct_done;
  assign m2ahV_2_1_d = {m2ahV_2_destruct_d[16:1],
                        (m2ahV_2_destruct_d[0] && (! m2ahV_2_destruct_emitted[0]))};
  assign m2ahV_2_2_d = {m2ahV_2_destruct_d[16:1],
                        (m2ahV_2_destruct_d[0] && (! m2ahV_2_destruct_emitted[1]))};
  assign m2ahV_2_destruct_done = (m2ahV_2_destruct_emitted | ({m2ahV_2_2_d[0],
                                                               m2ahV_2_1_d[0]} & {m2ahV_2_2_r,
                                                                                  m2ahV_2_1_r}));
  assign m2ahV_2_destruct_r = (& m2ahV_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_2_destruct_emitted <= 2'd0;
    else
      m2ahV_2_destruct_emitted <= (m2ahV_2_destruct_r ? 2'd0 :
                                   m2ahV_2_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2ahV_3_2,Pointer_QTree_Int) > (m2ahV_3_2_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ahV_3_2_bufchan_d;
  logic m2ahV_3_2_bufchan_r;
  assign m2ahV_3_2_r = ((! m2ahV_3_2_bufchan_d[0]) || m2ahV_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_3_2_bufchan_d <= {16'd0, 1'd0};
    else if (m2ahV_3_2_r) m2ahV_3_2_bufchan_d <= m2ahV_3_2_d;
  Pointer_QTree_Int_t m2ahV_3_2_bufchan_buf;
  assign m2ahV_3_2_bufchan_r = (! m2ahV_3_2_bufchan_buf[0]);
  assign m2ahV_3_2_argbuf_d = (m2ahV_3_2_bufchan_buf[0] ? m2ahV_3_2_bufchan_buf :
                               m2ahV_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_3_2_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ahV_3_2_argbuf_r && m2ahV_3_2_bufchan_buf[0]))
        m2ahV_3_2_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ahV_3_2_argbuf_r) && (! m2ahV_3_2_bufchan_buf[0])))
        m2ahV_3_2_bufchan_buf <= m2ahV_3_2_bufchan_d;
  
  /* fork (Ty Pointer_QTree_Int) : (m2ahV_3_destruct,Pointer_QTree_Int) > [(m2ahV_3_1,Pointer_QTree_Int),
                                                                      (m2ahV_3_2,Pointer_QTree_Int)] */
  logic [1:0] m2ahV_3_destruct_emitted;
  logic [1:0] m2ahV_3_destruct_done;
  assign m2ahV_3_1_d = {m2ahV_3_destruct_d[16:1],
                        (m2ahV_3_destruct_d[0] && (! m2ahV_3_destruct_emitted[0]))};
  assign m2ahV_3_2_d = {m2ahV_3_destruct_d[16:1],
                        (m2ahV_3_destruct_d[0] && (! m2ahV_3_destruct_emitted[1]))};
  assign m2ahV_3_destruct_done = (m2ahV_3_destruct_emitted | ({m2ahV_3_2_d[0],
                                                               m2ahV_3_1_d[0]} & {m2ahV_3_2_r,
                                                                                  m2ahV_3_1_r}));
  assign m2ahV_3_destruct_r = (& m2ahV_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_3_destruct_emitted <= 2'd0;
    else
      m2ahV_3_destruct_emitted <= (m2ahV_3_destruct_r ? 2'd0 :
                                   m2ahV_3_destruct_done);
  
  /* buf (Ty Pointer_QTree_Int) : (m2ahV_4_destruct,Pointer_QTree_Int) > (m2ahV_4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ahV_4_destruct_bufchan_d;
  logic m2ahV_4_destruct_bufchan_r;
  assign m2ahV_4_destruct_r = ((! m2ahV_4_destruct_bufchan_d[0]) || m2ahV_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2ahV_4_destruct_r)
        m2ahV_4_destruct_bufchan_d <= m2ahV_4_destruct_d;
  Pointer_QTree_Int_t m2ahV_4_destruct_bufchan_buf;
  assign m2ahV_4_destruct_bufchan_r = (! m2ahV_4_destruct_bufchan_buf[0]);
  assign m2ahV_4_1_argbuf_d = (m2ahV_4_destruct_bufchan_buf[0] ? m2ahV_4_destruct_bufchan_buf :
                               m2ahV_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ahV_4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ahV_4_1_argbuf_r && m2ahV_4_destruct_bufchan_buf[0]))
        m2ahV_4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ahV_4_1_argbuf_r) && (! m2ahV_4_destruct_bufchan_buf[0])))
        m2ahV_4_destruct_bufchan_buf <= m2ahV_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (m2ai5_goMux_mux,Pointer_QTree_Int) > (m2ai5_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t m2ai5_goMux_mux_bufchan_d;
  logic m2ai5_goMux_mux_bufchan_r;
  assign m2ai5_goMux_mux_r = ((! m2ai5_goMux_mux_bufchan_d[0]) || m2ai5_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ai5_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (m2ai5_goMux_mux_r)
        m2ai5_goMux_mux_bufchan_d <= m2ai5_goMux_mux_d;
  Pointer_QTree_Int_t m2ai5_goMux_mux_bufchan_buf;
  assign m2ai5_goMux_mux_bufchan_r = (! m2ai5_goMux_mux_bufchan_buf[0]);
  assign m2ai5_1_argbuf_d = (m2ai5_goMux_mux_bufchan_buf[0] ? m2ai5_goMux_mux_bufchan_buf :
                             m2ai5_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) m2ai5_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((m2ai5_1_argbuf_r && m2ai5_goMux_mux_bufchan_buf[0]))
        m2ai5_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! m2ai5_1_argbuf_r) && (! m2ai5_goMux_mux_bufchan_buf[0])))
        m2ai5_goMux_mux_bufchan_buf <= m2ai5_goMux_mux_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronahX_2_2,MyDTInt_Int_Int) > (op_kronahX_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronahX_2_2_bufchan_d;
  logic op_kronahX_2_2_bufchan_r;
  assign op_kronahX_2_2_r = ((! op_kronahX_2_2_bufchan_d[0]) || op_kronahX_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_2_2_bufchan_d <= 1'd0;
    else
      if (op_kronahX_2_2_r) op_kronahX_2_2_bufchan_d <= op_kronahX_2_2_d;
  MyDTInt_Int_Int_t op_kronahX_2_2_bufchan_buf;
  assign op_kronahX_2_2_bufchan_r = (! op_kronahX_2_2_bufchan_buf[0]);
  assign op_kronahX_2_2_argbuf_d = (op_kronahX_2_2_bufchan_buf[0] ? op_kronahX_2_2_bufchan_buf :
                                    op_kronahX_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_kronahX_2_2_argbuf_r && op_kronahX_2_2_bufchan_buf[0]))
        op_kronahX_2_2_bufchan_buf <= 1'd0;
      else if (((! op_kronahX_2_2_argbuf_r) && (! op_kronahX_2_2_bufchan_buf[0])))
        op_kronahX_2_2_bufchan_buf <= op_kronahX_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_kronahX_2_destruct,MyDTInt_Int_Int) > [(op_kronahX_2_1,MyDTInt_Int_Int),
                                                                       (op_kronahX_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_kronahX_2_destruct_emitted;
  logic [1:0] op_kronahX_2_destruct_done;
  assign op_kronahX_2_1_d = (op_kronahX_2_destruct_d[0] && (! op_kronahX_2_destruct_emitted[0]));
  assign op_kronahX_2_2_d = (op_kronahX_2_destruct_d[0] && (! op_kronahX_2_destruct_emitted[1]));
  assign op_kronahX_2_destruct_done = (op_kronahX_2_destruct_emitted | ({op_kronahX_2_2_d[0],
                                                                         op_kronahX_2_1_d[0]} & {op_kronahX_2_2_r,
                                                                                                 op_kronahX_2_1_r}));
  assign op_kronahX_2_destruct_r = (& op_kronahX_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_2_destruct_emitted <= 2'd0;
    else
      op_kronahX_2_destruct_emitted <= (op_kronahX_2_destruct_r ? 2'd0 :
                                        op_kronahX_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronahX_3_2,MyDTInt_Int_Int) > (op_kronahX_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronahX_3_2_bufchan_d;
  logic op_kronahX_3_2_bufchan_r;
  assign op_kronahX_3_2_r = ((! op_kronahX_3_2_bufchan_d[0]) || op_kronahX_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_3_2_bufchan_d <= 1'd0;
    else
      if (op_kronahX_3_2_r) op_kronahX_3_2_bufchan_d <= op_kronahX_3_2_d;
  MyDTInt_Int_Int_t op_kronahX_3_2_bufchan_buf;
  assign op_kronahX_3_2_bufchan_r = (! op_kronahX_3_2_bufchan_buf[0]);
  assign op_kronahX_3_2_argbuf_d = (op_kronahX_3_2_bufchan_buf[0] ? op_kronahX_3_2_bufchan_buf :
                                    op_kronahX_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_kronahX_3_2_argbuf_r && op_kronahX_3_2_bufchan_buf[0]))
        op_kronahX_3_2_bufchan_buf <= 1'd0;
      else if (((! op_kronahX_3_2_argbuf_r) && (! op_kronahX_3_2_bufchan_buf[0])))
        op_kronahX_3_2_bufchan_buf <= op_kronahX_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_kronahX_3_destruct,MyDTInt_Int_Int) > [(op_kronahX_3_1,MyDTInt_Int_Int),
                                                                       (op_kronahX_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_kronahX_3_destruct_emitted;
  logic [1:0] op_kronahX_3_destruct_done;
  assign op_kronahX_3_1_d = (op_kronahX_3_destruct_d[0] && (! op_kronahX_3_destruct_emitted[0]));
  assign op_kronahX_3_2_d = (op_kronahX_3_destruct_d[0] && (! op_kronahX_3_destruct_emitted[1]));
  assign op_kronahX_3_destruct_done = (op_kronahX_3_destruct_emitted | ({op_kronahX_3_2_d[0],
                                                                         op_kronahX_3_1_d[0]} & {op_kronahX_3_2_r,
                                                                                                 op_kronahX_3_1_r}));
  assign op_kronahX_3_destruct_r = (& op_kronahX_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_3_destruct_emitted <= 2'd0;
    else
      op_kronahX_3_destruct_emitted <= (op_kronahX_3_destruct_r ? 2'd0 :
                                        op_kronahX_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronahX_4_destruct,MyDTInt_Int_Int) > (op_kronahX_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronahX_4_destruct_bufchan_d;
  logic op_kronahX_4_destruct_bufchan_r;
  assign op_kronahX_4_destruct_r = ((! op_kronahX_4_destruct_bufchan_d[0]) || op_kronahX_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_kronahX_4_destruct_r)
        op_kronahX_4_destruct_bufchan_d <= op_kronahX_4_destruct_d;
  MyDTInt_Int_Int_t op_kronahX_4_destruct_bufchan_buf;
  assign op_kronahX_4_destruct_bufchan_r = (! op_kronahX_4_destruct_bufchan_buf[0]);
  assign op_kronahX_4_1_argbuf_d = (op_kronahX_4_destruct_bufchan_buf[0] ? op_kronahX_4_destruct_bufchan_buf :
                                    op_kronahX_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronahX_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_kronahX_4_1_argbuf_r && op_kronahX_4_destruct_bufchan_buf[0]))
        op_kronahX_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_kronahX_4_1_argbuf_r) && (! op_kronahX_4_destruct_bufchan_buf[0])))
        op_kronahX_4_destruct_bufchan_buf <= op_kronahX_4_destruct_bufchan_d;
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronai7_2_2,MyDTInt_Int_Int) > (op_kronai7_2_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronai7_2_2_bufchan_d;
  logic op_kronai7_2_2_bufchan_r;
  assign op_kronai7_2_2_r = ((! op_kronai7_2_2_bufchan_d[0]) || op_kronai7_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_2_2_bufchan_d <= 1'd0;
    else
      if (op_kronai7_2_2_r) op_kronai7_2_2_bufchan_d <= op_kronai7_2_2_d;
  MyDTInt_Int_Int_t op_kronai7_2_2_bufchan_buf;
  assign op_kronai7_2_2_bufchan_r = (! op_kronai7_2_2_bufchan_buf[0]);
  assign op_kronai7_2_2_argbuf_d = (op_kronai7_2_2_bufchan_buf[0] ? op_kronai7_2_2_bufchan_buf :
                                    op_kronai7_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_2_2_bufchan_buf <= 1'd0;
    else
      if ((op_kronai7_2_2_argbuf_r && op_kronai7_2_2_bufchan_buf[0]))
        op_kronai7_2_2_bufchan_buf <= 1'd0;
      else if (((! op_kronai7_2_2_argbuf_r) && (! op_kronai7_2_2_bufchan_buf[0])))
        op_kronai7_2_2_bufchan_buf <= op_kronai7_2_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_kronai7_2_destruct,MyDTInt_Int_Int) > [(op_kronai7_2_1,MyDTInt_Int_Int),
                                                                       (op_kronai7_2_2,MyDTInt_Int_Int)] */
  logic [1:0] op_kronai7_2_destruct_emitted;
  logic [1:0] op_kronai7_2_destruct_done;
  assign op_kronai7_2_1_d = (op_kronai7_2_destruct_d[0] && (! op_kronai7_2_destruct_emitted[0]));
  assign op_kronai7_2_2_d = (op_kronai7_2_destruct_d[0] && (! op_kronai7_2_destruct_emitted[1]));
  assign op_kronai7_2_destruct_done = (op_kronai7_2_destruct_emitted | ({op_kronai7_2_2_d[0],
                                                                         op_kronai7_2_1_d[0]} & {op_kronai7_2_2_r,
                                                                                                 op_kronai7_2_1_r}));
  assign op_kronai7_2_destruct_r = (& op_kronai7_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_2_destruct_emitted <= 2'd0;
    else
      op_kronai7_2_destruct_emitted <= (op_kronai7_2_destruct_r ? 2'd0 :
                                        op_kronai7_2_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronai7_3_2,MyDTInt_Int_Int) > (op_kronai7_3_2_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronai7_3_2_bufchan_d;
  logic op_kronai7_3_2_bufchan_r;
  assign op_kronai7_3_2_r = ((! op_kronai7_3_2_bufchan_d[0]) || op_kronai7_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_3_2_bufchan_d <= 1'd0;
    else
      if (op_kronai7_3_2_r) op_kronai7_3_2_bufchan_d <= op_kronai7_3_2_d;
  MyDTInt_Int_Int_t op_kronai7_3_2_bufchan_buf;
  assign op_kronai7_3_2_bufchan_r = (! op_kronai7_3_2_bufchan_buf[0]);
  assign op_kronai7_3_2_argbuf_d = (op_kronai7_3_2_bufchan_buf[0] ? op_kronai7_3_2_bufchan_buf :
                                    op_kronai7_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_3_2_bufchan_buf <= 1'd0;
    else
      if ((op_kronai7_3_2_argbuf_r && op_kronai7_3_2_bufchan_buf[0]))
        op_kronai7_3_2_bufchan_buf <= 1'd0;
      else if (((! op_kronai7_3_2_argbuf_r) && (! op_kronai7_3_2_bufchan_buf[0])))
        op_kronai7_3_2_bufchan_buf <= op_kronai7_3_2_bufchan_d;
  
  /* fork (Ty MyDTInt_Int_Int) : (op_kronai7_3_destruct,MyDTInt_Int_Int) > [(op_kronai7_3_1,MyDTInt_Int_Int),
                                                                       (op_kronai7_3_2,MyDTInt_Int_Int)] */
  logic [1:0] op_kronai7_3_destruct_emitted;
  logic [1:0] op_kronai7_3_destruct_done;
  assign op_kronai7_3_1_d = (op_kronai7_3_destruct_d[0] && (! op_kronai7_3_destruct_emitted[0]));
  assign op_kronai7_3_2_d = (op_kronai7_3_destruct_d[0] && (! op_kronai7_3_destruct_emitted[1]));
  assign op_kronai7_3_destruct_done = (op_kronai7_3_destruct_emitted | ({op_kronai7_3_2_d[0],
                                                                         op_kronai7_3_1_d[0]} & {op_kronai7_3_2_r,
                                                                                                 op_kronai7_3_1_r}));
  assign op_kronai7_3_destruct_r = (& op_kronai7_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_3_destruct_emitted <= 2'd0;
    else
      op_kronai7_3_destruct_emitted <= (op_kronai7_3_destruct_r ? 2'd0 :
                                        op_kronai7_3_destruct_done);
  
  /* buf (Ty MyDTInt_Int_Int) : (op_kronai7_4_destruct,MyDTInt_Int_Int) > (op_kronai7_4_1_argbuf,MyDTInt_Int_Int) */
  MyDTInt_Int_Int_t op_kronai7_4_destruct_bufchan_d;
  logic op_kronai7_4_destruct_bufchan_r;
  assign op_kronai7_4_destruct_r = ((! op_kronai7_4_destruct_bufchan_d[0]) || op_kronai7_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_4_destruct_bufchan_d <= 1'd0;
    else
      if (op_kronai7_4_destruct_r)
        op_kronai7_4_destruct_bufchan_d <= op_kronai7_4_destruct_d;
  MyDTInt_Int_Int_t op_kronai7_4_destruct_bufchan_buf;
  assign op_kronai7_4_destruct_bufchan_r = (! op_kronai7_4_destruct_bufchan_buf[0]);
  assign op_kronai7_4_1_argbuf_d = (op_kronai7_4_destruct_bufchan_buf[0] ? op_kronai7_4_destruct_bufchan_buf :
                                    op_kronai7_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) op_kronai7_4_destruct_bufchan_buf <= 1'd0;
    else
      if ((op_kronai7_4_1_argbuf_r && op_kronai7_4_destruct_bufchan_buf[0]))
        op_kronai7_4_destruct_bufchan_buf <= 1'd0;
      else if (((! op_kronai7_4_1_argbuf_r) && (! op_kronai7_4_destruct_bufchan_buf[0])))
        op_kronai7_4_destruct_bufchan_buf <= op_kronai7_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1abW_destruct,Pointer_QTree_Int) > (q1abW_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1abW_destruct_bufchan_d;
  logic q1abW_destruct_bufchan_r;
  assign q1abW_destruct_r = ((! q1abW_destruct_bufchan_d[0]) || q1abW_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1abW_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1abW_destruct_r) q1abW_destruct_bufchan_d <= q1abW_destruct_d;
  Pointer_QTree_Int_t q1abW_destruct_bufchan_buf;
  assign q1abW_destruct_bufchan_r = (! q1abW_destruct_bufchan_buf[0]);
  assign q1abW_1_argbuf_d = (q1abW_destruct_bufchan_buf[0] ? q1abW_destruct_bufchan_buf :
                             q1abW_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1abW_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1abW_1_argbuf_r && q1abW_destruct_bufchan_buf[0]))
        q1abW_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1abW_1_argbuf_r) && (! q1abW_destruct_bufchan_buf[0])))
        q1abW_destruct_bufchan_buf <= q1abW_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1ai1_3_destruct,Pointer_QTree_Int) > (q1ai1_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1ai1_3_destruct_bufchan_d;
  logic q1ai1_3_destruct_bufchan_r;
  assign q1ai1_3_destruct_r = ((! q1ai1_3_destruct_bufchan_d[0]) || q1ai1_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ai1_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1ai1_3_destruct_r)
        q1ai1_3_destruct_bufchan_d <= q1ai1_3_destruct_d;
  Pointer_QTree_Int_t q1ai1_3_destruct_bufchan_buf;
  assign q1ai1_3_destruct_bufchan_r = (! q1ai1_3_destruct_bufchan_buf[0]);
  assign q1ai1_3_1_argbuf_d = (q1ai1_3_destruct_bufchan_buf[0] ? q1ai1_3_destruct_bufchan_buf :
                               q1ai1_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1ai1_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1ai1_3_1_argbuf_r && q1ai1_3_destruct_bufchan_buf[0]))
        q1ai1_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1ai1_3_1_argbuf_r) && (! q1ai1_3_destruct_bufchan_buf[0])))
        q1ai1_3_destruct_bufchan_buf <= q1ai1_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q1aic_3_destruct,Pointer_QTree_Int) > (q1aic_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q1aic_3_destruct_bufchan_d;
  logic q1aic_3_destruct_bufchan_r;
  assign q1aic_3_destruct_r = ((! q1aic_3_destruct_bufchan_d[0]) || q1aic_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aic_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q1aic_3_destruct_r)
        q1aic_3_destruct_bufchan_d <= q1aic_3_destruct_d;
  Pointer_QTree_Int_t q1aic_3_destruct_bufchan_buf;
  assign q1aic_3_destruct_bufchan_r = (! q1aic_3_destruct_bufchan_buf[0]);
  assign q1aic_3_1_argbuf_d = (q1aic_3_destruct_bufchan_buf[0] ? q1aic_3_destruct_bufchan_buf :
                               q1aic_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q1aic_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q1aic_3_1_argbuf_r && q1aic_3_destruct_bufchan_buf[0]))
        q1aic_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q1aic_3_1_argbuf_r) && (! q1aic_3_destruct_bufchan_buf[0])))
        q1aic_3_destruct_bufchan_buf <= q1aic_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2abX_1_destruct,Pointer_QTree_Int) > (q2abX_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2abX_1_destruct_bufchan_d;
  logic q2abX_1_destruct_bufchan_r;
  assign q2abX_1_destruct_r = ((! q2abX_1_destruct_bufchan_d[0]) || q2abX_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2abX_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2abX_1_destruct_r)
        q2abX_1_destruct_bufchan_d <= q2abX_1_destruct_d;
  Pointer_QTree_Int_t q2abX_1_destruct_bufchan_buf;
  assign q2abX_1_destruct_bufchan_r = (! q2abX_1_destruct_bufchan_buf[0]);
  assign q2abX_1_1_argbuf_d = (q2abX_1_destruct_bufchan_buf[0] ? q2abX_1_destruct_bufchan_buf :
                               q2abX_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2abX_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2abX_1_1_argbuf_r && q2abX_1_destruct_bufchan_buf[0]))
        q2abX_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2abX_1_1_argbuf_r) && (! q2abX_1_destruct_bufchan_buf[0])))
        q2abX_1_destruct_bufchan_buf <= q2abX_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2ai2_2_destruct,Pointer_QTree_Int) > (q2ai2_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2ai2_2_destruct_bufchan_d;
  logic q2ai2_2_destruct_bufchan_r;
  assign q2ai2_2_destruct_r = ((! q2ai2_2_destruct_bufchan_d[0]) || q2ai2_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ai2_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2ai2_2_destruct_r)
        q2ai2_2_destruct_bufchan_d <= q2ai2_2_destruct_d;
  Pointer_QTree_Int_t q2ai2_2_destruct_bufchan_buf;
  assign q2ai2_2_destruct_bufchan_r = (! q2ai2_2_destruct_bufchan_buf[0]);
  assign q2ai2_2_1_argbuf_d = (q2ai2_2_destruct_bufchan_buf[0] ? q2ai2_2_destruct_bufchan_buf :
                               q2ai2_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2ai2_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2ai2_2_1_argbuf_r && q2ai2_2_destruct_bufchan_buf[0]))
        q2ai2_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2ai2_2_1_argbuf_r) && (! q2ai2_2_destruct_bufchan_buf[0])))
        q2ai2_2_destruct_bufchan_buf <= q2ai2_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q2aid_2_destruct,Pointer_QTree_Int) > (q2aid_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q2aid_2_destruct_bufchan_d;
  logic q2aid_2_destruct_bufchan_r;
  assign q2aid_2_destruct_r = ((! q2aid_2_destruct_bufchan_d[0]) || q2aid_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aid_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q2aid_2_destruct_r)
        q2aid_2_destruct_bufchan_d <= q2aid_2_destruct_d;
  Pointer_QTree_Int_t q2aid_2_destruct_bufchan_buf;
  assign q2aid_2_destruct_bufchan_r = (! q2aid_2_destruct_bufchan_buf[0]);
  assign q2aid_2_1_argbuf_d = (q2aid_2_destruct_bufchan_buf[0] ? q2aid_2_destruct_bufchan_buf :
                               q2aid_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q2aid_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q2aid_2_1_argbuf_r && q2aid_2_destruct_bufchan_buf[0]))
        q2aid_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q2aid_2_1_argbuf_r) && (! q2aid_2_destruct_bufchan_buf[0])))
        q2aid_2_destruct_bufchan_buf <= q2aid_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3abY_2_destruct,Pointer_QTree_Int) > (q3abY_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3abY_2_destruct_bufchan_d;
  logic q3abY_2_destruct_bufchan_r;
  assign q3abY_2_destruct_r = ((! q3abY_2_destruct_bufchan_d[0]) || q3abY_2_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3abY_2_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3abY_2_destruct_r)
        q3abY_2_destruct_bufchan_d <= q3abY_2_destruct_d;
  Pointer_QTree_Int_t q3abY_2_destruct_bufchan_buf;
  assign q3abY_2_destruct_bufchan_r = (! q3abY_2_destruct_bufchan_buf[0]);
  assign q3abY_2_1_argbuf_d = (q3abY_2_destruct_bufchan_buf[0] ? q3abY_2_destruct_bufchan_buf :
                               q3abY_2_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3abY_2_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3abY_2_1_argbuf_r && q3abY_2_destruct_bufchan_buf[0]))
        q3abY_2_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3abY_2_1_argbuf_r) && (! q3abY_2_destruct_bufchan_buf[0])))
        q3abY_2_destruct_bufchan_buf <= q3abY_2_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3ai3_1_destruct,Pointer_QTree_Int) > (q3ai3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3ai3_1_destruct_bufchan_d;
  logic q3ai3_1_destruct_bufchan_r;
  assign q3ai3_1_destruct_r = ((! q3ai3_1_destruct_bufchan_d[0]) || q3ai3_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ai3_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3ai3_1_destruct_r)
        q3ai3_1_destruct_bufchan_d <= q3ai3_1_destruct_d;
  Pointer_QTree_Int_t q3ai3_1_destruct_bufchan_buf;
  assign q3ai3_1_destruct_bufchan_r = (! q3ai3_1_destruct_bufchan_buf[0]);
  assign q3ai3_1_1_argbuf_d = (q3ai3_1_destruct_bufchan_buf[0] ? q3ai3_1_destruct_bufchan_buf :
                               q3ai3_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3ai3_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3ai3_1_1_argbuf_r && q3ai3_1_destruct_bufchan_buf[0]))
        q3ai3_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3ai3_1_1_argbuf_r) && (! q3ai3_1_destruct_bufchan_buf[0])))
        q3ai3_1_destruct_bufchan_buf <= q3ai3_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q3aie_1_destruct,Pointer_QTree_Int) > (q3aie_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q3aie_1_destruct_bufchan_d;
  logic q3aie_1_destruct_bufchan_r;
  assign q3aie_1_destruct_r = ((! q3aie_1_destruct_bufchan_d[0]) || q3aie_1_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aie_1_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q3aie_1_destruct_r)
        q3aie_1_destruct_bufchan_d <= q3aie_1_destruct_d;
  Pointer_QTree_Int_t q3aie_1_destruct_bufchan_buf;
  assign q3aie_1_destruct_bufchan_r = (! q3aie_1_destruct_bufchan_buf[0]);
  assign q3aie_1_1_argbuf_d = (q3aie_1_destruct_bufchan_buf[0] ? q3aie_1_destruct_bufchan_buf :
                               q3aie_1_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q3aie_1_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q3aie_1_1_argbuf_r && q3aie_1_destruct_bufchan_buf[0]))
        q3aie_1_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q3aie_1_1_argbuf_r) && (! q3aie_1_destruct_bufchan_buf[0])))
        q3aie_1_destruct_bufchan_buf <= q3aie_1_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4abZ_3_destruct,Pointer_QTree_Int) > (q4abZ_3_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4abZ_3_destruct_bufchan_d;
  logic q4abZ_3_destruct_bufchan_r;
  assign q4abZ_3_destruct_r = ((! q4abZ_3_destruct_bufchan_d[0]) || q4abZ_3_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4abZ_3_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4abZ_3_destruct_r)
        q4abZ_3_destruct_bufchan_d <= q4abZ_3_destruct_d;
  Pointer_QTree_Int_t q4abZ_3_destruct_bufchan_buf;
  assign q4abZ_3_destruct_bufchan_r = (! q4abZ_3_destruct_bufchan_buf[0]);
  assign q4abZ_3_1_argbuf_d = (q4abZ_3_destruct_bufchan_buf[0] ? q4abZ_3_destruct_bufchan_buf :
                               q4abZ_3_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4abZ_3_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4abZ_3_1_argbuf_r && q4abZ_3_destruct_bufchan_buf[0]))
        q4abZ_3_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4abZ_3_1_argbuf_r) && (! q4abZ_3_destruct_bufchan_buf[0])))
        q4abZ_3_destruct_bufchan_buf <= q4abZ_3_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4ai4_destruct,Pointer_QTree_Int) > (q4ai4_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4ai4_destruct_bufchan_d;
  logic q4ai4_destruct_bufchan_r;
  assign q4ai4_destruct_r = ((! q4ai4_destruct_bufchan_d[0]) || q4ai4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ai4_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4ai4_destruct_r) q4ai4_destruct_bufchan_d <= q4ai4_destruct_d;
  Pointer_QTree_Int_t q4ai4_destruct_bufchan_buf;
  assign q4ai4_destruct_bufchan_r = (! q4ai4_destruct_bufchan_buf[0]);
  assign q4ai4_1_argbuf_d = (q4ai4_destruct_bufchan_buf[0] ? q4ai4_destruct_bufchan_buf :
                             q4ai4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4ai4_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4ai4_1_argbuf_r && q4ai4_destruct_bufchan_buf[0]))
        q4ai4_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4ai4_1_argbuf_r) && (! q4ai4_destruct_bufchan_buf[0])))
        q4ai4_destruct_bufchan_buf <= q4ai4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (q4aif_destruct,Pointer_QTree_Int) > (q4aif_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t q4aif_destruct_bufchan_d;
  logic q4aif_destruct_bufchan_r;
  assign q4aif_destruct_r = ((! q4aif_destruct_bufchan_d[0]) || q4aif_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4aif_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (q4aif_destruct_r) q4aif_destruct_bufchan_d <= q4aif_destruct_d;
  Pointer_QTree_Int_t q4aif_destruct_bufchan_buf;
  assign q4aif_destruct_bufchan_r = (! q4aif_destruct_bufchan_buf[0]);
  assign q4aif_1_argbuf_d = (q4aif_destruct_bufchan_buf[0] ? q4aif_destruct_bufchan_buf :
                             q4aif_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) q4aif_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((q4aif_1_argbuf_r && q4aif_destruct_bufchan_buf[0]))
        q4aif_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! q4aif_1_argbuf_r) && (! q4aif_destruct_bufchan_buf[0])))
        q4aif_destruct_bufchan_buf <= q4aif_destruct_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf,CT$wnnz_Int) > (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) */
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  logic readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r = ((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d[0]) || readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= {115'd0,
                                                             1'd0};
    else
      if (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_r)
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_d;
  CT$wnnz_Int_t readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf;
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_r = (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]);
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0] ? readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf :
                                                           readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                               1'd0};
    else
      if ((readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r && readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0]))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= {115'd0,
                                                                 1'd0};
      else if (((! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r) && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf[0])))
        readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_buf <= readPointer_CT$wnnz_Intscfarg_0_1_argbuf_bufchan_d;
  
  /* fork (Ty CT$wnnz_Int) : (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb,CT$wnnz_Int) > [(lizzieLet19_1,CT$wnnz_Int),
                                                                                      (lizzieLet19_2,CT$wnnz_Int),
                                                                                      (lizzieLet19_3,CT$wnnz_Int),
                                                                                      (lizzieLet19_4,CT$wnnz_Int)] */
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done;
  assign lizzieLet19_1_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet19_2_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet19_3_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet19_4_d = {readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[115:1],
                            (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_d[0] && (! readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done = (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted | ({lizzieLet19_4_d[0],
                                                                                                                       lizzieLet19_3_d[0],
                                                                                                                       lizzieLet19_2_d[0],
                                                                                                                       lizzieLet19_1_d[0]} & {lizzieLet19_4_r,
                                                                                                                                              lizzieLet19_3_r,
                                                                                                                                              lizzieLet19_2_r,
                                                                                                                                              lizzieLet19_1_r}));
  assign readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r = (& readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_emitted <= (readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_r ? 4'd0 :
                                                               readPointer_CT$wnnz_Intscfarg_0_1_argbuf_rwb_done);
  
  /* buf (Ty CTf'_f'_Int_Int_Int_Int) : (readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf,CTf'_f'_Int_Int_Int_Int) > (readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTf'_f'_Int_Int_Int_Int) */
  \CTf'_f'_Int_Int_Int_Int_t  \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d ;
  logic \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r ;
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_r  = ((! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d [0]) || \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d  <= {99'd0,
                                                                             1'd0};
    else
      if (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_r )
        \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d  <= \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_d ;
  \CTf'_f'_Int_Int_Int_Int_t  \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf ;
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_r  = (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0]);
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d  = (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0] ? \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  :
                                                                           \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {99'd0,
                                                                               1'd0};
    else
      if ((\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r  && \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0]))
        \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= {99'd0,
                                                                                 1'd0};
      else if (((! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r ) && (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf [0])))
        \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_buf  <= \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_bufchan_d ;
  
  /* fork (Ty CTf'_f'_Int_Int_Int_Int) : (readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb,CTf'_f'_Int_Int_Int_Int) > [(lizzieLet23_1,CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet23_2,CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet23_3,CTf'_f'_Int_Int_Int_Int),
                                                                                                                            (lizzieLet23_4,CTf'_f'_Int_Int_Int_Int)] */
  logic [3:0] \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted ;
  logic [3:0] \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done ;
  assign lizzieLet23_1_d = {\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [0]))};
  assign lizzieLet23_2_d = {\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [1]))};
  assign lizzieLet23_3_d = {\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [2]))};
  assign lizzieLet23_4_d = {\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [99:1],
                            (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_d [0] && (! \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted [3]))};
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done  = (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  | ({lizzieLet23_4_d[0],
                                                                                                                                                       lizzieLet23_3_d[0],
                                                                                                                                                       lizzieLet23_2_d[0],
                                                                                                                                                       lizzieLet23_1_d[0]} & {lizzieLet23_4_r,
                                                                                                                                                                              lizzieLet23_3_r,
                                                                                                                                                                              lizzieLet23_2_r,
                                                                                                                                                                              lizzieLet23_1_r}));
  assign \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r  = (& \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  <= 4'd0;
    else
      \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_emitted  <= (\readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_r  ? 4'd0 :
                                                                               \readPointer_CTf'_f'_Int_Int_Int_Intscfarg_0_1_1_argbuf_rwb_done );
  
  /* buf (Ty CTf_f_Int_Int_Int_Int) : (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf,CTf_f_Int_Int_Int_Int) > (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int_Int_Int_Int) */
  CTf_f_Int_Int_Int_Int_t readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d;
  logic readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_r;
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_r = ((! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d[0]) || readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d <= {83'd0,
                                                                         1'd0};
    else
      if (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_r)
        readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d <= readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_d;
  CTf_f_Int_Int_Int_Int_t readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf;
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_r = (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0]);
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d = (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0] ? readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf :
                                                                       readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= {83'd0,
                                                                           1'd0};
    else
      if ((readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_r && readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0]))
        readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= {83'd0,
                                                                             1'd0};
      else if (((! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_r) && (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf[0])))
        readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_buf <= readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_bufchan_d;
  
  /* fork (Ty CTf_f_Int_Int_Int_Int) : (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb,CTf_f_Int_Int_Int_Int) > [(lizzieLet28_1,CTf_f_Int_Int_Int_Int),
                                                                                                                      (lizzieLet28_2,CTf_f_Int_Int_Int_Int),
                                                                                                                      (lizzieLet28_3,CTf_f_Int_Int_Int_Int),
                                                                                                                      (lizzieLet28_4,CTf_f_Int_Int_Int_Int)] */
  logic [3:0] readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_done;
  assign lizzieLet28_1_d = {readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[83:1],
                            (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet28_2_d = {readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[83:1],
                            (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet28_3_d = {readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[83:1],
                            (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet28_4_d = {readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[83:1],
                            (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_d[0] && (! readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted[3]))};
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_done = (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted | ({lizzieLet28_4_d[0],
                                                                                                                                               lizzieLet28_3_d[0],
                                                                                                                                               lizzieLet28_2_d[0],
                                                                                                                                               lizzieLet28_1_d[0]} & {lizzieLet28_4_r,
                                                                                                                                                                      lizzieLet28_3_r,
                                                                                                                                                                      lizzieLet28_2_r,
                                                                                                                                                                      lizzieLet28_1_r}));
  assign readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_r = (& readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_emitted <= (readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_r ? 4'd0 :
                                                                           readPointer_CTf_f_Int_Int_Int_Intscfarg_0_2_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm1ahU_1_argbuf,QTree_Int) > (readPointer_QTree_Intm1ahU_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm1ahU_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm1ahU_1_argbuf_r = ((! readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm1ahU_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm1ahU_1_argbuf_r)
        readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d <= readPointer_QTree_Intm1ahU_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm1ahU_1_argbuf_bufchan_r = (! readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm1ahU_1_argbuf_rwb_d = (readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm1ahU_1_argbuf_rwb_r && readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm1ahU_1_argbuf_rwb_r) && (! readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm1ahU_1_argbuf_bufchan_buf <= readPointer_QTree_Intm1ahU_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm1ahU_1_argbuf_rwb,QTree_Int) > [(lizzieLet13_1_1,QTree_Int),
                                                                             (lizzieLet13_1_2,QTree_Int),
                                                                             (lizzieLet13_1_3,QTree_Int),
                                                                             (lizzieLet13_1_4,QTree_Int),
                                                                             (lizzieLet13_1_5,QTree_Int),
                                                                             (lizzieLet13_1_6,QTree_Int),
                                                                             (lizzieLet13_1_7,QTree_Int),
                                                                             (lizzieLet13_1_8,QTree_Int),
                                                                             (lizzieLet13_1_9,QTree_Int)] */
  logic [8:0] readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Intm1ahU_1_argbuf_rwb_done;
  assign lizzieLet13_1_1_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet13_1_2_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet13_1_3_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet13_1_4_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet13_1_5_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet13_1_6_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet13_1_7_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet13_1_8_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet13_1_9_d = {readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[66:1],
                              (readPointer_QTree_Intm1ahU_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Intm1ahU_1_argbuf_rwb_done = (readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted | ({lizzieLet13_1_9_d[0],
                                                                                                             lizzieLet13_1_8_d[0],
                                                                                                             lizzieLet13_1_7_d[0],
                                                                                                             lizzieLet13_1_6_d[0],
                                                                                                             lizzieLet13_1_5_d[0],
                                                                                                             lizzieLet13_1_4_d[0],
                                                                                                             lizzieLet13_1_3_d[0],
                                                                                                             lizzieLet13_1_2_d[0],
                                                                                                             lizzieLet13_1_1_d[0]} & {lizzieLet13_1_9_r,
                                                                                                                                      lizzieLet13_1_8_r,
                                                                                                                                      lizzieLet13_1_7_r,
                                                                                                                                      lizzieLet13_1_6_r,
                                                                                                                                      lizzieLet13_1_5_r,
                                                                                                                                      lizzieLet13_1_4_r,
                                                                                                                                      lizzieLet13_1_3_r,
                                                                                                                                      lizzieLet13_1_2_r,
                                                                                                                                      lizzieLet13_1_1_r}));
  assign readPointer_QTree_Intm1ahU_1_argbuf_rwb_r = (& readPointer_QTree_Intm1ahU_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Intm1ahU_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm1ahU_1_argbuf_rwb_r ? 9'd0 :
                                                          readPointer_QTree_Intm1ahU_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_Intm2ai5_1_argbuf,QTree_Int) > (readPointer_QTree_Intm2ai5_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d;
  logic readPointer_QTree_Intm2ai5_1_argbuf_bufchan_r;
  assign readPointer_QTree_Intm2ai5_1_argbuf_r = ((! readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d[0]) || readPointer_QTree_Intm2ai5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_Intm2ai5_1_argbuf_r)
        readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d <= readPointer_QTree_Intm2ai5_1_argbuf_d;
  QTree_Int_t readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf;
  assign readPointer_QTree_Intm2ai5_1_argbuf_bufchan_r = (! readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_Intm2ai5_1_argbuf_rwb_d = (readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf[0] ? readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf :
                                                      readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_Intm2ai5_1_argbuf_rwb_r && readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_Intm2ai5_1_argbuf_rwb_r) && (! readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_Intm2ai5_1_argbuf_bufchan_buf <= readPointer_QTree_Intm2ai5_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_Intm2ai5_1_argbuf_rwb,QTree_Int) > [(lizzieLet6_1,QTree_Int),
                                                                             (lizzieLet6_2,QTree_Int),
                                                                             (lizzieLet6_3,QTree_Int),
                                                                             (lizzieLet6_4,QTree_Int),
                                                                             (lizzieLet6_5,QTree_Int),
                                                                             (lizzieLet6_6,QTree_Int),
                                                                             (lizzieLet6_7,QTree_Int),
                                                                             (lizzieLet6_8,QTree_Int),
                                                                             (lizzieLet6_9,QTree_Int)] */
  logic [8:0] readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted;
  logic [8:0] readPointer_QTree_Intm2ai5_1_argbuf_rwb_done;
  assign lizzieLet6_1_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet6_2_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet6_3_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet6_4_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[3]))};
  assign lizzieLet6_5_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[4]))};
  assign lizzieLet6_6_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[5]))};
  assign lizzieLet6_7_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[6]))};
  assign lizzieLet6_8_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[7]))};
  assign lizzieLet6_9_d = {readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_Intm2ai5_1_argbuf_rwb_d[0] && (! readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted[8]))};
  assign readPointer_QTree_Intm2ai5_1_argbuf_rwb_done = (readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted | ({lizzieLet6_9_d[0],
                                                                                                             lizzieLet6_8_d[0],
                                                                                                             lizzieLet6_7_d[0],
                                                                                                             lizzieLet6_6_d[0],
                                                                                                             lizzieLet6_5_d[0],
                                                                                                             lizzieLet6_4_d[0],
                                                                                                             lizzieLet6_3_d[0],
                                                                                                             lizzieLet6_2_d[0],
                                                                                                             lizzieLet6_1_d[0]} & {lizzieLet6_9_r,
                                                                                                                                   lizzieLet6_8_r,
                                                                                                                                   lizzieLet6_7_r,
                                                                                                                                   lizzieLet6_6_r,
                                                                                                                                   lizzieLet6_5_r,
                                                                                                                                   lizzieLet6_4_r,
                                                                                                                                   lizzieLet6_3_r,
                                                                                                                                   lizzieLet6_2_r,
                                                                                                                                   lizzieLet6_1_r}));
  assign readPointer_QTree_Intm2ai5_1_argbuf_rwb_r = (& readPointer_QTree_Intm2ai5_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted <= 9'd0;
    else
      readPointer_QTree_Intm2ai5_1_argbuf_rwb_emitted <= (readPointer_QTree_Intm2ai5_1_argbuf_rwb_r ? 9'd0 :
                                                          readPointer_QTree_Intm2ai5_1_argbuf_rwb_done);
  
  /* buf (Ty QTree_Int) : (readPointer_QTree_IntwstH_1_1_argbuf,QTree_Int) > (readPointer_QTree_IntwstH_1_1_argbuf_rwb,QTree_Int) */
  QTree_Int_t readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d;
  logic readPointer_QTree_IntwstH_1_1_argbuf_bufchan_r;
  assign readPointer_QTree_IntwstH_1_1_argbuf_r = ((! readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d[0]) || readPointer_QTree_IntwstH_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d <= {66'd0, 1'd0};
    else
      if (readPointer_QTree_IntwstH_1_1_argbuf_r)
        readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d <= readPointer_QTree_IntwstH_1_1_argbuf_d;
  QTree_Int_t readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf;
  assign readPointer_QTree_IntwstH_1_1_argbuf_bufchan_r = (! readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf[0]);
  assign readPointer_QTree_IntwstH_1_1_argbuf_rwb_d = (readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf[0] ? readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf :
                                                       readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
    else
      if ((readPointer_QTree_IntwstH_1_1_argbuf_rwb_r && readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf[0]))
        readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf <= {66'd0, 1'd0};
      else if (((! readPointer_QTree_IntwstH_1_1_argbuf_rwb_r) && (! readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf[0])))
        readPointer_QTree_IntwstH_1_1_argbuf_bufchan_buf <= readPointer_QTree_IntwstH_1_1_argbuf_bufchan_d;
  
  /* fork (Ty QTree_Int) : (readPointer_QTree_IntwstH_1_1_argbuf_rwb,QTree_Int) > [(lizzieLet4_1,QTree_Int),
                                                                              (lizzieLet4_2,QTree_Int),
                                                                              (lizzieLet4_3,QTree_Int),
                                                                              (lizzieLet4_4,QTree_Int)] */
  logic [3:0] readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted;
  logic [3:0] readPointer_QTree_IntwstH_1_1_argbuf_rwb_done;
  assign lizzieLet4_1_d = {readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted[0]))};
  assign lizzieLet4_2_d = {readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted[1]))};
  assign lizzieLet4_3_d = {readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted[2]))};
  assign lizzieLet4_4_d = {readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[66:1],
                           (readPointer_QTree_IntwstH_1_1_argbuf_rwb_d[0] && (! readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted[3]))};
  assign readPointer_QTree_IntwstH_1_1_argbuf_rwb_done = (readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted | ({lizzieLet4_4_d[0],
                                                                                                               lizzieLet4_3_d[0],
                                                                                                               lizzieLet4_2_d[0],
                                                                                                               lizzieLet4_1_d[0]} & {lizzieLet4_4_r,
                                                                                                                                     lizzieLet4_3_r,
                                                                                                                                     lizzieLet4_2_r,
                                                                                                                                     lizzieLet4_1_r}));
  assign readPointer_QTree_IntwstH_1_1_argbuf_rwb_r = (& readPointer_QTree_IntwstH_1_1_argbuf_rwb_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted <= 4'd0;
    else
      readPointer_QTree_IntwstH_1_1_argbuf_rwb_emitted <= (readPointer_QTree_IntwstH_1_1_argbuf_rwb_r ? 4'd0 :
                                                           readPointer_QTree_IntwstH_1_1_argbuf_rwb_done);
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (sc_0_10_destruct,Pointer_CTf'_f'_Int_Int_Int_Int) > (sc_0_10_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_10_destruct_bufchan_d;
  logic sc_0_10_destruct_bufchan_r;
  assign sc_0_10_destruct_r = ((! sc_0_10_destruct_bufchan_d[0]) || sc_0_10_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_10_destruct_r)
        sc_0_10_destruct_bufchan_d <= sc_0_10_destruct_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  sc_0_10_destruct_bufchan_buf;
  assign sc_0_10_destruct_bufchan_r = (! sc_0_10_destruct_bufchan_buf[0]);
  assign sc_0_10_1_argbuf_d = (sc_0_10_destruct_bufchan_buf[0] ? sc_0_10_destruct_bufchan_buf :
                               sc_0_10_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_10_1_argbuf_r && sc_0_10_destruct_bufchan_buf[0]))
        sc_0_10_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_10_1_argbuf_r) && (! sc_0_10_destruct_bufchan_buf[0])))
        sc_0_10_destruct_bufchan_buf <= sc_0_10_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (sc_0_14_destruct,Pointer_CTf_f_Int_Int_Int_Int) > (sc_0_14_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_14_destruct_bufchan_d;
  logic sc_0_14_destruct_bufchan_r;
  assign sc_0_14_destruct_r = ((! sc_0_14_destruct_bufchan_d[0]) || sc_0_14_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_14_destruct_r)
        sc_0_14_destruct_bufchan_d <= sc_0_14_destruct_d;
  Pointer_CTf_f_Int_Int_Int_Int_t sc_0_14_destruct_bufchan_buf;
  assign sc_0_14_destruct_bufchan_r = (! sc_0_14_destruct_bufchan_buf[0]);
  assign sc_0_14_1_argbuf_d = (sc_0_14_destruct_bufchan_buf[0] ? sc_0_14_destruct_bufchan_buf :
                               sc_0_14_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_14_1_argbuf_r && sc_0_14_destruct_bufchan_buf[0]))
        sc_0_14_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_14_1_argbuf_r) && (! sc_0_14_destruct_bufchan_buf[0])))
        sc_0_14_destruct_bufchan_buf <= sc_0_14_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (sc_0_6_destruct,Pointer_CT$wnnz_Int) > (sc_0_6_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_bufchan_d;
  logic sc_0_6_destruct_bufchan_r;
  assign sc_0_6_destruct_r = ((! sc_0_6_destruct_bufchan_d[0]) || sc_0_6_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_d <= {16'd0, 1'd0};
    else
      if (sc_0_6_destruct_r)
        sc_0_6_destruct_bufchan_d <= sc_0_6_destruct_d;
  Pointer_CT$wnnz_Int_t sc_0_6_destruct_bufchan_buf;
  assign sc_0_6_destruct_bufchan_r = (! sc_0_6_destruct_bufchan_buf[0]);
  assign sc_0_6_1_argbuf_d = (sc_0_6_destruct_bufchan_buf[0] ? sc_0_6_destruct_bufchan_buf :
                              sc_0_6_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((sc_0_6_1_argbuf_r && sc_0_6_destruct_bufchan_buf[0]))
        sc_0_6_destruct_bufchan_buf <= {16'd0, 1'd0};
      else if (((! sc_0_6_1_argbuf_r) && (! sc_0_6_destruct_bufchan_buf[0])))
        sc_0_6_destruct_bufchan_buf <= sc_0_6_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (scfarg_0_1_goMux_mux,Pointer_CTf'_f'_Int_Int_Int_Int) > (scfarg_0_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  scfarg_0_1_goMux_mux_bufchan_d;
  logic scfarg_0_1_goMux_mux_bufchan_r;
  assign scfarg_0_1_goMux_mux_r = ((! scfarg_0_1_goMux_mux_bufchan_d[0]) || scfarg_0_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_1_goMux_mux_r)
        scfarg_0_1_goMux_mux_bufchan_d <= scfarg_0_1_goMux_mux_d;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  scfarg_0_1_goMux_mux_bufchan_buf;
  assign scfarg_0_1_goMux_mux_bufchan_r = (! scfarg_0_1_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_1_argbuf_d = (scfarg_0_1_goMux_mux_bufchan_buf[0] ? scfarg_0_1_goMux_mux_bufchan_buf :
                                  scfarg_0_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_1_argbuf_r && scfarg_0_1_goMux_mux_bufchan_buf[0]))
        scfarg_0_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_1_argbuf_r) && (! scfarg_0_1_goMux_mux_bufchan_buf[0])))
        scfarg_0_1_goMux_mux_bufchan_buf <= scfarg_0_1_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (scfarg_0_2_goMux_mux,Pointer_CTf_f_Int_Int_Int_Int) > (scfarg_0_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t scfarg_0_2_goMux_mux_bufchan_d;
  logic scfarg_0_2_goMux_mux_bufchan_r;
  assign scfarg_0_2_goMux_mux_r = ((! scfarg_0_2_goMux_mux_bufchan_d[0]) || scfarg_0_2_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_2_goMux_mux_r)
        scfarg_0_2_goMux_mux_bufchan_d <= scfarg_0_2_goMux_mux_d;
  Pointer_CTf_f_Int_Int_Int_Int_t scfarg_0_2_goMux_mux_bufchan_buf;
  assign scfarg_0_2_goMux_mux_bufchan_r = (! scfarg_0_2_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_2_1_argbuf_d = (scfarg_0_2_goMux_mux_bufchan_buf[0] ? scfarg_0_2_goMux_mux_bufchan_buf :
                                  scfarg_0_2_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_2_1_argbuf_r && scfarg_0_2_goMux_mux_bufchan_buf[0]))
        scfarg_0_2_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_2_1_argbuf_r) && (! scfarg_0_2_goMux_mux_bufchan_buf[0])))
        scfarg_0_2_goMux_mux_bufchan_buf <= scfarg_0_2_goMux_mux_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (scfarg_0_goMux_mux,Pointer_CT$wnnz_Int) > (scfarg_0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_d;
  logic scfarg_0_goMux_mux_bufchan_r;
  assign scfarg_0_goMux_mux_r = ((! scfarg_0_goMux_mux_bufchan_d[0]) || scfarg_0_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) scfarg_0_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (scfarg_0_goMux_mux_r)
        scfarg_0_goMux_mux_bufchan_d <= scfarg_0_goMux_mux_d;
  Pointer_CT$wnnz_Int_t scfarg_0_goMux_mux_bufchan_buf;
  assign scfarg_0_goMux_mux_bufchan_r = (! scfarg_0_goMux_mux_bufchan_buf[0]);
  assign scfarg_0_1_argbuf_d = (scfarg_0_goMux_mux_bufchan_buf[0] ? scfarg_0_goMux_mux_bufchan_buf :
                                scfarg_0_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((scfarg_0_1_argbuf_r && scfarg_0_goMux_mux_bufchan_buf[0]))
        scfarg_0_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! scfarg_0_1_argbuf_r) && (! scfarg_0_goMux_mux_bufchan_buf[0])))
        scfarg_0_goMux_mux_bufchan_buf <= scfarg_0_goMux_mux_bufchan_d;
  
  /* buf (Ty Int) : (v'aib_1,Int) > (v'aib_1_argbuf,Int) */
  Int_t \v'aib_1_bufchan_d ;
  logic \v'aib_1_bufchan_r ;
  assign \v'aib_1_r  = ((! \v'aib_1_bufchan_d [0]) || \v'aib_1_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aib_1_bufchan_d  <= {32'd0, 1'd0};
    else if (\v'aib_1_r ) \v'aib_1_bufchan_d  <= \v'aib_1_d ;
  Int_t \v'aib_1_bufchan_buf ;
  assign \v'aib_1_bufchan_r  = (! \v'aib_1_bufchan_buf [0]);
  assign \v'aib_1_argbuf_d  = (\v'aib_1_bufchan_buf [0] ? \v'aib_1_bufchan_buf  :
                               \v'aib_1_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aib_1_bufchan_buf  <= {32'd0, 1'd0};
    else
      if ((\v'aib_1_argbuf_r  && \v'aib_1_bufchan_buf [0]))
        \v'aib_1_bufchan_buf  <= {32'd0, 1'd0};
      else if (((! \v'aib_1_argbuf_r ) && (! \v'aib_1_bufchan_buf [0])))
        \v'aib_1_bufchan_buf  <= \v'aib_1_bufchan_d ;
  
  /* fork (Ty Int) : (v'aib_destruct,Int) > [(v'aib_1,Int),
                                        (v'aib_2,Int)] */
  logic [1:0] \v'aib_destruct_emitted ;
  logic [1:0] \v'aib_destruct_done ;
  assign \v'aib_1_d  = {\v'aib_destruct_d [32:1],
                        (\v'aib_destruct_d [0] && (! \v'aib_destruct_emitted [0]))};
  assign \v'aib_2_d  = {\v'aib_destruct_d [32:1],
                        (\v'aib_destruct_d [0] && (! \v'aib_destruct_emitted [1]))};
  assign \v'aib_destruct_done  = (\v'aib_destruct_emitted  | ({\v'aib_2_d [0],
                                                               \v'aib_1_d [0]} & {\v'aib_2_r ,
                                                                                  \v'aib_1_r }));
  assign \v'aib_destruct_r  = (& \v'aib_destruct_done );
  always_ff @(posedge clk)
    if ((reset == 1'd1)) \v'aib_destruct_emitted  <= 2'd0;
    else
      \v'aib_destruct_emitted  <= (\v'aib_destruct_r  ? 2'd0 :
                                   \v'aib_destruct_done );
  
  /* buf (Ty Int) : (vai0_destruct,Int) > (vai0_1_argbuf,Int) */
  Int_t vai0_destruct_bufchan_d;
  logic vai0_destruct_bufchan_r;
  assign vai0_destruct_r = ((! vai0_destruct_bufchan_d[0]) || vai0_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai0_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vai0_destruct_r) vai0_destruct_bufchan_d <= vai0_destruct_d;
  Int_t vai0_destruct_bufchan_buf;
  assign vai0_destruct_bufchan_r = (! vai0_destruct_bufchan_buf[0]);
  assign vai0_1_argbuf_d = (vai0_destruct_bufchan_buf[0] ? vai0_destruct_bufchan_buf :
                            vai0_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai0_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vai0_1_argbuf_r && vai0_destruct_bufchan_buf[0]))
        vai0_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vai0_1_argbuf_r) && (! vai0_destruct_bufchan_buf[0])))
        vai0_destruct_bufchan_buf <= vai0_destruct_bufchan_d;
  
  /* buf (Ty Int) : (vai8_2_2,Int) > (vai8_2_2_argbuf,Int) */
  Int_t vai8_2_2_bufchan_d;
  logic vai8_2_2_bufchan_r;
  assign vai8_2_2_r = ((! vai8_2_2_bufchan_d[0]) || vai8_2_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_2_2_bufchan_d <= {32'd0, 1'd0};
    else if (vai8_2_2_r) vai8_2_2_bufchan_d <= vai8_2_2_d;
  Int_t vai8_2_2_bufchan_buf;
  assign vai8_2_2_bufchan_r = (! vai8_2_2_bufchan_buf[0]);
  assign vai8_2_2_argbuf_d = (vai8_2_2_bufchan_buf[0] ? vai8_2_2_bufchan_buf :
                              vai8_2_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_2_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vai8_2_2_argbuf_r && vai8_2_2_bufchan_buf[0]))
        vai8_2_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vai8_2_2_argbuf_r) && (! vai8_2_2_bufchan_buf[0])))
        vai8_2_2_bufchan_buf <= vai8_2_2_bufchan_d;
  
  /* fork (Ty Int) : (vai8_2_destruct,Int) > [(vai8_2_1,Int),
                                         (vai8_2_2,Int)] */
  logic [1:0] vai8_2_destruct_emitted;
  logic [1:0] vai8_2_destruct_done;
  assign vai8_2_1_d = {vai8_2_destruct_d[32:1],
                       (vai8_2_destruct_d[0] && (! vai8_2_destruct_emitted[0]))};
  assign vai8_2_2_d = {vai8_2_destruct_d[32:1],
                       (vai8_2_destruct_d[0] && (! vai8_2_destruct_emitted[1]))};
  assign vai8_2_destruct_done = (vai8_2_destruct_emitted | ({vai8_2_2_d[0],
                                                             vai8_2_1_d[0]} & {vai8_2_2_r,
                                                                               vai8_2_1_r}));
  assign vai8_2_destruct_r = (& vai8_2_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_2_destruct_emitted <= 2'd0;
    else
      vai8_2_destruct_emitted <= (vai8_2_destruct_r ? 2'd0 :
                                  vai8_2_destruct_done);
  
  /* buf (Ty Int) : (vai8_3_2,Int) > (vai8_3_2_argbuf,Int) */
  Int_t vai8_3_2_bufchan_d;
  logic vai8_3_2_bufchan_r;
  assign vai8_3_2_r = ((! vai8_3_2_bufchan_d[0]) || vai8_3_2_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_3_2_bufchan_d <= {32'd0, 1'd0};
    else if (vai8_3_2_r) vai8_3_2_bufchan_d <= vai8_3_2_d;
  Int_t vai8_3_2_bufchan_buf;
  assign vai8_3_2_bufchan_r = (! vai8_3_2_bufchan_buf[0]);
  assign vai8_3_2_argbuf_d = (vai8_3_2_bufchan_buf[0] ? vai8_3_2_bufchan_buf :
                              vai8_3_2_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_3_2_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vai8_3_2_argbuf_r && vai8_3_2_bufchan_buf[0]))
        vai8_3_2_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vai8_3_2_argbuf_r) && (! vai8_3_2_bufchan_buf[0])))
        vai8_3_2_bufchan_buf <= vai8_3_2_bufchan_d;
  
  /* fork (Ty Int) : (vai8_3_destruct,Int) > [(vai8_3_1,Int),
                                         (vai8_3_2,Int)] */
  logic [1:0] vai8_3_destruct_emitted;
  logic [1:0] vai8_3_destruct_done;
  assign vai8_3_1_d = {vai8_3_destruct_d[32:1],
                       (vai8_3_destruct_d[0] && (! vai8_3_destruct_emitted[0]))};
  assign vai8_3_2_d = {vai8_3_destruct_d[32:1],
                       (vai8_3_destruct_d[0] && (! vai8_3_destruct_emitted[1]))};
  assign vai8_3_destruct_done = (vai8_3_destruct_emitted | ({vai8_3_2_d[0],
                                                             vai8_3_1_d[0]} & {vai8_3_2_r,
                                                                               vai8_3_1_r}));
  assign vai8_3_destruct_r = (& vai8_3_destruct_done);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_3_destruct_emitted <= 2'd0;
    else
      vai8_3_destruct_emitted <= (vai8_3_destruct_r ? 2'd0 :
                                  vai8_3_destruct_done);
  
  /* buf (Ty Int) : (vai8_4_destruct,Int) > (vai8_4_1_argbuf,Int) */
  Int_t vai8_4_destruct_bufchan_d;
  logic vai8_4_destruct_bufchan_r;
  assign vai8_4_destruct_r = ((! vai8_4_destruct_bufchan_d[0]) || vai8_4_destruct_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_4_destruct_bufchan_d <= {32'd0, 1'd0};
    else
      if (vai8_4_destruct_r)
        vai8_4_destruct_bufchan_d <= vai8_4_destruct_d;
  Int_t vai8_4_destruct_bufchan_buf;
  assign vai8_4_destruct_bufchan_r = (! vai8_4_destruct_bufchan_buf[0]);
  assign vai8_4_1_argbuf_d = (vai8_4_destruct_bufchan_buf[0] ? vai8_4_destruct_bufchan_buf :
                              vai8_4_destruct_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) vai8_4_destruct_bufchan_buf <= {32'd0, 1'd0};
    else
      if ((vai8_4_1_argbuf_r && vai8_4_destruct_bufchan_buf[0]))
        vai8_4_destruct_bufchan_buf <= {32'd0, 1'd0};
      else if (((! vai8_4_1_argbuf_r) && (! vai8_4_destruct_bufchan_buf[0])))
        vai8_4_destruct_bufchan_buf <= vai8_4_destruct_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (lizzieLet13_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet13_1_argbuf_d = (writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf :
                                   writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((lizzieLet13_1_argbuf_r && writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! lizzieLet13_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet0_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet20_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet20_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet20_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet20_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca2_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_1_argbuf_d = (writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca2_1_argbuf_r && writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca2_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet20_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet21_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet21_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet21_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet21_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca1_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_1_argbuf_d = (writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca1_1_argbuf_r && writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca1_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet21_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet22_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet22_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet22_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf :
                                                       writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet22_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca0_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_1_argbuf_d = (writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((sca0_1_argbuf_r && writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! sca0_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet22_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf,Pointer_CT$wnnz_Int) > (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]);
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf :
                                                      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CT$wnnz_Int) : (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb,Pointer_CT$wnnz_Int) > (sca3_1_argbuf,Pointer_CT$wnnz_Int) */
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  logic writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r = ((! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d[0]) || writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_r)
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_d;
  Pointer_CT$wnnz_Int_t writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf;
  assign writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_r = (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_1_argbuf_d = (writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0] ? writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf :
                            writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                              1'd0};
    else
      if ((sca3_1_argbuf_r && writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0]))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                1'd0};
      else if (((! sca3_1_argbuf_r) && (! writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf[0])))
        writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_buf <= writeCT$wnnz_IntlizzieLet5_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > (writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d  <= {16'd0,
                                                                         1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_d  = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf  :
                                                                       \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
    else
      if ((\writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_r  && \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf  <= {16'd0,
                                                                             1'd0};
      else if (((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_r ) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) > (sca3_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                             1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf [0]);
  assign sca3_1_1_argbuf_d = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
    else
      if ((sca3_1_1_argbuf_r && \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                                 1'd0};
      else if (((! sca3_1_1_argbuf_r) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet11_2_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > (writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_d  = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf  :
                                                                     \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((\writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_r  && \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_r ) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) > (lizzieLet6_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf [0]);
  assign lizzieLet6_1_1_argbuf_d = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf  :
                                    \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((lizzieLet6_1_1_argbuf_r && \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! lizzieLet6_1_1_argbuf_r) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet17_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > (writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_d  = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  :
                                                                     \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((\writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_r  && \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_r ) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) > (sca2_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0]);
  assign sca2_1_1_argbuf_d = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((sca2_1_1_argbuf_r && \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! sca2_1_1_argbuf_r) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet24_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > (writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_d  = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  :
                                                                     \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((\writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_r  && \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_r ) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) > (sca1_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0]);
  assign sca1_1_1_argbuf_d = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((sca1_1_1_argbuf_r && \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! sca1_1_1_argbuf_r) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet25_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) > (writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d  <= {16'd0,
                                                                       1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf [0]);
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_d  = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf  :
                                                                     \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf  <= {16'd0,
                                                                         1'd0};
    else
      if ((\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_r  && \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf  <= {16'd0,
                                                                           1'd0};
      else if (((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_r ) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_bufchan_d ;
  
  /* buf (Ty Pointer_CTf'_f'_Int_Int_Int_Int) : (writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb,Pointer_CTf'_f'_Int_Int_Int_Int) > (sca0_1_1_argbuf,Pointer_CTf'_f'_Int_Int_Int_Int) */
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d ;
  logic \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_r ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_r  = ((! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d [0]) || \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_r );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d  <= {16'd0,
                                                                           1'd0};
    else
      if (\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_r )
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_d ;
  \Pointer_CTf'_f'_Int_Int_Int_Int_t  \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf ;
  assign \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_r  = (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf [0]);
  assign sca0_1_1_argbuf_d = (\writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf [0] ? \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf  :
                              \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d );
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                             1'd0};
    else
      if ((sca0_1_1_argbuf_r && \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf [0]))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf  <= {16'd0,
                                                                               1'd0};
      else if (((! sca0_1_1_argbuf_r) && (! \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf [0])))
        \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_buf  <= \writeCTf'_f'_Int_Int_Int_IntlizzieLet26_1_argbuf_rwb_bufchan_d ;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_d = (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf :
                                                                 writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_r && writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) > (sca3_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]);
  assign sca3_2_1_argbuf_d = (writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((sca3_2_1_argbuf_r && writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! sca3_2_1_argbuf_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet15_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_d = (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf :
                                                                 writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_r && writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) > (lizzieLet10_1_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet10_1_1_argbuf_d = (writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf :
                                     writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((lizzieLet10_1_1_argbuf_r && writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! lizzieLet10_1_1_argbuf_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet18_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_d = (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf :
                                                                 writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_r && writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) > (sca2_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]);
  assign sca2_2_1_argbuf_d = (writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((sca2_2_1_argbuf_r && writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! sca2_2_1_argbuf_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet29_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_d = (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf :
                                                                 writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_r && writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) > (sca1_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]);
  assign sca1_2_1_argbuf_d = (writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((sca1_2_1_argbuf_r && writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! sca1_2_1_argbuf_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet30_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) > (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= {16'd0,
                                                                   1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]);
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_d = (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf :
                                                                 writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                     1'd0};
    else
      if ((writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_r && writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= {16'd0,
                                                                       1'd0};
      else if (((! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_CTf_f_Int_Int_Int_Int) : (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb,Pointer_CTf_f_Int_Int_Int_Int) > (sca0_2_1_argbuf,Pointer_CTf_f_Int_Int_Int_Int) */
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  logic writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_r = ((! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d[0]) || writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                                       1'd0};
    else
      if (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_r)
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d <= writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_d;
  Pointer_CTf_f_Int_Int_Int_Int_t writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf;
  assign writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_r = (! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]);
  assign sca0_2_1_argbuf_d = (writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0] ? writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf :
                              writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                         1'd0};
    else
      if ((sca0_2_1_argbuf_r && writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0]))
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                           1'd0};
      else if (((! sca0_2_1_argbuf_r) && (! writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf[0])))
        writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_buf <= writeCTf_f_Int_Int_Int_IntlizzieLet31_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_r = ((! writeQTree_IntlizzieLet10_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_r)
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_d = (writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet10_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet10_1_argbuf_rwb_r && writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet10_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet10_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet4_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet10_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet10_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet4_1_1_argbuf_d = (writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet4_1_1_argbuf_r && writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet4_1_1_argbuf_r) && (! writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet10_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_r = ((! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_1_argbuf_r)
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet12_1_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d = (writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf :
                                                       writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r && writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet12_1_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet12_1_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet5_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d <= {16'd0,
                                                             1'd0};
    else
      if (writeQTree_IntlizzieLet12_1_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet12_1_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet5_1_1_argbuf_d = (writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
    else
      if ((lizzieLet5_1_1_argbuf_r && writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                                 1'd0};
      else if (((! lizzieLet5_1_1_argbuf_r) && (! writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet12_1_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet14_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_argbuf_r = ((! writeQTree_IntlizzieLet14_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_argbuf_r)
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet14_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_d = (writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet14_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet14_1_argbuf_rwb_r && writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet14_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet14_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet14_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet7_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet14_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet14_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet7_1_1_argbuf_d = (writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet7_1_1_argbuf_r && writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet7_1_1_argbuf_r) && (! writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet14_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_r = ((! writeQTree_IntlizzieLet16_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_r)
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_d = (writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet16_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet16_1_argbuf_rwb_r && writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet16_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet16_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet9_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet16_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet16_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet9_1_1_argbuf_d = (writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((lizzieLet9_1_1_argbuf_r && writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! lizzieLet9_1_1_argbuf_r) && (! writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet16_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet27_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet27_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet27_1_argbuf_r = ((! writeQTree_IntlizzieLet27_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet27_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet27_1_argbuf_r)
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet27_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet27_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_d = (writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet27_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet27_1_argbuf_rwb_r && writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet27_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet27_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet27_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet27_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet27_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet27_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_1_1_argbuf_d = (writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_1_1_argbuf_r && writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_1_1_argbuf_r) && (! writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet27_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_r = ((! writeQTree_IntlizzieLet32_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_r)
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_d = (writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf :
                                                     writeQTree_IntlizzieLet32_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet32_1_argbuf_rwb_r && writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet32_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet32_1_argbuf_rwb,Pointer_QTree_Int) > (contRet_0_2_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet32_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet32_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]);
  assign contRet_0_2_1_argbuf_d = (writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf :
                                   writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                             1'd0};
    else
      if ((contRet_0_2_1_argbuf_r && writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= {16'd0,
                                                               1'd0};
      else if (((! contRet_0_2_1_argbuf_r) && (! writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet32_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_r = ((! writeQTree_IntlizzieLet7_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_r)
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_d = (writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet7_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet7_1_argbuf_rwb_r && writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet7_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet7_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet1_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet7_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet7_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet1_1_1_argbuf_d = (writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet1_1_1_argbuf_r && writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet1_1_1_argbuf_r) && (! writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet7_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_r = ((! writeQTree_IntlizzieLet8_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_r)
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_d = (writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet8_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet8_1_argbuf_rwb_r && writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet8_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet8_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet2_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet8_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet8_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet2_1_1_argbuf_d = (writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet2_1_1_argbuf_r && writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet2_1_1_argbuf_r) && (! writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet8_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf,Pointer_QTree_Int) > (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_r = ((! writeQTree_IntlizzieLet9_1_argbuf_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_r)
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]);
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_d = (writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf :
                                                    writeQTree_IntlizzieLet9_1_argbuf_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((writeQTree_IntlizzieLet9_1_argbuf_rwb_r && writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= {16'd0, 1'd0};
      else if (((! writeQTree_IntlizzieLet9_1_argbuf_rwb_r) && (! writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (writeQTree_IntlizzieLet9_1_argbuf_rwb,Pointer_QTree_Int) > (lizzieLet3_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  logic writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_r = ((! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d[0]) || writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= {16'd0, 1'd0};
    else
      if (writeQTree_IntlizzieLet9_1_argbuf_rwb_r)
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d <= writeQTree_IntlizzieLet9_1_argbuf_rwb_d;
  Pointer_QTree_Int_t writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf;
  assign writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_r = (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]);
  assign lizzieLet3_1_1_argbuf_d = (writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0] ? writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf :
                                    writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((lizzieLet3_1_1_argbuf_r && writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0]))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= {16'd0, 1'd0};
      else if (((! lizzieLet3_1_1_argbuf_r) && (! writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf[0])))
        writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_buf <= writeQTree_IntlizzieLet9_1_argbuf_rwb_bufchan_d;
  
  /* buf (Ty Pointer_QTree_Int) : (wstH_1_goMux_mux,Pointer_QTree_Int) > (wstH_1_1_argbuf,Pointer_QTree_Int) */
  Pointer_QTree_Int_t wstH_1_goMux_mux_bufchan_d;
  logic wstH_1_goMux_mux_bufchan_r;
  assign wstH_1_goMux_mux_r = ((! wstH_1_goMux_mux_bufchan_d[0]) || wstH_1_goMux_mux_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wstH_1_goMux_mux_bufchan_d <= {16'd0, 1'd0};
    else
      if (wstH_1_goMux_mux_r)
        wstH_1_goMux_mux_bufchan_d <= wstH_1_goMux_mux_d;
  Pointer_QTree_Int_t wstH_1_goMux_mux_bufchan_buf;
  assign wstH_1_goMux_mux_bufchan_r = (! wstH_1_goMux_mux_bufchan_buf[0]);
  assign wstH_1_1_argbuf_d = (wstH_1_goMux_mux_bufchan_buf[0] ? wstH_1_goMux_mux_bufchan_buf :
                              wstH_1_goMux_mux_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1)) wstH_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
    else
      if ((wstH_1_1_argbuf_r && wstH_1_goMux_mux_bufchan_buf[0]))
        wstH_1_goMux_mux_bufchan_buf <= {16'd0, 1'd0};
      else if (((! wstH_1_1_argbuf_r) && (! wstH_1_goMux_mux_bufchan_buf[0])))
        wstH_1_goMux_mux_bufchan_buf <= wstH_1_goMux_mux_bufchan_d;
  
  /* buf (Ty CT$wnnz_Int) : (wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) > (lizzieLet21_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d;
  logic wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_r;
  assign wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_r = ((! wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d[0]) || wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d <= {115'd0,
                                                                                              1'd0};
    else
      if (wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_r)
        wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d <= wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_d;
  CT$wnnz_Int_t wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf;
  assign wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_r = (! wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf[0]);
  assign lizzieLet21_1_argbuf_d = (wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf[0] ? wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf :
                                   wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                1'd0};
    else
      if ((lizzieLet21_1_argbuf_r && wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf[0]))
        wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf <= {115'd0,
                                                                                                  1'd0};
      else if (((! lizzieLet21_1_argbuf_r) && (! wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf[0])))
        wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_buf <= wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int1) : [(wwstK_2_destruct,Int#),
                                (lizzieLet19_4Lcall_$wnnz_Int2,Int#),
                                (sc_0_4_destruct,Pointer_CT$wnnz_Int),
                                (q4abZ_2_destruct,Pointer_QTree_Int)] > (wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1,CT$wnnz_Int) */
  assign wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_d = Lcall_$wnnz_Int1_dc((& {wwstK_2_destruct_d[0],
                                                                                                               lizzieLet19_4Lcall_$wnnz_Int2_d[0],
                                                                                                               sc_0_4_destruct_d[0],
                                                                                                               q4abZ_2_destruct_d[0]}), wwstK_2_destruct_d, lizzieLet19_4Lcall_$wnnz_Int2_d, sc_0_4_destruct_d, q4abZ_2_destruct_d);
  assign {wwstK_2_destruct_r,
          lizzieLet19_4Lcall_$wnnz_Int2_r,
          sc_0_4_destruct_r,
          q4abZ_2_destruct_r} = {4 {(wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_r && wwstK_2_1lizzieLet19_4Lcall_$wnnz_Int2_1sc_0_4_1q4abZ_2_1Lcall_$wnnz_Int1_d[0])}};
  
  /* buf (Ty CT$wnnz_Int) : (wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0,CT$wnnz_Int) > (lizzieLet22_1_argbuf,CT$wnnz_Int) */
  CT$wnnz_Int_t wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d;
  logic wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_r;
  assign wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_r = ((! wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d[0]) || wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_r);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d <= {115'd0,
                                                                                               1'd0};
    else
      if (wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_r)
        wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d <= wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_d;
  CT$wnnz_Int_t wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf;
  assign wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_r = (! wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf[0]);
  assign lizzieLet22_1_argbuf_d = (wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf[0] ? wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf :
                                   wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d);
  always_ff @(posedge clk)
    if ((reset == 1'd1))
      wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                 1'd0};
    else
      if ((lizzieLet22_1_argbuf_r && wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf[0]))
        wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf <= {115'd0,
                                                                                                   1'd0};
      else if (((! lizzieLet22_1_argbuf_r) && (! wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf[0])))
        wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_buf <= wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_bufchan_d;
  
  /* dcon (Ty CT$wnnz_Int,
      Dcon Lcall_$wnnz_Int0) : [(wwstK_3_destruct,Int#),
                                (ww1XuL_1_destruct,Int#),
                                (lizzieLet19_4Lcall_$wnnz_Int1,Int#),
                                (sc_0_5_destruct,Pointer_CT$wnnz_Int)] > (wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0,CT$wnnz_Int) */
  assign wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_d = Lcall_$wnnz_Int0_dc((& {wwstK_3_destruct_d[0],
                                                                                                                ww1XuL_1_destruct_d[0],
                                                                                                                lizzieLet19_4Lcall_$wnnz_Int1_d[0],
                                                                                                                sc_0_5_destruct_d[0]}), wwstK_3_destruct_d, ww1XuL_1_destruct_d, lizzieLet19_4Lcall_$wnnz_Int1_d, sc_0_5_destruct_d);
  assign {wwstK_3_destruct_r,
          ww1XuL_1_destruct_r,
          lizzieLet19_4Lcall_$wnnz_Int1_r,
          sc_0_5_destruct_r} = {4 {(wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_r && wwstK_3_1ww1XuL_1_1lizzieLet19_4Lcall_$wnnz_Int1_1sc_0_5_1Lcall_$wnnz_Int0_d[0])}};
  
  /* op_add (Ty Int#) : (wwstK_4_1ww1XuL_2_1_Add32,Int#) (ww2XuO_1_destruct,Int#) > (es_6_2_1ww2XuO_1_1_Add32,Int#) */
  assign es_6_2_1ww2XuO_1_1_Add32_d = {(wwstK_4_1ww1XuL_2_1_Add32_d[32:1] + ww2XuO_1_destruct_d[32:1]),
                                       (wwstK_4_1ww1XuL_2_1_Add32_d[0] && ww2XuO_1_destruct_d[0])};
  assign {wwstK_4_1ww1XuL_2_1_Add32_r,
          ww2XuO_1_destruct_r} = {2 {(es_6_2_1ww2XuO_1_1_Add32_r && es_6_2_1ww2XuO_1_1_Add32_d[0])}};
  
  /* op_add (Ty Int#) : (wwstK_4_destruct,Int#) (ww1XuL_2_destruct,Int#) > (wwstK_4_1ww1XuL_2_1_Add32,Int#) */
  assign wwstK_4_1ww1XuL_2_1_Add32_d = {(wwstK_4_destruct_d[32:1] + ww1XuL_2_destruct_d[32:1]),
                                        (wwstK_4_destruct_d[0] && ww1XuL_2_destruct_d[0])};
  assign {wwstK_4_destruct_r,
          ww1XuL_2_destruct_r} = {2 {(wwstK_4_1ww1XuL_2_1_Add32_r && wwstK_4_1ww1XuL_2_1_Add32_d[0])}};
  
  /* dcon (Ty Int,
      Dcon I#) : [(xap7_1lizzieLet0_1_1_Add32,Int#)] > (es_0_1_1I#,Int) */
  assign \es_0_1_1I#_d  = \I#_dc ((& {xap7_1lizzieLet0_1_1_Add32_d[0]}), xap7_1lizzieLet0_1_1_Add32_d);
  assign {xap7_1lizzieLet0_1_1_Add32_r} = {1 {(\es_0_1_1I#_r  && \es_0_1_1I#_d [0])}};
  
  /* op_add (Ty Int#) : (xap7_destruct,Int#) (arg0_2_1Dcon_main1_3I#_1_argbuf_2,Int#) > (xap7_1lizzieLet0_1_1_Add32,Int#) */
  assign xap7_1lizzieLet0_1_1_Add32_d = {(xap7_destruct_d[32:1] + \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [32:1]),
                                         (xap7_destruct_d[0] && \arg0_2_1Dcon_main1_3I#_1_argbuf_2_d [0])};
  assign {xap7_destruct_r,
          \arg0_2_1Dcon_main1_3I#_1_argbuf_2_r } = {2 {(xap7_1lizzieLet0_1_1_Add32_r && xap7_1lizzieLet0_1_1_Add32_d[0])}};
endmodule